PK                      checkpoint/data.pklFB ZZZZZZZZZZZ�}q (X   epochqM�X	   optimizerq}q(X   stateq}q(K }q(X   stepqctorch._utils
_rebuild_tensor_v2
q((X   storageq	ctorch
FloatStorage
q
X   0qX   cpuqKtqQK ))�ccollections
OrderedDict
q)RqtqRqX   exp_avgqh((h	h
X   1qhM�tqQK K9K�qKK�q�h)RqtqRqX
   exp_avg_sqqh((h	h
X   2qhM�tqQK K9K�qKK�q�h)Rqtq Rq!uK}q"(hh((h	h
X   3q#hKtq$QK ))�h)Rq%tq&Rq'hh((h	h
X   4q(hMStq)QK KKK�q*KK�q+�h)Rq,tq-Rq.hh((h	h
X   5q/hMStq0QK KKK�q1KK�q2�h)Rq3tq4Rq5uK}q6(hh((h	h
X   6q7hKtq8QK ))�h)Rq9tq:Rq;hh((h	h
X   7q<hKKtq=QK KK�q>K�q?�h)Rq@tqARqBhh((h	h
X   8qChKKtqDQK KK�qEK�qF�h)RqGtqHRqIuK}qJ(hh((h	h
X   9qKhKtqLQK ))�h)RqMtqNRqOhh((h	h
X   10qPhMqtqQQK KK�qRKK�qS�h)RqTtqURqVhh((h	h
X   11qWhMqtqXQK KK�qYKK�qZ�h)Rq[tq\Rq]uK}q^(hh((h	h
X   12q_hKtq`QK ))�h)RqatqbRqchh((h	h
X   13qdhKtqeQK K�qfK�qg�h)RqhtqiRqjhh((h	h
X   14qkhKtqlQK K�qmK�qn�h)RqotqpRqquK}qr(hh((h	h
X   15qshKtqtQK ))�h)RqutqvRqwhh((h	h
X   16qxhJH� tqyQK M�K��qzK�K�q{�h)Rq|tq}Rq~hh((h	h
X   17qhJH� tq�QK M�K��q�K�K�q��h)Rq�tq�Rq�uK}q�(hh((h	h
X   18q�hKtq�QK ))�h)Rq�tq�Rq�hh((h	h
X   19q�hM�tq�QK M��q�K�q��h)Rq�tq�Rq�hh((h	h
X   20q�hM�tq�QK M��q�K�q��h)Rq�tq�Rq�uK}q�(hh((h	h
X   21q�hKtq�QK ))�h)Rq�tq�Rq�hh((h	h
X   22q�hM�tq�QK M��q�K�q��h)Rq�tq�Rq�hh((h	h
X   23q�hM�tq�QK M��q�K�q��h)Rq�tq�Rq�uK}q�(hh((h	h
X   24q�hKtq�QK ))�h)Rq�tq�Rq�hh((h	h
X   25q�hM�tq�QK M��q�K�q��h)Rq�tq�Rq�hh((h	h
X   26q�hM�tq�QK M��q�K�q��h)Rq�tq�Rq�uK	}q�(hh((h	h
X   27q�hKtq�QK ))�h)Rq�tq�Rq�hh((h	h
X   28q�hMTotq�QK K9M��q�M�K�qˉh)Rq�tq�Rq�hh((h	h
X   29q�hMTotq�QK K9M��q�M�K�q҉h)Rq�tq�Rq�uK
}q�(hh((h	h
X   30q�hKtq�QK ))�h)Rq�tq�Rq�hh((h	h
X   31q�hK9tq�QK K9�q�K�q߉h)Rq�tq�Rq�hh((h	h
X   32q�hK9tq�QK K9�q�K�q�h)Rq�tq�Rq�uuX   param_groupsq�]q�}q�(X   lrq�G?PbM���X   betasq�G?�������G?�����+�q�X   epsq�G>Ey��0�:X   weight_decayq�K X   amsgradq�X   maximizeq�X   foreachq�NX
   capturableq��X   differentiableq��X   fusedq�NX   paramsq�]q�(K KKKKKKKKK	K
euauX   model_state_dictq�h)Rq�(X   input_embeddings.weightq�h((h	h
X   33q�hM�tq�QK K9K�q�KK�r   �h)Rr  tr  Rr  X"   attention.attention.in_proj_weightr  h((h	h
X   34r  hMStr  QK KKK�r  KK�r  �h)Rr	  tr
  Rr  X    attention.attention.in_proj_biasr  h((h	h
X   35r  hKKtr  QK KK�r  K�r  �h)Rr  tr  Rr  X#   attention.attention.out_proj.weightr  h((h	h
X   36r  hMqtr  QK KK�r  KK�r  �h)Rr  tr  Rr  X!   attention.attention.out_proj.biasr  h((h	h
X   37r  hKtr  QK K�r  K�r   �h)Rr!  tr"  Rr#  X   linear.weightr$  h((h	h
X   38r%  hJH� tr&  QK M�K��r'  K�K�r(  �h)Rr)  tr*  Rr+  X   linear.biasr,  h((h	h
X   39r-  hM�tr.  QK M��r/  K�r0  �h)Rr1  tr2  Rr3  X   normalize.weightr4  h((h	h
X   40r5  hM�tr6  QK M��r7  K�r8  �h)Rr9  tr:  Rr;  X   normalize.biasr<  h((h	h
X   41r=  hM�tr>  QK M��r?  K�r@  �h)RrA  trB  RrC  X   output.weightrD  h((h	h
X   42rE  hMTotrF  QK K9M��rG  M�K�rH  �h)RrI  trJ  RrK  X   output.biasrL  h((h	h
X   43rM  hK9trN  QK K9�rO  K�rP  �h)RrQ  trR  RrS  u}rT  X	   _metadatarU  h)RrV  (X    rW  }rX  X   versionrY  KsX   input_embeddingsrZ  }r[  jY  KsX	   attentionr\  }r]  jY  KsX   attention.attentionr^  }r_  jY  KsX   attention.attention.out_projr`  }ra  jY  KsX   flattenrb  }rc  jY  KsX   linearrd  }re  jY  KsX	   normalizerf  }rg  jY  KsX
   activationrh  }ri  jY  KsX   outputrj  }rk  jY  KsusbX   token_decoderrl  }rm  (K X   
rn  KX    ro  KX   !rp  KX   'rq  KX   ,rr  KX   -rs  KX   .rt  KX   :ru  KX   ;rv  K	X   ?rw  K
X   Arx  KX   Bry  KX   Crz  KX   Dr{  KX   Er|  KX   Fr}  KX   Hr~  KX   Ir  KX   Jr�  KX   Lr�  KX   Mr�  KX   Nr�  KX   Or�  KX   Pr�  KX   Rr�  KX   Sr�  KX   Tr�  KX   Ur�  KX   Vr�  KX   Wr�  KX   Yr�  KX   ar�  K X   br�  K!X   cr�  K"X   dr�  K#X   er�  K$X   fr�  K%X   gr�  K&X   hr�  K'X   ir�  K(X   jr�  K)X   kr�  K*X   lr�  K+X   mr�  K,X   nr�  K-X   or�  K.X   pr�  K/X   qr�  K0X   rr�  K1X   sr�  K2X   tr�  K3X   ur�  K4X   vr�  K5X   wr�  K6X   xr�  K7X   yr�  K8X   zr�  uX   char_encoderr�  }r�  (jn  K jo  Kjp  Kjq  Kjr  Kjs  Kjt  Kju  Kjv  Kjw  K	jx  K
jy  Kjz  Kj{  Kj|  Kj}  Kj~  Kj  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  Kj�  K j�  K!j�  K"j�  K#j�  K$j�  K%j�  K&j�  K'j�  K(j�  K)j�  K*j�  K+j�  K,j�  K-j�  K.j�  K/j�  K0j�  K1j�  K2j�  K3j�  K4j�  K5j�  K6j�  K7j�  K8uX   hyperparametersr�  }r�  (X   context_lengthr�  K
X   embedding_dimr�  KX   n_tokensr�  K9X   n_attn_headsr�  KX	   n_neuronsr�  M�uu.PKr�?m      PK                      checkpoint/byteorderFB ZZZZZZZZZZZZZZZZZZZZZZZZZZlittlePK�=�      PK                     ; checkpoint/data/0FB7 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     = checkpoint/data/1FB9 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�q6�6�6 ��2M߆6Bku6H�;�@�
�H��t�6��6FMO6���5dĶ4��ɵ�G�6��!�6$m�� ?r�N}7�64��5c@(6Z�
7܎d����7�`)�>�71�8<^1��T���o�6��з;�6���6�`�7���75�m7�7
(-7��߶
�H���6��ҷ��ӷP�t��J7�& 8�{7��η(7�!z�@c1�v ���̳��3 U4��4����"4���v����D��[��4��x��3{��4j��@�³��0�)4Jڳ�"���<�j�}�]�%��9E�b�3���Y�w5&*�4�<5�i�42���sf����w�h��53�l��O4��T5.QC5��쵱$5G` 5�Ȱ�Ic������z�5�:��vɳ5�o"��6X\����k6B��ح�5c�6`+J4�	5�{6��:�!q��ص���6
-Q��{�5\8�5�(��1�2�W`6� 6�r56G�����16�rܳJ�)�m6��X|$�@�|����TV�4w4E�54���nNo5_y5�ͳѥ�4����ӡ���n]��s
��ߘ��G����H�>��-5��ʴJ�5�7δ��A30|^�j
���\^�J����0��r��3�5����|��5?� ��[n5�54,05D5�w75� ����@���z�/6���5�2I��ۿ����ݼ5��54ʞ�����*6yQN6�\ٵ���5��ȵ��i5�K$6�ص5�J7�]��9M6I�t���5Z�U6~���"��4 I��&V��`�"�B�2��4ku����ֳ ��1��0��wo2�y�}^����5lQ23���4�ܳ��3
e�4�Xb1��4�E���X��0�A�e��4i	��0)4�K3�y�J�06����0�5�'-�]����dʵ�C���H58����6�O� �5Wµ}j��c�TFS�Vf���ڢ5 x�����3J\5��D5�ά�P"4��tU�$��4�b�wE��W�4⮘5�E$5,Ѵ���5�.����1Ϻ5<�5����n5Z��4,tq�5Z��)ʵ2��4�0�c����"�5���f��4���4(�4��Yͳ���1�-'�,oL�����7��Vf4�FP2�MY��%3%��3 ��3�'n���3}�0����h�����zk-3��I��*���IJ4\/�3 �!4�_�~߽5��5�RW6�H�6GZ 6�{"��b�����L�Y���%�x�4���ؐ���$66y
��w���z�G�n5 �����t6�D�6K#��䡏���|�w>�2Y���N^3�4r3��t\���31ɟL�G���Td���2M �3.J2��W3R�W��m3����t�F�.��2�v���\�2tE3�;2�_-3�阱�u�5����	�5G[�D2�5���l{�.k�B�$�'_66x�T�v�򵒮�3&յ������^�5Z*�5C	4�d6�
rõ�65O�96��6������?�4������C4�C&3�ճ̥�Gf
� w�������ߴtT�4�5��[��u��3����L_4�5u4w.�4�^ܳ�M���g4�����.�� ��4�[(�o-�ϒ۴,����
�&5�5�>�`i��<�4��5}�?5��2A�5넶��-q���:5o� 4E6�4-&�WM46ą��%�a��o�5�ܾ5_>I�ɦ�D��>��5� 6.�85���V1���4T06�U��3�/���2��&t75��ݵ�j�����)W�H�H5<9���=���ߵ��(����5��]�Q��5s��2FT��.����K1Ҥ�2����¾X�~q	3�ӱR�2j�V��!��"5�1
�k1���2�Y�0�.2v�;�7�26T�2Yk3��3@�+�P�Y2u�N3��2XU�04ޝ�MyP3�Q���j���1���"س�ѥ3�D�1�������1��]2��J3�ب�|=�333�[�3�(��W�3\�˳Ð2�2Y�'N�3�ޙ5Oʙ5���L�vfX�S�5�W�5΄5���"�5�ϵ9t/���5ݏ�5� �"�85�W5�\�3L�5��C5��4�C���`�i��4����06�A 3-�X6����f�6�!�5�b���6V�6�n�5P�@6&F� ��1S�˵,��5�����M5:��5�޾5���5!��5��43�)5�c(6^-��>�sZ����4��j5�F�҉F5�a36r������g45�4�ꑳf�"�wA�5CN��.�`5ܱ15�o4"��Nz��ĸl5t���&6�`5F�z�N�3�Ͳ���2ó��rd3%��2Ь�o?x�b/�2�3_3��R����2ª�]m�2��2����35��ƅ2���1�:3�*3��j����2ѿk2L�&12D�	��F �J,=5b�\4rF���`�K�5o��h�4����w$��)X�X��5Ⱥ�4�R��^�4`�5	�ⵘA.�^6�!>s�9��5fB5.��õ��˵�����K��x-)6H?`6��7�Z=85 U65Rҙ����5�~5���3(�5��6֌�5��4��M6�n5(逴N���0C6���5T� 5�;Q6�LH6j��5yI�5H��5�5Q���"m�5 �ߴ�6̧*�l�ն<T�5v{�5��6�	,��gG6x��5��M�`w��5[6�ŷ5LU^6F�$6|J)�M�^��Ԉ5�
�@8��~�5�:6A�ڵ�q�4n0$4]�44<*5[A�5/�5��n��w��������6'��5R�I���!6�)��.}$�R4�#еP]�4�/�2}�3ST�24Y����ϲ� ���ʙ��Q�2:�����
g��<`�3�p�3�.�3�f�3"%i�ĕ63ڌ���+�3��y28v�ўL��3�O�S����2p� 6L��5p��Z��6^= ��(��´�n
5�t�5Ȥp�����B�Gj6�!&6��6�۵�6p��N+���ҍ����46+����5�?7��K����S�9SųU�4m��	�ֲ��t4~�մ�r4���4�ޱ�f"����3x;	4�Qo�A�3�;5���@�$���>5(����G�vmv�v�4[{54��t4��Z7��O�!��Q$�"�7`��4���6wC�6��-�x����XF7L�H�PT�5�ϛ��4�6��6J����N���77��7��&7���@�61���5({��7bO�����M�4��`3�6��5'Ie�jo�������紎� 70J�6A�׵�o�4U�����5tc6T^6�f:6Kܭ3M�Y��f��k�Y6�M�6_�J�x6�Ȓ5�Nw��������յ�X޶�����C�6��7���6�>9��0ʶ 7j��6e�J���z6�qk3��ӵ��4h[� ���P�4X��Q8P�~���d�6���6��46�6`�6x�2d96��}6��6l}e���5��/6GP �ܶ2�&T���-�5�[��@5�{��h��6��6"�ѶF6�Ŕ�2T��"� ���i5�4� �3"��6h3�Z�>6�)�6�`7.�|6i��6�V7���������l6xF�5�]K7�8����7�>��H����Q6LW~��<���,�������8�r�6��5;���0�5��6f�4���hd�5L!�����[��5\n85d���u�6U�C6�m���ӵ?]1�Z����궼k�6x��5��4���5ᜁ�"�����y5z�
ͽ5N&n6�蟶�[�5��5�+�6�>x4('���Nc�5!4vԙ6��6h�&�ɔ��|_E6&�E7 �e3�%6�@4���6�����k�6@s5|���N6�C�����3H?���޶�F�6F��5��6&
�6�u6�w����5�8�5�E����ٵ����ӶF��x�6���5���6�̂��T6�6��zU�5BB �45k�h�w6�,T57�����5�H����5�6>ܣ��j6(��x�k�TR����xܵ6ͮ�3�=ڲ ��4��3��'3<�3����;2Pj3,���k�2$F1����2��۲*S 3rSV3�̲T�S�/I����C��,���Բ9Z3�Z����A���4��4�д�՘��a)4���4���4TDӳ���s�� ��l]� �4����U�����\�o3)�д�%'�A54A&�k�5��B5�Z13���5�j6?�׵�\4�2��|R6��u��؁6��5���5b��68z�R�4�N�7Μ6 6� �P1~�\�]\L�!��06RӀ5��	6Dr��9þ��Y�����wr�5��%5��6���hѳ3"��4 �)��66S���	6�x�5��*��@�5*T!�C�:�wZF6��5y�ڪ����v���5H76�e��ּ5�R��l�D��I�5��6��6�S6>%!�� 7P�6:��6,�6^+ٶD	�~#=7297�g����F�(��p�=�!`G�1h��m�����66���k�7�Y\�Ʈ6��6ݟ�fw6�	�60L7��6�2z7ʣH��c�����Z�Ƕ~�ٶ|
*5`�
5T���W7���6�!���6b��6���-!�5`}�4 �"���un�����5�>A5���5��5	��4��5�G�4?��5�$�TK5��P��[6��6��׵p��H[u��l��r�>5<<23���a�F�v&�3�2u�t2�� ��г�����>�30��'��3_O���D(4��T3�T;4SY�^d����s13U*�"ז��C��?; 3br4;�3�~0(y��ʴ�6���4�e���;5��Ƕ�e��նY�7�t60a�6 �X7)(�`��4�X�J'��������������s68���y�5�O6�2�H̴67���"6���5��4�8��6�
7����v��6��7^���O����6e�:7�d�[~����5[�6��(��ET�x�w6\ɯ5�ў���X7�x9����5��*�W����6��f6���'Q��_3�!�^���N x�ny7�D7a��6�!�Py�>���5�=�6��"6��0��G�M�7�B�7{/�6�D5t��� Ѳ��w6Sr4�H��5�~�6��)6�z5#O6�Kd��+�4񉴼�O�{ؼ��r�4�M]6��b4�}\5b'F�с��hk6�6P�'�P�;�2�q5�2�4� 6Ĕ�5�� �e6R���(6�����w]�|���\a�XW1����4�j�@Kl3��5��54�	�5�������5:.�>9�5��\�)��FV5��:6t���̰5d冴��ϵ��3\g#62��5 Ҝ��d�Al�6��)��L�5�I�55��6 /6Ԇ��è�=C6�ە�>�N5~V��<2�v&3d�@��>j���C2`�23�h�3��3t(o��w3�#4��J3TG������T�2yP��셍3B�8��6ܲb�W3z��3\:�04��2������&�F3�5�5��5�U�evy6NM����(6�=��Q�A�2����n4�\�4��6��56*�6`�=6>�]�ۦ�6�f�5 E�5�𱶮��6Pg�;D�6��H��F���5�GB6�>5��s�f��³���*���6ժ1�t�E5�=i���l��*���p6 ��3j��5M��䴤47��#p��ǵA����{�PK*���D  D  PK                     < checkpoint/data/10FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���64*�����5��[7ƒ�܍)��ᡷ��� �*���-��.7Ё`���8u
������57"�(=���ڷ��.�x2�7���6���b5������.� ��6�娵���7��7��#6�7��v 5�05zy97��7ڨ���A7�b�JdI7��7�[\7�l�&
ö@�9��{7\l�7���7d�>7cSg7�BW���[7P� �3�0�5h��4A� f�4x���B�5����r�Z��6��7j�u6q(X7��	4�g|��7�#_��Q�6���d7�ʶ| 16��'��Kr7�U
�P����,����	7/������0+L6���7����M�7>���$�6�"h7ʵ����7�_�OE�J�6��7"ط����eD��S�7���6��3���v勺2[c7��N7 �ҵf�G��υ7Xj57��k�q��6-�۷̹�60�o���Զ���7p'G4�/��p�7+����~-v7.C�v��r�	8[��>h�7�{�7�.8�*+6l}�۰��te{6��|�j��7\��� �3��[5j����9�6h�
|�7��ȶ�KB�.Ff���Y6|l�N4d6��6�뇷^ ������K:�����:77X8�|��G6D����7�r17Ȁ8:څ6�7�7�+
5rC�Cn��މ�dL{6��57��97�"
68w����i7SLd7=ܶ�5��7$ځ6�E���c�J�ūS���%58���ݚ�\��  �l�@���6�%���6[컷^6S��A7����o�����ڌt�Ջ0756a7�"�5��8u�6��6�~27�ȷ�M��!A��\i7'�17&P\���ʶ��!8t!���L��rpp7D�7�l��<�79�^7Vh7�������7�E%���c��~�5N��6�ʓ7* 7�5P��c�����3!�7P�$64�~e.��!6��8�7ж�7<�#5R�6��.7Zg�N�{6��L��N 7������]72l�6�W���Jm6XK7(��6����d4�o9��Xu���S�5��?6 �W4�B�lG7 ��4O��<�7!a�5ʽ[7.�6Z��7ٔ7~��6�;E7V�7V��� Q��85'uv6H�����6Gҷ\έ� >��� 7���أ7��5Y��7�8��.	7��p��ℷ��.7��7��
5_[�
�7~*�5���6�a��6�Ҷ��1�ğ�5nB�6�b�tK	6^���|�y��5�7�K�
P����e���>�/	�6VŲ���6j�5���@u����e7��r��X�Ͷ�F�7:�y���	��@K��ܚ���q�2а���C6�4Ӷ����Ws6x(@6��7�f�XO7p����٨�rh�.N������\r�7d�Ӷ�ȷJ�������e� �k�t�07~�J6�$���)�����6@ �7��-6�n\7n-97@8��O���9�� C���^�7��8�f06l�W�4���s���~7Oj7 ��4 엵�v 7P��5�����Hֶ��7��N�xd	7'M�7(�6��6���6��7�$�6�Yn7��DQ�6`�4��G6�WE���74�q�m�����5,,6��޶��87q^D�h�k7n�p8N�8�c6��Ķ�G�5�mK7���6~]�7q��Lb�7<�5J���,8��	7
�77ـD6��z�Aζ��7�o�4t��7����k䈷�i�7H�ֵv�s1���u:7 ���䈶����6��7g�6#��7k⮷\dX7v_7x����6\�6T0O7�[68��7ӹ�7
�/��7t��ͽ75�7�� 8�c7��[7��7YfѶ��7���6�ͷ��1 8 �4���7Z��7�k�p�����ط��7|E������0'����7 �47�9t7��J648�'�6�
��P$���X77�P@8��5R�	��74P
�p����L�U��6�[���i!7��7t�,8*�<���O7`�u5.w�6:�"7(�N�*��7��صl��6@�4< ���S� �U�D�7�����B��I�7���7���7�:W���7�c<7�����52ݟ��׶���7��7u27��/�J�?��W��W���`3�6F�U6 � 60��O}	7״�7�3�6.y�7�ԇ�lk0���6����6>�27r/!8+չ5�7J��6�}m���6H�����G7��i5���7 ����̷X�*�����-N7bDO7v|�r�G������6}V˷��7z刷�7^7P74:�6Fc�{q緀��`?�j�`��Ѥ����a��+&�7`q��N�6c�7�a����d�����i��������.e.7s'���q5�h�7���¾��(�ǷA�v����s�¶8&>4�A϶��0�B�|��z`�H��� ��7�87�t8��
7k
7� 8(��6�+�6XZ57d;����5څo�?�p7���V۵L����L6dƶ5����6ՙ6F�÷���63̫� �+6PKW<љ�	  �	  PK                     < checkpoint/data/11FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ/6���5��w5��5��6\հ5�K76���5��65��%5Vֳ5�%)6%�5H$m5�9~5ϡ5�y�6Թ�58��5��#5���4)g55��5W�5ߛM5!�5
<�5Q�5���5��5���5��6#1�5��4_ח5��5
�s6��u5)!_5�OC5�qW5�1&6��%5�2�5E5�=15��#5.C$5a�B5P�t59�5 L5��@5�~�5	6(P5��5sp^5� 5�A+5؃�5��_6��_5�5nA5��5�`�5�V�4 5�m5TC�4#&b5>�5́@5��5���5�{�5h��5�s5O~�5r��5���5⎿5E2@5��5sO�5~�6 ��5�d85��h5�};5�^6�Z�5�5���5
�5`X5x�y5��S5�ߋ5�!�5k�5�:/5w��5u��5m�576��}5	�5NYD5� �5��'6�dq5lbd5��5Y�;5�V6{�5��~5ys�5q\�4w�c5�Ҡ5��5���5d�g6wT�5SE�5 �5z��5�;�5K�6��5�e�5�15HM�5���5�a�5��}5�]5��5	�76Җx5�z�5�؍5s�5��5in5"�4# *5J�76��5�d5�m45��}5��:5�/6�`�5%CF515k�5ɾ�5�̀5�Wf5�щ5S!w5��R6�+z5�s�5�5��4.e-5�i5�75?�5���5���5���5��5f� 6p�5\��5�c�5��G5�iI5�A�5t� 6�3z5�P5r��5�^D5�7B6��\5x�{5H7<5�Z�4D5eH05~)5��%5��6B\�5��5�]�5e�$6A,5PΚ5ɡ�5(�(5/95�1a5i�5��5e�5
?5��85��-6Zʋ5&��5QZf5��5�'5��5ID@5�Q&5UF�5нK5���5��5S�/6,�5�W�5(�5b5��4gYT5�6�؃5�D�5RQf5D�5a*6&g�5ov�5�A5�)
5�45��5^�_55F5-c�5㐟5`�O5i2�5H9
6�a�5}�#6ɵ5�t5� 5�7�5���5:��5��?5�,'5�0X5�5Q�5c
�5f�h5ֵ�4/u:5�)5�	W5sbn5���5�5RL5��N5�6���5�� 6��Q5�b�4�5�M5���5@��5+Y5��}5u(5�&6T,Y5��5D7.5|�5�y5zN!5"�4��5���5�Ư5��;5��5!u 6�B�5�M�5���5+z�4��E5�5�:6
�`5��X555�5PlG6��5�Q�5*3A5�>�42�85��,5595&E15���5abk5�&5'��5+�5��5=�5��}5��5BJ
5~�u5�+�5\	k5fOn5��4O�4p 6�a5�'5�#5[Y�4��[5w��4��5�F5̸�5B�5��-5<ɩ5��6�֢5��5��5��5Fa 5�}�5���5VU5�FN5�Oh5XS5ؕ*6�f5�D�5�O5	�
5­U5(�;52�75�H%5�*6��V5v��51U�5G�5�$�5��r6�0�5��>5��F5+*�5NK�5OK5�
�5)�J5C�J5�!S6�U�5�l�5�^\5� 	5�4z5gI:5��J5�vC5�Vu6���5%��5���5U6�J�5i�6p��5ÑW5'�`5�o6Z%�6?�d5��5Λ�5M��4���6�,Z5�U�5�j�5&.J5��5��5c�52|5	 �5���5��
5�^�5$� 6[s5ia 6��V5"�(5��55�,5إ�5�Qu5���5�5I�4Wk�5�D5��75�L5�H5<�$5^5�"�4��l5NB.6R=�5cYq5�/y56���5>x�5
�6�s5$��5nr�5�k�6>H�5�Ľ5��5��5��6���5U1�52A5Z�+5�Ȥ5:5SEi5��c5Ʀ�5�5�q55�R5���5�z�5�0�5�aD53P�4�	P5R��5�5�5�9x51%5�5n`5���5�B5��5Xzr5�5�M5�.&5Z�56�5V� 6�O�5�+i5[1�5؞�5Z �5�*�5�5�G5n5��5�*�5�5�P"5�B5��j5ڳ�5��Y5/"�5k��4M55�k5}oW5��*5~"L5$e#6݂x5�[O5���5+W�5E#�5�e�5�W�5�>5��\5%*�50C#6�w5�5�5Y5�j5r�6Bϓ5�5�5��4}JZ5�[5�oK5CD{5���5� 69t5o��5�0�5�w�5��5Y��5��N5�B;5bB�5��6�F�5X��5+�5ѽ`5f'6�Mv5�Y�5�]�5��H5RP5��5�45�tT5s��5���5@��5�5�z6� 67��5)w�55%5KaM5�X5���6	
�5�K�5��5r�5�y@6��D5"��5��P5p55v.5_G5s�5��5�y�5UW�5="5{^5@&�5�s5(Z�5Y��5-�	5��5�m�5�ӆ5 8�5�5�;5�i:5^�6��4�ZF5�"�5cO5
�!5�9%5�@J5?5PK�5���	  �	  PK                     < checkpoint/data/12FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/13FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ5z�7D~a���X�E�7��j7b��@)��97z�*� ��)�7߱�7g��7��]7.470��HN����θP��Sn6���7�ӱ�X7488�#�PK��˦d   d   PK                      checkpoint/data/14FB ZZZZZZZZZZZZZZZZZZZZZZZZR�6�6�d�60T�6�6��7Q��6*��6��6���6�/�6A�k6 9�6n�6���6aq	7m�n7U/�6-��6�.G6]1�6$��6�Dz6R"�6��{6PK��%kd   d   PK                      checkpoint/data/15FB ZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/16FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�����e6��7��2E��Ӛ�^��62$�58��6�5��֝��k3�å��)/���t6z�45��N� "C6B�4i6��{���γ��,��4����"���s�eۃ� �F+6Q�96xJ;6����p��I���0G4�i�5*3׵��r5�'��5�5u��T~�5�5r�L�ʵ�
5&c��޵���̪����&����4�7���W���5���6��+�ج�5�N�5hچ4H��������H��\6�op6��NDW���.�-�����4����`7�3:�D5��N���`εz��5F��6�Z�6��FO��`k6~6X���� �5��j��,ĵn@(6d�6
ζ P�6z��5 �� �7I�f60J_5˘�lE�6�ׯ��_O��9"����t ��\0�>��5�H�4)��4Ф���ҵwh_�a*H6j~�6�mc�B�4�3�O76fڊ��A�6�
�����4�|�e[6�Pݶ"��w���5�5<v��j�5	.6�L�5N�5�?��G��5�>��H����4\�6�Q�5�8L4)']�v�@��cG4�2��E�r���9���ֵd����k�4ަ���q51A�5JY68�7-�����u5pݴLg���g��ⶲ�50�*5R�6�/��lW�N��5<G�5��6@�*�>�5��4ڹ\�4�6H��6n,�5z1�1q�P�g�@-���6�7Z���Д6�Ʒ54	}��P'�xx�B���lL[�CB��@J5wb6 +�5�(��h�)�~F}�d����s6�N6x=<�J������6D�6p��5���5��D6�r95���4]ŵ�)�6DU��l�6�+g�Av��s������ h��^�`M �Isŵ�S46���5Vs 6�X�48�4��p5�6�/U�gc_6붯�X�4���4k�5����摵�Xl��a���S6��A4j�56|g6� �5ڿ��I
6&���J�R5ji6�u� ��30�6T�65 �����`�/�Պ��^굎ꁶ��6֋��v����)
�c��5��6���5��R�6�.&4GUV�R��-�zC����-�o45�l�5���� ��$��5��84�K�6+y�^���x�Ե��K6 X��OK����{5 �6�,V
�h?6z5�FP� �4<�6�%ǵ�{���]�JR�x���6��S5[`�<v@6Xd6
}��3�5y��p�4���1�|5Ը�5(#�����\A�XO��/������1��3��A�}6��#��赎s%6��6V+�5�Z�6�\�6/�D5�� �:P�f;ص�^T�8kc5ٓT������۽3�:K�X�V��6�X>�������5�뽵��5����a�60��m
��86(5<����6頊6��3Dp,5++��p�B��#��.�n6�]j5��4�ɍ4	*���Y_6L4�5��6Tm��f�5[	�5�<򵀯0���?�d��5d7|5^26�`�����5E���6Xgj51���V�5T�5t~�����5H�����5R�5�����5,d[�X����=m�����W�z6(��4��5 ��5L�����@6�06��6,�9��S�?�6�$6,!�5��õ�ԃ5 �0?��u�۵�t�6���5U92��)�m"X6��=5 ^��I
�5ޱ&6�(�\HZ��v� ""�yU䵔��6�ٲ��ꐶ���5�+[���G�6�m�"���|،������>��_8��
�y6��\5l䏴�r�HU��P<���ڵ��Ķ<��I�A65��5@�n3b{���J6$$�5\����C�5�Ƴ"U^5,����̲�� ��5tC�6q�4��26�n6
��$,26в9�H�<:#����44�������5�nx����5xn5���5��ڵ9��5�m6�w�!�4��6��S�4eܴ	q5�R5�5��8�5�;�4�$�R1A6i\6z�5ܪ7��Z���������m5�|$7��f4�V
����4J�d5��7zF�Z
�6܈4|&��⑨��#ɶ��O�(ɱ��3��]/�d-.7�^�6莙6�6n��6�I�6��?��~R5*��5��6�ƶ�gɷo���<l6�ӝ7�æ��76�Ԉ7s�t7_%7v�73;��ӎf7�N�7�}�z7�ǯ
�;��@�7����M�6�9�rv�6�6X�Ƕ"��6N�Ͷ{�L6b1���\7�h�5�`�6����bö�xy6�5�L6�����4F7b��5�6�7�S�p�qZD����6L�A��c�5U��5����$���17�v6�>���=� ��68�6�)�6Dr�5�&W��' 6�W��HOߵ֡���¶!� 5�m��J�6x
�JK�6��6ԑն����T�e6;��6n� ���4�E���@��|����:7g�ⶤ㖶������P��4�)��:�0���g5�')�H�5.��4�n7�I�5�]Ŷ�K2���5�����6�4��6�n	`��`��1���S�5Ә6A�Ƶ�4BK�5R�$����=�������_!�`�6e*׶(v���!?���ҵ�e�6A��5@��z�>�5�76%�6J����p��3���*�$�.G�5��6{&6�O���HgR��)7|Ax6?�A��{=6�w����P7�:��,J6|�6^R�6�]e���6�<�~�@6�*��"q7�5�6�HO�Ĭ�6�灶w#7.��6D�q��R�6��A6*� �g6)���̎J7�g��P�ٵbc�6�R7"��4�k(5���5cI�D��|���k�K50�6�	86LK��=r5�W���7mS��FK7�i#��[R�A���k���F	7���6�9��.74��5*��\>7O�/����50�u6�W�6G<�\���4�.�Ǵ��64}�`����?�n�6�מ6���6>�6e�+��۵�J6�Ȳ���6��ڶ�c��7$�b�0�)6*����q�K6l>n�7](6������6c��7�A��?j6�
 �
ȵڑV6���̿6�<����6���4i�6��r5��4���6l:;7�,��|9��|�6�,t��$�6@�n3x�Y���B�jY�6@�E6�T%���W�bQ7�W3�����?6���#7��6�S��@��5����$��'�L7.Ի�@�X6�C�I�6 ��6�#:5��8�0W6�6�d�����6P߬60xU4����g�5<e�5��M5�/7a�\�^�6`��3��1��0s;��![� =_���4&�=�컸�˜�$��K[%7�]�N!�6d�����6�:U6�k����26	���Q�\�׶3�c���\3粵 ��x2�6��'���ڵp'54ۦ�����r�K�#6g��6 I�л��6&�'��D����6/����}���y��bu6�$�z�L6
N:�����7��նr�E�cXC��D�6�F�M��߶�~�6O:��kǩ�6��5��C�����<Z���˯����6^��4*���B1�;�6l�y6�U�6��v����U,U����6�ж@u�4�S�6��׵3d
6�=�t����ŶC�7r7�q�5:�E�x�ŵ R����|6ƨ6�����5�Ҵ�Wx6*г�Ě�6��״�հ��>�5)���P�6�1���D[6��t6�>5��*�J7��W6��6"����6�p��i۶��7�A�4-9�5��N�J#T�ޭX6!��wضw�x6(�p� �����6���da����6��&7��-6BN����v�c6���4��6���4�L�6���U��5	 �HT�M����!X7�����P[�i*�<��5�J7u���=D�6�6�6�vk����6�6�����9ҵ��ݴL�b6�`�6���sڗ��G���G��z�C�>v��f�6���6@m\5���6�b��~yE��#���j���4��^��|��5���3�4Ķ���6�XN� #ʶ��ֶ���y5`F�4����繶��h�2����<���ٶ���B�a7����F6��6΅����5PC�4�J?�P�ܥ�.q7H�Ե�W��^6XvK7�|�7ސ�6p�4�$�F�)70:�3W�L�Ha��`��a �6��6�?v���y�60ˁ�/�Ҷ�37ӝV� =4��7��l��|�ƕѶ�Kٵ�W�}��6ӏ6ֺ�6�?;�lf�
�%��d�7���6ފ���6�g�6���_��6Q2�6�h�e
7M�'5��׶~�]�آ7!x���i7�M6f���^7La�T�'56\N���60p6΍���x'7���5E�6�7�	�.O�5��7����Īo�L7������278�6֢�6j��$ȵ�m7Z@�7�wL4b�O60u��¹B�(�7���w�� ����
�4`ӧ�8A6~<77����5U𝶂ݮ6SK6xq6�g���	7��'��G��
'70)6t�
6ۙ�6@��6��50]���9j7ep'6 �ʴ����x���gs���X:��z�64]�6��ƶU'�6�2�Y�PJ��.���9�,����ℵ	�X���Z�L�����5�v%5�4!��*L��iO5f}���ζT�R�3=�6��7^��6n��5�#ݵd�쵠����ֻ������¹�;����6�_e�L����������6�ց7�iö��5�Ѩ6R0��A��yw���	�� ���b���|�6b����qٶvl�6�����6j�>7�%���6��ʶ��v�N���\�6 %ֳ<T��$��^}�=�U ��-��J� 6���5��m7}���4ε(��	v9�lLյX7+Q���57627�K�6�WJ�R��0
���7�6�P6���1�d!m6�P66��޵���4��53_��m"�7�}7����r\6kT˵�R7�"��j7k��6����z~5<��6�ȅ�ɞ����6���|iM6o�5�iA6��55�ٶ��574�z�@�W6(&��b�6l��6n�ʵ�Lv6Ŭ ������m�5 ��4���68�i��RE68G7.�=5:�6��+(�6���5��56[fB�_,����4�䵀���x���:�6
T�64�����H�v5,�7vk6����@�ĳ0��ܵd7�6d66�dF5�52�6'��b�(�G5��6�L�tp�6tf86��5`˶df6��6��m6�l�6�7`6���5X��0�4���5n5�$5!��5fj�l���.e�܍�6�H�������K���6|���j�5���5��k� �e6d5�~g�%�õdM�5P�3��m6M^n6��!���b�ǵ/����y�5�>)��f6�N���3��5ױG�R�N60f{6�X���!5�Z����V*-6�g���?5؏��h'ƵL�~�dlS5H�"���v6غ[6��d����:�<���D����w06�B������B$�"�C� �5����6ݳ���Z��T��4�G}����5�~f6�ĶX�5��^5$���H�66B�J6�魳h��6��J6Zĵ#$�[uP��T�6��6J��5xT�5���h/i6Xǹ� yA�%��6rg$�?S"6\�k��s5�3m^6�84��)��;�6��$����6�%b���6�3�6��6�5ܶ0e��ױ��*�5:���M37�-���}C�LW-544"�����I7�����6Y�6�*���6dH��@3�6�B�6hLǴHϵ&[�6���6�Eյ}�X�������58���J8��*q�������+d��F�62_���N�69�ᵅ�p�씟�P�A���v�����)7<ʓ5qN�5���5�n�5�'��(3�5b0�6إ�w(6p�4������4ɴ�j[;� �w�|HƶlA�Ⱥ(���"7{��5@<�5��,60�I�����@��4��J�Z�ŵI�%�r1g����o����ŶK�5�y6 �̲l�A6(Ȗ�	W\�[ڶ���6H[6�յr "5?�E���$������|ʶQ�7pw�l�Ŷ;����u6g���W���6�*��m���/I6��p���5��[���9s6�D$�УD�2��6jf!6�H��,K7���*sO� ��4l�}��� �i4���6:�R6 <�6�tZ�3�'6��%���%�4M�j��Q��nV�6ߴ6F����s�L7��}6Ƃ�6b��6D����7(�p�Te����6��^60�Ҷ>T6�1d6��鴀�(4��5��3�	s�6�Ѷ�4���[6��^��S�6�I 7u2�6�����9��&7���6�/출[F�M�A��'6S��6"s��EM�6^�62�I�~}�6��6�]���󶆅�5�]6�#������ֶ�_ܶ�A���+��Iܟ6����6�I76Rɷ`�#��Q����3�@Zf���]6V�3ʱ�6{V�6�5a�tm��tY>��M	�݆S��1k4p21��P6��W��w�
6�6��۶�߶JN�6l�	6M�(P�88� x����S�h��Ԩ��$��?��Ĝ�5�k�6(x�5�悶���5j��6t�6Ly��w����ֽ߶��`%���³&�6@�6 ��2B/��?m���G!7���4����v�5�%ҵ��6��5�D{w6�C7���6t�4ׅݶ�[7���6`�A 6hՉ�.�)7���5�B�5h�G�1��;Ƕ�>g6������k�^T7��5���l� ��7�"��0|���C6�糶�@D6�Y��"�3�⳶(�6
�;���~6Z��6���������L�P��������ն�G��x�5� ԶF17�(�6�<���v6�d0�8�¶P<�J����@�6���5:�66��#$5>l�^��>?޶pa`6�C5��6S��6��t6��u6��붐L˵=q�6�-���6�ᇶ܆}��W�5Dy�5U��5�a�5�s�5��A�h��3K�h��$$@!5���rX5]F�lt5J{��d�5���5�ᴟ*�6�ܴɰ,��`3 F4��Ƒ�Ɲ����>6t�z������6�ND6���64��9W5~g7d���y"��x����5��|ߑ5�X���(�5І6���5�H��E��|PĶ)��6���5��I6�?��ԫ4���&5AdI6��)�D%75�G6anC�hu*��6��5 ���J�嶛EU6���$�C��Z����6&��6P%�4<�ʶގŶ!��5$�6�~���Љ4��f5��k4$�I5ð�����h�\���ŶV���a0�6rY85(�ܶdi5�ߖ����5��5��16�2�55�6v̶�������bSr6��(4&�b��4-7qE68W6�wz�kY�V��5�	��k�6ʔ�6(r�`�e�	��6��M�P����s�f�E���6��25�z�A�6@�4$)��y���Vw��#�ռx6 f�3uψ5�J*6�"{�%�Ҷ�S6���=�,΋��/-�	M�6�o�y��6$:Y��'�6F�!6\Ю�q��#5�l5�@�W6lOz�^3Q6����16za	6@p�4P�5L��������6�ѹ6�h6$��L��s7 �K��T��蓮�Ɇ϶�(���K�����4j�F4�2�5����6)6�4C�6@��sz6���6/["��2�6%���96�.�6lW��p����|!�����r�5���6}6����N�E|6��ⵈ+)�ɜ�6�j���w36+k�1����6N���6��X���~6��H���޵��γ ��6ƶBk�̯����A�׶8��5�Z��Pߴ+���7��V��4�� y6�@6NcS6�i��}�5��}��?!�4�_5�Q���գ5+��e椶��.6�6�x6<O�6ĝV��}�4vݗ6��a�4�M5 01w};5�Dl6L�� \6�-��.$5H��42"{69�8�H,_6�(�g)�6u\��>�E��1J6�\�6K��5��&���z6�@?5��5̯K6�׵kn�60��v(��r��6�7��5���5�!��Jb6�����5T�6�W�؊�5r�6|�[4�4NT���\�����6X|5����*�6u�5> 6��|�D��}D�,D=5�8q4[��l���C�2�~�3��(�5�Zh4�{e�}C��墆6Z0�m�=67(��[��+�6X!ӳX��4x�G5���4`�6�o6�U�>j�4e���&��uT 5 �6l
�j85^ 	�u�*�|�E;���T�6+X´���5|[�ނ6A 6r��6;b��6��"`U��A5}��$�|5 p�Þ��[&�6����6�F�j�7�k�4��6D?�]����5�s�5��5dS6k�9�@hN3Xt�5��"�Zy�5�OA5��B��,5�k����66�6||*6��r60w���6R+���7�v6�'w��O�6�D�5޳�����4�M5'p6�5��0�FA:6Wx��K��6�öd�Y5L�3���U5�µ/�Ƕ���*)��S� 6�Ob��4����M��%�$ML����4=M�6u	���e�cL6?��0�ֵ�����g9��&��蕉�#�5�X�{�("x�S���J��f�C6 (�(o�4$�I5N})���4r�I����6
�(���˵��Y6Y������&��2�5?��6�>��SJ��|=6_;^6��T6��˶#�6PVb�kyx��"�f�5\R�G��6!�5�^��h������6�26�l#3�`�5�/.��"�ʫ�4ҥ6��|6�Ŷ�Q�6w�е*N��L��6 �;�͵�	�5�oe6%d�d.�4�5�>a6��$5�X�5d	�5��5M��56�1�cx5��*6{(5���5x�a6��Ķ�A�5�óh�h69�Q��.�4�u�xC˶�0�6Ԡ,5�Id�}�7d���ƺ5��M6�#��oO56���3,�~�/:6��d� �t5���62�5��!6�6"�0�2~/4͖��*c6��I��X��j���5��V5�ib���F�j�|69��6%��zg�6gJ���f6 5��,�4��T�xҧ3%+5��6Bv���5���5��_�H[�ը���5��R5���q��5�B�6�X451��X��55e�4��-�g��\�ö�,K��[�6b&�L�5���s:h64� 6��O6s`d5�
r6ոr6�$�r6��gYB6�L�n�q6$M)6;�5R�>6�����4��6��޳�H6p�51$�5���w�)6�O�Z~
��@6X�;4��6���6 �e5���5JY�����61����6倉�Rݵ8��E�5#�7����:����4�;5B�I��d���b���5�F?�$\&6���5{��-B6��6����ս��)�!F����-58�6�7#�gH6щ�6���5Ъ���x6-P�4��4��6���5m�5^뢶��5�sS6�$�h�x5WDҵz��55{�ᾚ�ikS�Ѭ&���6�f�ރ�����6EE&���е�6Lh�430����B6�3I��k�5�X��5���X
6����]��6܀^�KJ��c6��c4�]��������rj�t<�6j(?�Kރ���'6�f���Oc�x4����5묋6�"�̗G��r��:��:� 6:���%d�5n#����tkĴYa6�>�6q�ε X6�����lܴ��k6�n$��5��1�[n�6�	\�8w+���?�@�E5ך��@��6��@�񞏶4P��x�����4L~��d[+6�R�5ٴ��/�r5.�ǵj�16 ]T5�6;�P6�/<���w5$ܴ5\�k��_��e����]q��G	������^�5x ��sZ�*�#���_���4���5� F5e�� �ͱ��_�����qs5R̵q&��55�[E��EG�����P��R56SZ�UJ*���5V`5�f15s�6ӫ�
��,IǶJ맶.J�6�7��Y+k��{�xɳ�RܵӞ涔su����5���4������I%6pJL5V���k����5ɰ)�����B�6�#l�◞6EMT��J�5^%�6X��������a��˵�G�P^5Z���4";5���6�:���6�5�B�5U^ŵG��6���6Xñ�D//6��C3hN�+�5���xc5���6��5���5�ҵ�D*6D_���6*A@��[�4���6���6`x´}o�6,=5Y#�6v�(�D���^\� .�1<�m5@&�D�µe�6Xn-6 ��0��B%?��uS4\�鶓c���1��(�6���5�d����/ұ����6�ts�t!�5��6�9z����T.��G6fʫ5���4$ː���A6����������62~R��@���g���66Ԕ6��6�h6xد5H�v�3,�5�,Ӷ�
|4+{6)�3���5T>7��۵���5LF�5Pڽ�$r�5��D�5!r@�0���N������J�5��t�b��5W�>6�/]5�CY�ʰ�5̹P�\x������R�T`�5�6�~�5���5�Iv���J��3]7��50ᑴ��~����4��x5$Yk6��������0j� ��)�Fy��hϵ�r-6
��6���+!<5,�4��Z6+5�PЮ��78���������J�J�6��>5�V��@e6M=µP�Y4�S�6�5ɥݶ��I��������oZ����5J�P6 �4Th�����0$�5�?�풶�5���|��0��.T����ҵV��4h��5�Z"6�6P���ڵHHT��µPյ�R���g��耒��5�7ƶ	�6u�26<o�W��d/r�8K����6����p���n�P6��6�6�FP�ZT�6�`7����h�W4$D�5f�6��'6�{��$�����S��(�54̈5��Y6�9�5�u�6Lu7d6Ó��0��4�F��������5'n���26)�5��
����X$�����5EUB6�s���6���z496bXR57P��]r6��k��Kw5��76Gŋ�Ee�6&i6�Z����	�=B6$'V5��<���5re��*6�z�5R�S��r��D����C��h�����6����/6Q��4�4�;6��q6��µ>:q6*X�.5~5�j_6+�鵪�.��◵z��6U�u��:��Fp�6��55+.���d5l�M������5�2��}��6��<��_�68v5�����I� 6��5G�H6���V�6e�5jL6RE��Ji���ɵ��<6V�Y5ȅN5�������y5]����X�5��N5��X6pj#�Ӆ�|U5cf�5�F�4$��Y�6���1t�4���4�Q 6�h!6�q=�Ex��J�/6	[�5tR�����2��'�s�!�ʧ�~�񵹾e�Yz�6N��^@5Mj6`c�И��C�56j,�x,��2M@68�������	6�[5`�?J<4��6'�A6�����5گ۵���58"�6'㪵��ߴ�k�4�qo6�L5D`�5����5�N6�IA�y���#�	6���6 ?"5�������� �5N�5�s�P6�T���ș�r-�糝6zЍ5�?�5��a6�*l�<xc6rä��O6zEp�Ц!6��H�4�;���d6�恶K�5&��5��6"��g�%6����ߣ�����6�[M6��ص���6Ʌ3��=鵔�´�n�����$���677[6��ʵ��
X|5b�E6B���j�h5��4�DO6�k�*Ѣ6ʻ �b��5�Κ�0@*�q�k5]uC5���B1߶t	6V��8�6��3�F��va6�9�6�������p�N9
�,!�4J�N�R�˴_vz�zS�5w,W5�r\4�D��p��5��8��C��l�5��6˶�5ܗ\��;�53�68E���36�
�M�;5�~�5&5���5��T5y�)��0"6����p� ��v��)�(���5sV�5h��H��5�Z� Mw4� �5 �m��Lȶ�DZ����l��̮~5���6�x6ٴ6�`��t��ٶ@m���6"ă�{/�6Z�66���6%�6��#����=>�6�O�5Ȭ@5�Rw�5�ʶ�[���i5�5�P�� UO�<��6�͊6~�ڵ�s���@ص �5�2��<m6{h����5Bg���'���6����O�\b~�XAE���6� ��T�����l6cD(����5X�5 ��V=-6�B�5f�B��/�6����$6�w����M��/5?�-6���Z��5t��5R`ɶ�'�w6��6p�#5�6[ϵ�l�5�����r?6}q�_�4|�6��
�r�����6�vN���6�6�46�C�5�9�pt52O5aa5d|��ҥ��@�����62��]]�6��5kQ�6k�5��6��%���5 ��3U��/�7 .�4���4�	����5�÷6p��5�b5�/�5 6󦻶�����5��5T~ʵ�1���̴�ٶ�Q6ol�Ju�6�Ag6@b��E��6�D6�;��wLb6��9�����6k=��Ǫ����5i=R6 �4PK5���6��5�ߵ�W_�4��_7l��)̌6��Z6�����B�3.�6��z5��;6b���h�6��76�C��"��54�t5-P)6�76\;!5P������zj�50_�4h��5���6o�����"�b䙵�C�4�	9����5Kv��!o���/6��5@'v�sS6�K�4�d�6�V���׬6e��6�n����6)��4SF�6�ܶ �L6��b�h����!6Aq�6|x�5�)6���V﵄s����0�9⧵�26�y�5T��z�6b5��6p��6�����@�6L
͵�T*6������6 �n5��"���5�۵�v�6�{׵�N56$�;�=6��6������5UW�6 �ǵJ��6���6��a65K1�5  6�M�5��6N-6�2	�gw��Sx6�~�6�=68"5���5�,q5�oŴDk�6�﮵\9�5�t�4�B6X�4��5
Ɯ��jݴh�'�d�6\���M_��Z􎶨�6{/6N�5�V�-6Q� �ԎеmƦ6'|u� �{�LE�6ĭ#6����r^�6 i|4��[66�5@�~�o�ε(��60[���J�k����#�1�6X��$���,�0�5Dl�5�E���ܵC�6��Z�y�+���3��5E*�5ϛ`�>!���]��HR�?��
t�5�|7)ϵ�4���M��Q.���i&6J���V��J6���{�����63�E6:l�Z������6>rY~��є5��6���ε��=6�����Jv��r�5�a¶^��6��#5��6=��0�c4��6:�
6��6�)5�9�6�4\��ƌ��ѓ6qN�57��6�6� �4h�6Z�5ݖõZ��5|,v����������16���4��6>��5�8N��Չ�i6v7��ב�[ �5x�6P{���6]�B�8�f6��5藓6�-��"�r�|��5ʀ�6�v�Ӈ�5،v6:��,�p�h�f�Dg6�4'6��6��ݵ7��Yh6�����5PX�3"��5KV�5��^�Y5����~��H5V�=�B��56�A6j�W�ok6p#���`�6$h����ɶ�+��P�Y6�h�6&�D�Ȕ����#1�4�2��V�\�o6x�R��!ʳ +���iU5�a�d$���6Nu�� � �`��6�IW6��5V.X6PW���S>4�%6}^�5��6�K���"7%$6p��56�6D�e5�9˶��69�5����5�"7O_�5T�6dR�6@�ȳ�>i�߉6dt"��?��AԴ�_6��;67�6��o6�ᶴ�Ū3 6C6x���D��o��	%�Β6 r02���6��ᶶ����2�T6��
s�5W{��J��e��.�6�����6%~�6�c5�3���!���l6��78�;5?�|6�N����x�z�Ƕ�478��6���t��6����4��7��C��m|5�Y�6���6a�5n�ж0�6�T�59���;7E8��996��4�����
6�O6T�յՋb6�#ζt��6���6rG�6 t����ֶ�q��Td6�M���6p��5T��5Q�_����5����%��6.�B6DH�6�h�ȩ�z� 6��8�:�5$?��ؐ�d�����6����~ڪ����6Wɐ���7�:f�5��D3BH�6�R4�@���6^-$�� 6�B^7�:6����YǶ�;�6�?6��Y�����44�V5�Ü�ӷ�5��6���5�@��?�6ȟZ6f=p6�k5�S��O��в�5wq�5����Ԥ���F��u/�~�6�y�6�Y�2(6��Զ�Wp6��F6�1j�JE��7p���z�:��؀��M����5��7J��4���mA�4��_�E�6��� ��3�5(7��������6˜���j6Z�w�t�(�ue[6\�o5�B�6(��6ik�]r�62����d��?�h�y޶����e�7�E�z���6��3�`�[6�R07�ޖ�����G�5y�$��R�-�N�Ŷ��� �Y�{G��[��W��H�60��4��~Y�6�"�4��;sv6��W��D
6�ڗ5`?1�T?����6pr����ǵ������7`J��a<6�w 7ڍ'�]ʶ^��R�6!�X��Գ5ﵧ�+7�	����5���
૶2�U5 �p5���.̶�-s�2(d6m��6ҿ���)7�����5l���c�6��p&7lO5<�!�̵��嶹P����5�D\6&��6�1��I�'��柶 &/���o6�"]��'�6K�~;)���6�h����5�h����,6�M/�bjݵ+i�3�b�4�_"63%����6�ա6`������3�+�)8�4!M�D�"��<J��x:���}��6�i�2Z��ߛ$6��6��6l�3�F�~�����(9����� �\���L6N�26��p(����� �I2<p���������h^�5�P5n�5�����H��93 T�d���V���e5�:6�j;�J�6�����V��K¶�!�������f���&��-��F5��Ύ�5�F>��L�6~�U��̻�ܡ��8�7���-5^���F���8$@64=3��^y4H�/��5
�@5�Ij6 ���-c6��(� �W��LR62�.�tԼ4�i��F�6Tq5��s˵7	�?o���1�5^��5dn74��.*�5��[����6<�5�l4\���d6�X-�T��6ԛ'���З05��ڶB �X{_�PV�5���5�C6�<��S�5H�s���?63�����5F:����5���6���3U�?6�㫶���5`m����76Pr$6P�A5��5�96�P6�.B5���4�[�4B�=4sW��p:l�b\�5�]6���m	6�>v�x(6赀l3�V����5(�贖�6��)���{�����П�4��6�� 5��ٵ�5����9��J2شܦ�4��46�/�(A}��.���L56~���`��6V~�6`k6֝O6����`{6�x/�(�6O�\��5��@422µ
�5p�5����ݴ�e6���6���6*�I5`ꂵ�+56a�o6�յ��.�w>��c76�ٵE���md	6կ�6<=����&�T8��6�/�5�m2���"��55�H����:���50`X4 k�4?�ŵ ����5��5uv�5"[f5:A�5�߯5�:'�"��6H[�5��s�P�'�C�&6R�������^�6�"��~�5 E��e;�946�s6�뵞��6��]���]��ڈ�	=�5 "�5ޓδ�C�6�O�5|��4f�4 �g�\e6 �3`(6��~��l��S5��,�&�?����5��85 ��4���E\�ww5�(�@.�2������u!��a���96�?75��4":6���6Q�66�&����|H6b�����6Bʵ��´���6���4�=6=�6��;�1�58'���F�5dy¶��T��$q��z�6:p6_V{5��'6mQ϶����6�[�6�q6�!�7��'��p��D!6�_��6�qw6c�����u�5���^�6t�94��$6 ��4�5J����N��~ϳ϶�4��3��ಡ��6����ze��L �4G{�5��7��,����/���Զu�5�˵>A66��7w��������z6K�
��~����a4di��g6���5���5��6�5����D�����Ķf�^�>Ro�@a4h��5B�����x6���C4��6����l�5�.��5��6�4�)��5\���rx5�16����	�6}8��}I��qa6 ^#6X�����6��:�^�3521�6q��"5��/5/O��a:����Td��c�6Ȧ^3���4�����6�f���A���6n�Y�(�ض�
�6�|d6���6�x�5n�5�)��B6�S��{�a3��ߵ��5���6�O�5e�0�,_5{A�6�}86�7B7Ş�5Dp������@��~*�����4\�6gX6�i��e�6|䨵��,6.O�X��4��26Y�t6�Җ�(F�5��N6��5-,6��.6�8�z��������-��r*6���4���P^�5��4�j6j5$��5��8��	�����
n�����5�p�3a�t��DH6�>q6G�iy6zL�6N��6<�5��=� Ot���:6�+;7�/�6��l�6)�e6"ͶpC�4���4�	��mJ7PZ�5־�5�l�6 �)�J���!B�6������@Gt6xj��e�6��|3��O69_26L�a��Y�6$]���04>�"�Ft��LB60�o4�y�4Y���~5�<�5H:6�3`�@�6J��4�`�<�6�޲4����,`,7�t�5��m6��5� C�~��6/�6�)���O�����Ԃ�6�t̵T�&��t�3 �94�u%���=��Pݶc72��EG�N h�5,��^F��!\��浰X6�d6B�*�/�F6�p6��h6����I}&�X�65� 
�`���ȵ��G�X�b��N[5�cY��t� ���϶5�|�ٌ�
6�)�6@ �F�d�.��5��6��P�!4ꗮ�/沴�047�}D�2�n5��ε�!]6�S5���5J��6�8H��j�6��4�}j�m��5��5�&�4�[�6�A86����.��"�5�816�r���,v6&;6��J���.�L6��#6 �j4"��⵶L��6��7* 6��1��v6(s]6H��3 S�3L��#�Y���5�H5�M�6+����A�M���5�<�v���9ڶ�r54�W���%��` 6Dե5��}4�86p�4�� �G6�撵��*5'��6�ѯ�Pml����6ִ#6~|��0^���`��I����P�6���5����n�6�fi6W~`�_�޶��6@xV5D�us�9u����6@��4��BH�6�ം3�5��6v��4���H�4���6��B4&[>6�m��wp����5��%��"�6Gd�����&��6�.6�߶͌�]�>�R��5�Ǘ6��������5`6�}���9;6�_5k��6������ܶ�b_6�*M4 �� �m5��n6�����iT��9:5}��6(Fĳw��6��е���,��6��6z�}�+n+����6�t��FI��ȶ��B6�}6l��6(�p4�PH����45�#���
4��$5c�#6L��4�Ȓ�JĆ�봶`����"�Skg5(`�3�nԶ��R6��6ƾ{�H0¶	��5��� -a��И5.���f��5��6��Ǵ��],���?�5��H��p�"�5I96 ���`׆���O��dY����54#�5��5��5<w��h�5��6��5�7�_6(;���P���^!6Py5��ص���X����6jPζJ����8�6愅6�e�6A�6L�ᶸ`(7)$9���c��s\�P�0��U�蝮5|������������#�	K�5�a7J�,7�DW5VDǶ��	�߄�6�K���<���z��ضd䋷1�6���9���c;���D1m�W��6����ٵp�O��6j��n����D6�05��V4��_6H�6��N��6`���Oϳ�'�.7�v.6,2�58���DŶ]�]6�ZD64J�����F��6����B������B@S���6ϯ�7���4��6w���a��5"�ඍ�86`�55��l�������ᶼa��#g���g�69~�6�N�5��z6L%5م!��0���^�6-}e�T��6A�����6��6+�}6�ϼ6$)��f'6�Y�����6�̟5�Ӧ5X�{7@˴jj��7r4>70D�I�	7�s����*.�~#6�5�6eȜ��ĵvz ��|�6*im����l4�5ZKɵ�6��5��,��q6�zŵ{Z� .5 {���YF5��7���5�~ 5*���6B��5r4h�[9���5K��F�6�����ǵ��趄	7)��5�+C�K�Y�7��5��j���5��X�g�6@Ȃ6R���	뵌���u�6���6uΘ�L���w�5쾥��鴞N�5�"d6�ٙ��S�6bdB6̶��p}�6+��8���v�5烵�-��w16�w���}����7�D��6�����/5�6���@�M��K��-?�F�F���T6 ���no7j=B6��<��,�*� �f����_�����e�3;g�����Ŷ;EX6�"� i*��ai6���6��7j�6���5�5x�k5����/�96/�������6`����6�L	���Z��� �U�#�T.I5>{k�lw06���r6�Ρ6\�ص�N�4�i[���'4P$�5W����q3������������u��֊��-�6�~�5K�D6]}7N��5���r��6�6ճ��6��[�$K��ܦ6ǲ+�l@(7|��5��]5Sy6j�B����6���6�� ���#������ж	E6.���5^Q6�25�E�6�*�5��6r����v����6D˿6y�p7 ���v[Ѷ^����c��4J�쏃����6D�*6�f��uŞ6��b�$�D6��3f�626���h!�6��b�Nv6�&6�?�b���\6��6�KH6�����4$r�5�(��h�1��1����6�(�6�s�6>�6Œ����
��5ް_5�Hf�n/-�C�6%R>6pW��=�۶�5���5Z��5��Y���h6N�6(>�5��6��0�̱�e��6�r{5����C�8g�6{�6�������5� ��	�}�����/63˴6U�1�7��5*D� �o6�~H����6�$�6S�6Xg�ö�=m5���6(��6А@��յm�<1�z6��i��:���'ζ؆��6�uE4�6Ԃ�6ԙz��H��J��Ϝ6�75�1��n�6�b�S��6��t5 u�rV5$����5�,#6��V��v"6�ڥ2��޶䕆�_V6���6�ƶ1G��Ȁ�6v�z68�3�:�5<m�6�����]a�Te�5�@o5z���6Gᶄ��55��6X�"�'5�cc7g46�n𶷗l�WW3�>Sk6��*�[z�7�������6�V�4_�᯷6�h������i�6$��6���z66tX��܏�6�l�5	*76�I��Q	7���X�.��L�6g��5~�I7�v���X7u�����E7��26���6�>O�C^�6$5��5�6D�7�%o��$���zﶖ�6$Y����/��7��-7�t6o� 7<X�@%��$
��ɵ���5������6��*�k����6`��5U�L6���~������b��4�6O�[5���|�6+�In26%�36�����6ѵö�6�
�6l�������TJ��60Ki��;	���6��5`&��|�� �6��(�ݵ���J�54�񵎻R5��r6�Oo���n�x�5�J�'f�*F6X��	R������x�60��6&��6�q��,G�5B6P��5���5 K$24��5�s�A6�<���M����6ǵM��5��-64^ݶ�oo6fɴ��=S6 ��3�6I���q5@�ݴ�N_���6ޖ��y9϶��[5{C�6�5�����:��?�4V��2�:ע5���`��6)f6Y�6�5�w4���6���4w��
5���)���6���Gb6�J�6������L�#�7{�8�$��5����6�Hw�x{�4$޵��v6�n6��6�7��N5�T%6�e[5���G��6�c6��r�L#6������㰵��
6�ל6�D�4b�����5�5P*�69�4�f,6Sɵ��,5/:����6鶺6X7L5�fⵯ�ٶ�� ��b��id9���6��������4µ�4:�6H����\��~�b6TJ�����6�W�58+�4�z	7,/ߵ�!�5v;M��q�6��]�d�5/����;�잼5(r��fK55#��5Fv;6������j�ڒ�6�Z�s+_��@�6��K6Nf��ͽR6N��4��M6��Z5oO6Tn�5�"7g悶k��5 ���4{��,�V���*4(����6�Pi5�J�����6h#l��[�5��6��Z��3$�R	��O�g6X�L6"�M5��6�ܡ6��b��/b�֋ѵ��5�̼6���&꘵�㍵h�6��εЇ��o�쵒bе~6��A\7!�6O6�.6m��6�_%7�:9������F6z�56Ȅ
6��/6Mg��j`A6&$6 ~2�_�(nֵji#6��t�~�ȶ�a�6L�M6�25fE(�JQζ�	K�Jնy��6õ�6Hݹ�H77ƨ��30�6�Y���|�6Η6�/�6�-��J_�6ް�6�6@o6ȥ��f���>䶖��6Z]6��q5AO6b�6��R���#6�Y�5"�	�ѩ�5vP�5��5�W�4�-Y���#��b9��ʄ��E6�)U���k��$%�����l
��M	���5i�7n#�6�冶���77����P477�j��K��6̍6��6�-��x��_}��Ø6$�6F��5F;46�(��U��^R�6��)��+7|Z{�ܫ���.��|�X5,�o�H{#�G�6ԇ���6��k��Q�����~27e�5�G
6Rj����26Η�5��B�	���m7�%�6q��5�sS�`7R�^��6�u���e6$�h5w�/�ଶ� p�]T�����5��6G����Dn6�eӵ�g����6��6�,�����aP���0�2%6<zɶ c�4zr7�=6 ��64���Z����L07 y�6t5� (�3�N�6���6t�y�r�Z�6���4�mQ���I6��7�N��q��6�
/6 ⑴I�5R<��	6%�5�~5�Y�6K;� ����f����6��3��V�6�ţ5 s��<+7X�6t@x�z�Y�b86�ME�岵5�㶰����Y*�i��5{��ƕ�`��6��6��6��>���;5����8nE����7�xj6���}m)6a�"72����g�6�+7ڸ��g�K��$>6�.��Zt��Z7<Pt7�ۙ6nv��HFu��lնVM)7�Gֶ�6Ɖ5�'��$�6�í6�_�8J�5 i�4�6$�dX%5����d��6 ��4 ���?�v��Ԏ�8E��� 6��5q�6��6P�� w�e�̶AB���~�v��6��5�cj�hL%�<j��Cu7�J�P�`4�B7��>�D�c���\�3�+��>�N6��%����5`�	4W��6ϨJ5`������s�5���5�(7$7��|95�*��N<�6i�6�6�h64������.36.�߶���6�5HW5>�O7\���F��6!ɵ���J�6#(g5x"�4�{ϵ��� 1��̪5 Rm2@66�w�5���5 �?1=�l6T086�V�ozS6��)��I6�&¶��#�d?06�v56�r96��6��������j5�0`�6�B��K��5��A5<|1��:F6%i�������� �J6UG���x���5`6P5�華���3�����7��X6����M����"�6�3��hk�5���;W���e6�e��b��h[_���õV�86���`v�5b��5���4��2Z���D���G5���5jTr�������>�5� �,��U"f�|�t�$��4����4�е��Ua6����Uq���6p7<5��_��	6H�8�QQ�5��6���Mw5�u4�L��������f�|1�5z�a4��6왳5W��6�d�5�(��!�4� ���5��j5;ʗ5�=C5�C5�#�5�i��R4�M�5Do0�o�u6`J6�B6t��`+ʴ�5`��6r���錶R4b���y��9j��Z� �N4I6D�Դ0b�4��w�"�R��6��%���[5�*�5Ù��P�5��6������5����;�3���������t��+�5(%Z�(�i4�s6��.���5X�������r�%�))5�፶��6��޵%�޵V�ݵX�d��ڬ4��N�&6� B��5hѡ4E6'�5~��#޳%{��jh,5��T&ӵD��5�h鵘~����?6#��5]m�6�b6�d^4��v�>�c�6��U6�s�5�)���;�I�3�
6���5��6�v*�����L�v�X��4s��� 즴�w�P5��F����6�Vi�m�� B�k���5�]6�C��d��w36x�/5�z6.=�5��5�֙4|�5�
��w�����t��P��^ȅ�`�5: յ�N����{6�ng5$ް4���^�6��Ե]��5H\��S���B/6�5��	��.�\�}5��4��q6@�� ��͑��%��y���5�|���&.�,� ��h�5���5#����si6����ʹ������끶6�&6Su��'����6 �v1Ǆs6��q����6>��2r�h����&��ȗ6,�n��~m6T�X6s5��%���[5�{���0��\5�õ&�6��5M���)�69Ku6�����5<�ն�L�$lµ�)5��5&p�5�p�5>m���� 6&�6�b`�����&x�|����60򱵖��5c�6��3��[6ME�b��ر�4X}`�E��5<��5J�F��Ҭ�D��l16lW��k�5���5S�F�+���@�̲p��6 5H���6q8�ª�$;��4�����0�6�[ҵ��4*K��w����5Ą6l�5��R���5�JܳTM6_�5���m�5�����-�6��Ŵ�n6`U�4,6?)��|�p��Zq�d�h��;6�x������!�6�붵N�� ��6�!6�J@��b��4u��~[��C��ob�OR�6խ���N6�����hT�S�e�'��]��}�D��7��64$�5R䏶��6$�:�!�5P��di�
�r�6������nb6��Aж�y �;�I6P�6����t�4=/��PҬ�?T�U���=��1Rv�d(<6r����z�6v����2V"p5xp=75Nն� ���|5���5hu~4�ղ�<�;��-*6����E�5*�5���5=µ�ޒ5����`6ۮ�6,c��p�6#?o�j=P6�3�5�'ݶ��X6��ZP�8���v �>9�5��Զ��=�q����4� 6(�	���Է�6X�u� �D����4 #�4{�6֜<�t�5HZ���%�6բ16�5�o�/�Z󢶇����,���ϵ�_�5䉓6l�=66<ζ�R���"�7���:x�ס�!	��?ܩ����5�)a��l�6-2f�B�6�C:6���ty�3 �4%R�5Z?50X�����5�%5��Oٴ|�6XYq4 �Z3`K�����q:6�M�5�׵�^I6T���|����75���2j.5f����ί���5�_5}�ⵠ���J�5Z6�4��U5��׵���4��5@�Y4x��������#�z{����2���5�R��8�	5`¡4�(;5�n��1�5�Cv5w��و���s�Jہ�J' 6���W$�@|�Pe��,5񰵲�5��5t��� �i5��5F���F�3.�{6f���:�A6�H6�m����S��6d5���ЗF�p�Q��M����5e��5��B���!6�S57�53�^5 �A���N�H=6$��5MR��ĲD�r�<5�.�>_�,����s�5Օ��}45�)�5�0��r#5���� �5j�ٵ��5pI%6$~>�7��5f��5��j5�2W6 *�~/@�J��5@߈3�h�5^�L�~D4L�h5�'5zÑ6i5K�25�5گ5d+�5���5�oR��_�5���5���5�e[6��%3b=�5^-�6p"���5,��4��)6DB36��~6��r��C,6��5ZP�5�)�D��h������5�z�4DL��{�5oPY���4�ϵa�5��\6����W��5ڤ/6�`Ƶ�:� �Ե6�-5�/4J��4��5�wi4� 6 �25�v���-�>��5�)�1��5`E��(�����3�
L�6���5�f��)5�ܵڡ�5��\(.53��5���4F�#�8.:���`a\4�z66�8/� �e�hh�4k�A^&���44[5�:��^��dk6>�5�z�����쩑����5���8�'5�:�5��3�h�`�.��K�zf�:f�5�ʙ�L�8�(�a��5r�:6�/�4F1��V���g�4@� §1�ʵ@6c�5��5Ж53ZF�6�dµ�
6�B�5�84<+M6ߝ�f��5n��Ѻ����5�?3,55 ƻ4 VS��4B6����(Q5�j��%o6[�1��h6�,���� Զ1<��=,7u�̶�G�6R@���!5���6�6��5%Z����5 �,����ZI��n��R=6�7�6���2ě��\D��)6U��6�1���2��nI���ir���s� O
4��4_͵��#�Ѷ��Ƶ��/ĉ6;��6�����]���6��t�)�6Ӳ����/��Y6��ճjs���O����6���5"Bl�i7���5�5:6���� � 7�/�Ds�j��!7����26H��6����O�D���6�j���K6�+6}���-��6�s�5�B6�zQ�1�����0�}6N������5M�ݵAS6��h���6t�6�y��a57\<�6�6���-���D 6?y8��4�r5��nK�6�����S&7'�j6%F�6�+���܉���(6r���?%6 �	4�Q��WI����5�W�W�����6R����<�?���]�϶i6xiV6a���/�6n���IK��0#��6
�W6�	����M��D|ŵ��7Hɵ��Ĕնhs�5��ݴ�r�6�L\6f��5�-�� A�5<,��X��50�{6�b6��6��y�wzx�\�V��@ 6�H��E�6H6�6t�601f6ʀ	�X�5�_̵���6�X�6�.�U���a��5�G��Z�:���7�����Ӫ5���59����5���6\��4��8�FV,�5̶l�)6|�'68��5j�e6�޵��5Sƫ6�
7z�X6�_v7�m{6���UJ7�ȧ4��d�@s,�_v��o6���5r�I�H�ʶ���j7c���i6�_��8e���>˶��,]��x)7�h���X�ڹ�u��A�5p;5��	�Svj������k����{6��5l������6?������%�!�����RUl��)x6���5�%16x��6s��D���4���	72�6�u�fa�@���Ŷ���5�M6Ɵȵ�����6
�t�ţ��_���VD�5�ꄴ�O�6�c�}�8�r��ܤ�H�Q6�����xٵ<@5�(z��(��6�4� ��6��۴7|�x�3��V�8�	���V�D�6)=��㲀6��7�N^G6.�q5\YD��z6 j5�_"������"�6����$�L�N5���@6f��6付��25��6�8����w�h-g5��5/����W�6V�B6�~�lZ6�]�4�w6��o6�}�5n�6�:��@B��O�6��6l���37��c��+��?47$'B6�)��Ķ�7�Kn��)����5@��=�4���64��5��Ŷr�����䐵P!�4ߐ��_R͵
���$�{�����U��6�h��钵&�6�D�}?D�xJ�5Ў�]V������Y߶Y�c6U�t�b�7 �J6�Y�50u��G���'32�K���6�°6h����a��052��|j�����600��I�� �ru�5��6)6G��?��5��W6m��x��6��d�b-6�Jv6�5(A�#�5�����v6)��`;T6}R�66b��S_�6�5n3�����\4ֶ��6����5�2;6�Oᵪ��6�Ż�ά�7�@˵M�{6��*4��d����6��@�6��\6z������6����6�ż5 �ҵ���Ư���O�BH�6J����Q�5��4q��@"��m�58�4K96�c.�Y�����e6�>17����Ǩ������O>�6�W����\6�鶿|>6������S�[��5i�D� X�%��6Hq6�>6V*��/�\�2֡6��+5~��6�Z�����6h<�5�Wp6�̶P�r��nٴr~�6G������5�5�ޢd�+�s��@�����>�����6�5߶��:6%p�6��a�l�6�B�3��6���5�>�ߑ#�|�5�E�4�DǴ,-6���6S��6������60˔5l�x� �6������5�拶h�2�Ċ�6��6�+8�Mㄵ�t�5�8C��eb6`r6�@�آ�4��5�aY���6$�06�.6ʹʵ|<*6��&�D.0�LCN6�T�4Na��xB � �t���1�z��6'_A6���>j:6�6���K������=��̶�A����C���6aE)6�� 6�%���&6L�����V6{<>��9^6ߴ���6d@�5������6h���АD6��p6D�6�@�6C�f����6BNF��\R6��6���54~�5f�6���0'�6�j5<�ŵ�掴N���5�5��E5���5H�5��5�o��;�5�ހ6�8D�O���4�f5��H6�z�B�C��Ө�>zG���y6}66����%����7�����4�w�3JP��\m�6Lk5t��$�<� ��<6Рd5Pg�,�5A�쵈��5}C?5��w��6X�'4wA6��XH��\C6���5�3S6x_l���5o�96B󅶂S����{6А﵄�3�6N\6�56��õt����@<��j�5|�E�lZ5�O�50�����5]6����Z6��6ϯ9�Rf�6��5أ��P��6\fn6�lP4� �5tdx6���1�5ա�5��57�5\\5}e޵Њ�6h�5r680���+��mJ��	���ߵC�6�µ@�ݵ"V�5B�k6;�5ӛ(6"��6g\���5HUS6
�v�X��5zz@6S��I���OŴ,�5B���6v�06Ud�5��5��n5Ώ/��J�6�L�W6��� �92���6Jf����J6H�ٶjoP���5F����2���_4nMj6(�6�ڵC=��h)����h릶��N����5�`96�յέ���u趌6�L������6��M6 d�5T?�5W�� 6��4øH�缱5H���BMb�9�6XjL�@!I�s� lR585fk ������M�L���5�Y��6�g	��<�� vC��'�d��5�w��g?C���3P"�d�5pۀ6�E ��E0�Щ�4�#��c��Vk��P�\�@�ϳ1>���Z� k�5^��&�5X�,5�Ā�lf7��´�7�l��]�L6�饶�N���k�ʁ��&�4���X���408�6��6X)6��f6=���L�3��*ܶ�55�Z�`�޵��U���5 ��6nRK�Y>+�� 60[@5���5�OI�V�f5S6{�:6�!C��:��9K�6Q�Ҷ�_5���5��6(p�����y�^����ֲ7��5Ma�6dTm4,�x�5�K@6��*�����6 ��3�K?�zc�zPx����F!�6�-�5M�{�4766z�������@'�jc�5"75޺0�
$ڶ������>6pْ5p��5`V�6��5��ֳ�p�5�6����\��z5Z��4��j6{ʐ�@Z6q9T6Jp68I^6<������4��i��/�6`�ٴ�D)��j�6�K*6��PR�5�o�6�/E�Lb�5
6.�����VH�5%AŶ2�86�/Z6"h��&�Ѷ�k�5-�
��� �3W��~�m6��r�_ ��Ț5�l�5@���l�6�_l5��	�u�r6P�16����9�<S6�E^�'���4�V��5-�޶���\5n��5F�)6a���,�6RW���:�6��S6*;�lLA�@��6��6f-��/擵��ܶV���]6�w4�D�|KP6#5��͵se����U6�op5�6<�q��t�# }�i���4�5��6`��5�I�6�E��v�5D�z����3�h�D�5��2��ҵ�}�5q��
Ͷ�,�5x$=5jH��Ds�@-��^6�N��_��>ѽ�f�'�nR����94�W&��3o�@�i5"ˤ�s�y�D,�+�����5������`�(j6H:�6[0��w�$�.\6\�5p~���	H��54�>�S6X���ҥ�Ի�5V�8�#��� 8��)�6��,���o6lM�5�(�4��4@�����C�1P�l���h�
5�|���@�g�6< ���蕶��;7�8�5ts5�s�5$h�4��4��5�����^6�_66��5,�6>i���YF6%�5�ၵ`�i5�G�
ĭ��͠6Lƀ����5���56�B6ev��ػ�4��N*�箁4~'7����� �l� Nβ�͂���!�(�6 ���+�=i5�&ֶ��5��'6���n���ލ5ps�65�5�A�5��4B���?��"h`50� �󺱶R��[�6L��44c�5��1�e��6��6�[16�}��6�������4�0�*ѹ6�2!���H���t��5h6Q>16�։7��6?o��<�4j�'����go"�wP�6���5 �~��W�6������6�aR6���4l~o4z�P6�6��M���~�ܵ|O5�z�6��B5����0g�-.�6���8>������W53E6s��p�3@�ȵ�kD�2D>6��5~I�����K97�,ͶE/�5�605��|����6"j ��n26V��6�R4�ٵ���6�hT�A�6�6�y�6��5��58�5��X4t�L6)��M�6L�r��bz5*�N6�ն\�j��}����ڵО�4�1���5W_��)668��z�a�Jc�6B�{�7��5�e;67M�������6�R5 �h�z�J�6��_6�m4��6>	���L��]�T�z4�6p�?�����Q�6��B��#�l�d6��Ӷ<��6�^M�OƼ6|����kŶ XF4��5���63h �4{[�p�	����^5���邴��z%��M����:��pP��V�5,����6er�'��5��ʴX��=;�5��j����6�'a6J�¶�z�5�����$6�{�3��76�H�6ہ��i���� 6N�`6�-x6<��h��jf\5K*G��06���4T��6d��5s��5�\y5��u6d'z�V<^6�։6�ѫ6�v6�e4:����W6�=<��$6�.��z]6M踵Xxʴ怵6���KH)6��*6�Y6V�ŶI��5`/��1w������"�h���bŶ�
6��*��r 7����5�5Pp�5�a��F����ĵ�1�6����!������5�Q6 ���5W��6�ED�<Gt�1C�6��6�u$�����7���,������z��U�ٻ�WΡ6���5a���a6^�6��6��~532A�fP7$i��X�6�+����X��6	r��P*:6Bϋ6�>�6\�� �Y5��s�";55E�6j?A����6~��'��W��6T#�5��\���i4rP7_�36S�!�V�6d��6���6�6�D	6RB���^0��'a6Q�e�!�w�|�5��#�5H����6`�ȵ́�5���6�ᰵv��6v��5�[�6\G5ϡ׶�
��w�6���5�V=6e��6P�76�$�4 �4�O�"q��}'s6�-)6h_�6z���U<��7�6Ɛ6K�e6�p6�?5�6 ���K6]�t����~u 7��6c��6?�Եjf��K��4.�|Ю4�Q.�訉6~F��4߶�g�4��m6*a�6��N�t����Zȵ$��6���1ö`�)6N�\66s.6R0�5�`A�_�6M<6��3h(+7��SN����5n�%�%K�6���z6,��6�1ɶ�L�5Э��$
�6���4��M�6�6�"�6��6(d����6[8"6��6ʡ�ʺ
6�\B�E2�x=,��|M5�b�rjF5R��U 6*��6�]�6|/��c���7P.����06�ݶm��N6v��5g��6�K��3���k6�l]4���6xҤ��J�5p�4$|���5Ls5g�)6�qϵ��-��j���H6�w���<�I^6���d6�3�)a6���$�4�\�:5Jr6}ē�
4|�S^����`3�6$���4_�5jA�6�T4:>p�l��6{<5qq�6���7�M�"�t�O��4ø6o!'6qF.��]�6�b�6�6�:w5��$�
4^6���6�P06p~��B���y\��Ӷ���P�Y�?�$���?�L���jd6_?6jW�5¶H60������5<��5th��H+I��H����jo[���k�v��l��4P�ٶ�㭵ܰ�5Ү7��6��8�2Q���.��#���ȟն7����^�i����,6�<� K��5����[67.5>$�6���W�y̶0J�x<۴�#����5��p���/54E�4ys�6��(�?Z��4���!�4ޝ)7�ф�X֕��K׶o��6���� �6X]I4�>��i��V5I6�oضBӫ5��5�#��t/'7�? 5��J5Nq���L�68b@3`D���?��qs5�����6ӱ���1=6x�U���?��{86��6�8��L5��5�ft�̃6:�e5��6�Ǚ�;����<$6�7�6{��6 �˲�?6?j��P�6{W5HbT6�3t6��36�aC5���6��6���,6��4:'�5�Ķ��5��d6��6��\�Iꂴ>)ʶ�35���>a�5��5���>bk5H�4�	u5X��4v�϶�b5C]�5�I����B6p�(������?6��5�ْ��a�����ly��W4��������Q��ԉ�6jZڵ8��6�삶��6�+6Hߴ�����o6��6�I6�'���8�f�s6�ֻ6���qY� tS6�>�6*���P��6��)6i_7�E6ݞ9���O��
M�cV6m���M74>�y���0�m�EpK��wK�2�6�ц��[���ˋ�=S����υ�2B���E�5�ϐ��r62~R7g�c���l�vM��F�t��~�x+`66o�� h��w��t����ȶ�� 6R�/�4h��l�6��5P�Z4�Y�4^87�ړ2�d�P��v��5ʂ�!�ȶ��6΋���Em6�X�6��H6Id�5��ԵRw�4YU�6(q���8������%�5�݌3[����\�
7��µ���N:�4z����5o���Ĥ5��76ѿ6a	���P��|;6 Ε�6�7ﶁ�7oIT�&����6��ն�����V6O?ɶ��F6e�6��γ �e�@��6~��ß涗.\�=)��rO�.(�h�����C�� �5
�76 Nش��b6�T7B�6[Q5�O6��F7�k�����6
a�6�P5���6)ls���϶[�7�жН4�ݶ`�6��*���z�l����;�6�#Y�.%p6��Ŷا�����6`(�6��:6`Q��Ծ���{�z*��@���['6�	�6F��dgy�V��6�!�tL7��5�Z���^6ѽ��6�ۤ���6P�7�P�&���6��X7�ص��7��u�`w�3��������0�E���6(W7�%6�PV���6����N�6_;B7�B5?�Y�j"޶p��4�H�v<-5]��5B�i��Ǥ���|�.1�5D6"��[3�q�6Z�]��5�	����6���/૶Z�C�z.�6�jҵ2�6ɐx��a�6���5`c���K6�h�52Ƶ�5�s�5ɒ���#�6O�6��h��Y�62����ɶ�u66O˵�F����5 ���yO69X�V���0�6'sT��I�F���\�3�7���6�"�56|��x"���#7��6*u���I�5�d7Xb��*�ߵp|z���T  6��0������-4%:��#��.�6�o�� �6��E7c��5�6\�Ĵ(8k6𦵴*�.7��_���n� �5��2���?�F6�5aa%��g�6iw���6 ],7��5��5i!�� Z�\��6&$�Z��6!6A�g6佈���6��I�rh���47ͥ(6&_C5���6��P�>�϶�G��H5�s�M����C��6���hU6 m�5@��6�v7UI3�
2'6M��VX6��)�[�D6�����z�L8 6���5D�27�抶J�6�K���?����6�Զc���`%7 )ҵ�7W��6Z2��U6���6_w���������ڴ�c)6�?V�0��3�'!6݅��8kR���B6kuI6��6j��g5K�T5b����nе�ڵ�F 61娵�Ur3}u��`浠! 6ע���Y6�Q����5�<�6N��::-��畵�dõ�ݪ��mӵ�����u�4�%J4t�j�%̐�ʗ�4lܹ5N�56���5P�6�X63�a.�����5���	�ֶZ��5�2��6y3�5W�����ȦK����5`�44���dε"]��	
5�!6s����
���ڶ�&u6�:յ�Z�5��6��>�������.�o�.:��?@6lө��-6��T5����+�t��5��5��5�t�$�g6��4e����6�4,�!5��(��V�-+�6�'�6Ӧ^� ������̏6�_�2b0%���!6���(}�5���dN��266u#6ρ	�fa�4�u���<&5�Jz6�6�4�w�s8�5H����o�M�5 >����F���-�	61���u�h���5����6�7��'�̤#�F6E�
��5��7���4j�5�3�6k��6��6\	G��ٴ��46�6~g�5�=���5�KA�Z/�5�&35�S4�U���|Z���`6V=�&/���9�5�m��z��ȵ|���E6���&���<�6�s86�nS����5�E�5����4'5Ĝ<����6�<6NN��8X�5<� 6�
r�*�G��^3��j6����ej3�s���}賬��z���w���QW6���U�59�5�j15��� �:5��9� �:�p�=4>T�M#+�Q��i�5n3��!��ף���ٴ�����6�]C5�ƚ����%�25���X�<��N��dy��f|�i���$�x�>�h��Ì4���6s�n�\e�h9y4�k�3�e��S��v�74�l:�	ؿ��Oq���	����6����P�=5�hͳ����pH��4����6%7-����P)4 [��3��x���r��6֬���6y�p6͌�5�Q�6A6d�6�F���L�긮��=/6F���\�6�Q����	6ޔ�6�=�<��`��6T��6��Z6}�õ �ڱ��7���5j�
5*����8P�����6j�>��c�L^�5~)75��#6�� &<3�p6�v�5�g���7�R�(�Ί�6~g�5&b�6�
62=���J�6P'!��µkj6�3I�Go�5�5�j��6p�K6�H��,ey���6�8+5�2#����3�㥶@rJ5�5�53h�� ��4�2�5$$q�g5���4�[ж6�5S�06!	!5��4�%�}�*5�޵�kO5�+�214r�6��6����Xj�5�6ۗ�TG���τ������T��`��6H˵&x50f�h��6S�VC�⺈4����6H����i05�[6L�ڵvR��+6�,���J�1����o��5ž����O��l�6,�6h/��m����^����x�f����5���5$�����5H2�p�5_6F�����$��(368(�4�5�4��� 5�Cl4�g5l�5>�j�I�����4ă����5�[�5XzT�J�5��51��-m`6�F׵�U�6�>���/��J�6ر��6���6_��<㥴	��v�!6h$i�����_�=������_:�M�G�2w6��6�"�3l-��E% ��.�1�6$e�5��d��"�>-6i�4I��5:a6�_�5�57|%��	M�ڱ�6�^6Og���17���6lh����  l1XZ05?��#,����b6C¿�Nς5g�W6�&N4p�D�t8�6�|T5�r�5�ƹ5h'�6��a��+6$צ6����6�������5�đ4"Q��a67�{�V&�=�޵4n����5V���6�!6Ϝ6v�6R�6�=�5�Ş3�J �?�ٵ&����>Y�R`�5 ��5��b��6"��E26^;^6H�t5�575��6��i�5����d�6*�����D96��q���Z�lN�4�������~PW�J�˵�(�� �Դ\��6�y;�.�G6��-60U�4땔��%6B�t��v��mU5�K6<�˶���4��K�ܝ�5�.�6W���b@q6D����^6t�,�ꏸ����6�x���y6�\�5 ���q�5S肶:ڑ�b'��-��6(���dO�5���5�)���T��
a���W-�ۏ��a��(��5'�1�Lʷ�`8P6vv�6Ŏ5�Z�����dk�������M4 �2#��6�J�6�t��:�;��������6�wk�
��6�+M��$�6�6����q�f6�<�V�@�4
6�#�Լ�6� ���A�6��w� ]�n�5���$6��D��b=�F�6�����u6 af��͵���<��5�[e5m1o��q���U6����I����ta�5��`���������Q6�E�4x��5��4`�O4d�5c�}��5�=�5�O�����+5�:\�5J`"��DJ���6�'v6JL5N���7S�5o��6�>���g�5�]���<�l����@�6��5��=���
���^�ݴo�ؿ�5����Ł5@2��׶�De6x�`��5��i�Ƚ��
�T6����ɴ6@�5N?����R6l�6���68�J6d[5/Ru6K���RZ̵�M����>6����lo6�#w��˙��ɴ��(�t����86�BH6�l����6��6c�6 ��0�|��3�>�8����ƶO�66��Ͷ�>6��O4�`����5�q��*�~6��6��*��H6*��v�ҶVtY64���ྦྷ4t�6D�/6(Qڴ@2=�^۶�\���S6Z\06�b�����6��U�U!����3}�Aw�5 ؞3��6���a�\6,~�6dN�5!��6 �*�)ie6\��5�5@z��v:5E��6��5[�	6�{\6k\6Wdc��((6O��6� ��`x6�&���07� �c3��4o�6�W�6D�6<�6^e���C����I6���5J���A5L�6�mv�����4C�p3�65�;g��k����Ҷ�s6 �	��N�ll�5L�5Hc-��׊5��� }ߴ���5���6(�o��(�6B
6�i5�)�4`*ݶ��V4�U�5�����O��hr��⤶ ڱ=S��xŏ�C��5/��qĠ6�&�5���6*�\��E��׵�v�6L[6�'@��*!6I5N6Ay�6(#�6>U��(7�	s5�
6�U^6����%��6��2��2�6��`6�ZM5���6��5�#���{��o�����6�+��DR6���5��6�֢6p��5���5�c6�����L}�Z�?6�w73F�8'�5��5����6���q��w��6�G�6���5!?��ډ��D���6g�6�㧵�p5g�q�4��\6��2�u6#����6��6hᔶX˵sA�6u��� 75�������;����3�H��ޙ��b*5 O�2�JX6�K�T�{6 ��4rz�5C��64.f5����y���׶�� 7�!�5�徶�j�5���4d��bmx6�2�m�7�E'���by�d�Z6�j6
w�5�r�5�6�<�d=��A7��I6 , 4�k�6����Z^4Pew���5Ԓ�6�LD6v/8�dW6��6�o��	����y�5܌^6�|�6���XM �t~�6�L�4�Ƶ�;�L6���5�g6���\鐶@��6f6�D����6l\���#��t�}6�{������e��6@+���5�����B���]���F6ܸ4(��5y����5.�u6���<���%_���6$ME�ܑ 7��5�Z���3�5���g����xS����5�5uy6 yA�l㴾r<6L�87�g����5`Ѹ��|ζr&��������6��3�� 6��6���6�U�6�K6�"�d�4��`̴b>w�|Ͷx����6C���<�5l��6X��3(�ݶfE7���ƈ˵�o��A��63IC6��ȶ��e�Ps�����6z�A�O���N6Ё�(�6�䉶*�5��:��6F��6��<5p� ��:u�ꃨ6T���|�ö�I��֚6��6�#7h�K�h����5�d_7H��6�3�|��5�♶��[�BW���_B5��3��^���07�޶����,�7�Sd��c��F�6�}�oZ77�u�:k�6T�p���7<C]6-��6�炴���'7}�0��HJ�xT��#�6\޴��&��">�c;�5��6 <t1@�ֵ��6#@�6X�6�]�6�����6��S4Tjٵ�8�����656V5 �;�.L6���5�D��4eu��|յP6^�(j5\����>�]l6{[O6O�Q���5Ď��im�@4���n:���6+7H���Ƕ��Z��6l�.�r��5ρ6��\�[b��ү�����5*��66�����e6��5N(�53?�6���6��6
P
5 x涀�X4P߈����6��T60	�4�0x6{.H6����c��6p�48�j�TQw5P�������L�6Nr*�H���8557f�5�Q&6� 7۞����u��[�6�瀳<DL5����26\�56���5��6k۶��A6��=6���6�&M��7>��KA6�l	6 �D6*���k�]���7�5�`�j6�H�60WN5CV_7��m�7�6��6����
�K�a��6K���|o���g�������6��u6�҂��v�5�|�F�B�6<�5�o�¶L?�6vxc�,f�6�ߏ5�.��,��5I��6��C5��s�5�Fk��}7Q8�<ҫ6�}��#7��S�*�� >��FXS6�d�w`7��6�U_5�p�6��]7S%��Zت��̷�h+�5�2��P$��wf5ZW�!�36��6ҺC�(�6)ݩ6޻��Ts�5��5.e=��.7�p5�P:6~�J����l+ն�‶ ��6�NC6_~�P7ek�0*�4�Z�5е�Ac6Hԝ6���8n�5N��5���6n�6z�����5��y��|36~E���9�$��5�#���\,�G�еXiQ�����"�����n���F,6(��5(Qõ�F6f�����66�8���/6!T۶�mN�l���Y�v�6@6R�Q�bB:�V5|:��PѶx�c6���6d��5��5,�n5:��6?�Ƶ�h^���+����6����� w6�����0�k�6�a�6��k��66�X��~���Y6�5�4��6Y�����5F�<5�ɵcնbu2�����b���J���>���7���Z6h7��X���\�p?96;\T6Ī�3�����6 �m��� ����Y摶�{5�����A���%"6��~��y6�5�6B��� ��1%����͞6�-56�_˵��Ķ�:��I60C�4�/õ��ק#6s6�Aյ�o�5;���� �i��6z��P,��1)6��5֑6{(�6�)N���5�ʱ5�W���R���6��66�7�7��W4}��5pB�5b�B6z>��n��6)�~5HzƶK�5F�ڵ�R7b!�6���6�d6GUu�`{\��'���϶�06�*�6ᵈ~ǵ�4�15y�;6��S70�Զ"cȶ�<[6���6���3 f�3n���*۳��@�Y�Z71;�D������3��[6����f��6�����t��ZI6ለ5�r �j
x���5 +]6�s�6�l5��˴x�5_�6n ����&���6'�@ 
�Z���X�`�5�6���5P�<32L?��z(��]�5�}�����T(��(��6tu�6IU�5�D趵��6p��6jj6����� �6��6_���~6��`K��R�X�6��6l��O��6��6k~��{n7������\#�E/,��|��J 7`l��]�B6=�v6k8�6H%5v�t�������i5�˶ H\6'��6y���@;6���5���6 P��Z5�o�>��0�6��V�d#�+�47��r4bk��?��ë5��44�����;I6$�-5ђ6����7�{���L�k�m��6,2��ǧ6&:V6xg5[5�x��^�6�b�6Gۻ�l_$6�Ζ�Su�5�#<�� �z�5Z�64�K6B���/'��A� �ɵ
5��߲��~ 6ҋ69H5�Gִ��"����5��W��en��A�5����|�46-�6�]ѵb4$�
h|��"I6� �4"�6�eV6�=5_Ya��᭵$g�6ع�6
���5Kr����/-�� q5�F����0�p
6��60-:��<���2�����4��p�ż޵�ek�f�:6J�;��/6��3QN���0��f6�0A�*��5\>�5y'5����۔��ғ��y6:9���RR��C�5���5�_!�����H�4�!���C68�����6<�6�<Z��t�5XaA6<\�P^!6_I:6@����6� ��Nô6Rq�6�E�5@t���o?��%b�` ��b﵀���{��Ę4.�X5Ùy�F�6��I4bT(�]r����5j��G6�/�5��a�M����5����K5DX�53>/6�C{�P��ѫ��X�:���44;�pP/6Fu϶�j��~�)��{G6�ތ4]%��"/v6�o���b���5�]?4���6��5���Y��z�5�@ ��z���Ê4�EA��^�4��J��&�����5Ue����5�`+6��۾�Q�6�E�Y�6��I�6>��4�͢�?����6�b7�|���Sص~Xյ�0�6�k���-�6r��`v�6�g�6�E�����6mߵ�?���h)6(��5T'6�06b�W6�v�|&z6(��4�=\50@�6'H�6��P�61��5T(���'6�ǭ�>���4Ӛ�tF��8
���e6H ���@6��B�I��OT5p_޵h�h�6�C��#a�`d��p�5�L��Ƙ����մ X��,L_6<4�P��4l76���4��8��6��"z�5�K5�G 6XB�5��(�Z�6þ&�U��6nً6˩6�j���ܶn�63v�6��6�Zv6���'�6��F6aV3�#�6P�&5��#��/�5=�5��e�L�ʵ�9�6��鴕Ͱ�{8��v�5���5U6������j�|6&�16FV6ڜ��<�d5$�r6����⹢5�}���.�� �9��k���@u6�>6Ǳ0�Uf鴀����76Hw�6��h�S68�۴��=V�a6�v�5.������4'����例85B6�k���0858�5X���:�N5@�R���P��n�5��6�+��*M��Nj��b6�Ʋ6J��S<�6:3%��mm5r?���y�6�_>6��6ݿ��}!綾A�.��� ��3��<5А�6�/�6��5{�E۶�o� �/6�U\���5
�ܵ�憶�9дf�}6��N6@9D�J''6̚g5@l���
�8�6���6��17�����(6�I��ҙY�$M6`J�52��tpk�=����6|�p6z����5�ḵK�a�+��I�j�=b��q���\W6���3&m�5\��5�ں6���8iW6��5�N��#t�63�6z����r����6�.5��5z����	����6xdn��!5��5��,62eL�����;�z�d�ᵌN65��6�Fw�����Sl��͵,�q5��ROb54q�6x�5�U��{7��51�C5Jr6��)6yJ�!
E�d>������t��60P�5�x4��.6���3.���=87(�6 1\����55�#�f�5�+��V7Hm)�N���L�6`��U/w�`�N�[eS6R�6,4v���6��@���ж4�I��獵�U�4,�6G�1�K��<�5 ��1x$-���g6�678|:���s5p5T��^6�L��)�<�4TӴ73�6������5���L֦4ʁs4s�6�6�^�kp��~��\�6@�l��S5��g�Ԃ���h�6@�5����:��(5ap[�l�6�������~��5�3�46�%��4�P6�v6&ϵ��e�~��ޔ~6�2�6�"6Q�5��Ŷ={�6�':����+b����X5ZS�5iO6iF��L����8�63��X�5Ng[6p��5�nY�9�#��~ɶ������-��lۋ�?�5��{�� ��9�[�h����gӴ��5@�354��5��7����6 ߱�"����j6�5Y���6(��6�6В\4�U���0M6�򏴠* 2ᭆ6<�6l�56x��4�C���g5ӷ��Z�6=~5ݣ3�r�m���z6�'W6�G�4�5 �h3�5>����~��:�5�>g�����49z4ɳ���H�=ڮ���p6�g����5�1N�v�?6\<l��}6������b�@(6o��@��5��ȵ��.6R�6%�,��_�4\��4�y�����56�;�`[��"���&�63�Ͼ�����5�|6�����5���'�69� ��!������?c_6��
6b2,��m6�7�k̵��#�۩�5�C 6\�����6��ﴍ38�F�;����6�D60�,5,�����6@I|�|!6,lѶ���5�26��D�l-յ�b5`���u7� G4[�<6�k`��"4u�6�F�5����2,�Z�5�O�5�3�6��6�5��5���vO��y�7�Z���� �ؔ�4֡�6N;��-ƶ䫵T��6[�4�;6Q�4��7j5^s�qAQ5d�6u窶��ѵ��l�D��5H˫�`P�5�q�"�&�dX5��K5�?��@˴_*���1\50��3���_[�6a}���Q�KA�6t@�5kX~6 ����߼48U���-���t(6��"�^����ٵwr�5�.5 e�4�U6�K��'e�5_�V6(v���L5�-6���j5D�d4��6�"�+��5x�F���t��F� �23J��5���6t�6���4��5qlh������%6���6�_6��״�4x���H�p���o5���� A.�$d�5�例s	6}�6J����;�T^�4�Qĵ��ݴ��$�>�J6zfR5��4�q�5�gK���6����5)w��%��4���5 ��1&�@����5>�m��N8�5�6|V��¡��6 %�4�,�6ٯ�6	��5�
6̳�6%��6z�t6����;�]6.�\�. S���ж 986H�ֶ"�5�q�Q.��5h�����4MY�6�[��~���X6������6�aܶ�C��|Y06�� �2$ϵy�P6�~��J�6��&�؛6��%�3߁5|W׵�)�^?�6���5`!�6��H�va�486Hm|�t�M��L?6��5㷈6B㫵�*R5o+n5�52F�5neŶ�6����D��k6d#5�'�,EH5T�Z5�w�64Q?��6�6�C��6�w"6N5�6X���>4�6�3Gk�-�-���76�5>�6���68EW�L����6Q�d�z趠l6��<5��ε�$��U�s6S�o��N����+��2O5%s�����@!�5�ذ6���4�&�oѶ�K56�5B��QE���y6���h��5�M���ֵޑK��дz�n6�
���V�v\5C	5	��5�6��6�|&�!�4��5$�6l����5�6tY;3��5��µ�U�5��6� p��X5��6֦�/<"�-n*�Ĭ�4n66�*O���5Z�v5ȁ
�y4-6*�ʴ���a����k�6�Ι5���x��<J6z6�&Ҷ��J�^%�6��J60���:]68c7&&0���Y��5G4��5÷5+��5��6�(�6���E�� �O��ї3��7�i�4�5�!6�R6r�結��4�cY6�����r5�T6�n6Ǆ�6*>�6V�!�jK�5E��6�I��t'��0F����U��`?4�R���x_5�u5j��4�'��'��̸5�[���J6^�F6 �`�~N06��&��s/6�$�3>�T�0⣴��4PR�6�ֶ��6��5`�5(����n6k��6������{#� ��5�P�J�6���5e�d���7������T�Z�Y��
56|<�Q����x����'���:���I����5�,�6h��5"�6�nW6�EA6'�׶ص�� @� �5��=5��{����4��)5�U����5�>��J���X86�?p����@��j�6䤺��#6�����s�e��6~Ѝ5PS
59� ��5��x��`�
2U7���6��6C�5w��+v�6�ک��<p��_6�&ѵ�v�5����H��P:�6�7����=��d�no>6�ld�Xc-�\�)6a	�>t��7�#X�d����6z+��<{!5�=�l�z5|]��=���ɗ4ʦ�6`V<�p4�!n���q�4����=50P�6�6�x�4]��d�
7�a#5XƵ�#ԭ6��4h+86�)35���6&n����R6�	�6�g5d�4��$w5V��-�ڲ�60���,�2��6�e��B�5�6���6ή�6��aU����6�׏6wTw����5$zr5@� 4���6�ۥ���Ѷ^���]�n��4�G��'��My)6��5П{�`�δ���6k�?��Qǵ�Q����j���6%˥5@Q6��7S6h����ܳ�`?4,��Q�5E�� ����fd47�4�a�T�~6�>x��u��@���*�6 Р���6F�`���߶��=6p)7��������X���ͥ584J�� ����^���6fh6@���=��\�62�rZ�6��S��A	7��5���6؝j�ϵ���66:ƶg�U6�16�ZƵ����~�6��#��q�����5��Z�C5���MtN6�P�6�p�68�ǵ'�v5~g�F��6��5΄6��5`m��@Z�2(����6�m����6��ҵO0�@9�3������~5g����O5��d6V �pK���R�8�3��~^6�>�5�!���:���s�5<��5��Q�b6�~`�6u=]���x6��@��Z�6@h�5ɮJ���Ķ�疴��5��V�5�ch6*�&6���4� 66rc6�:��H�t�t\�6�	6V/���5gO*6�W�5�C����(5z/#6�6�m6maG6B�5��6zE�6���6�%���Դ��6�95��j��E�����#6��j�]�6�{[��^D6�Ǥ6�յ���6|]��ŵ>)���F62,���5Q�6N�Զ�k�Ŗ���5�_)5˗36O�4"�5�cM�6CM��'˵h&�6 �v�6���&k��|�(�5���5T�S6��Ƕ�+45^q6��!5r�5\����;k����6x��,�5�L	�Bо�^1M�)�e��p5/���A���e;�j�6T�Q5������5���5d~5�R�_l�?i6!�X6���5�6�4��Ѷ�)��s�6`�q��o]����h. ��> ��[���u�<P�6��59HX�zw=�a�X���4P�7s�p[�4�5��:�XO��|5�O16�t�5ay#5:G��P�w�Vȡ���4ց5���5�LM5VD6�����1��V����%U6d�=�T�56�d4�o9��wg6	;5Bu�5>���@Wb���j��#�s>.�4�
�P~�5 �����|�:5�76�����薶��ص0"4���4\.��ݬ�4�\5�'T�5�6I�56e�����5M},67�'6�q|6�T5~�5�죶��(6��5z�!�` 6_R��(��5��K6ʝ"5��յ�_��0(z6r6F{�Lڣ��>6@�5��x�ĵ�	����6P���X'��x�(��`��L��JR�6��5~����%�6��6�)��^m6�'1�?qĶ�]P5���lV�Z`ٵ(�5�A6��5�ߔ6y)8�^����3C�9�$�e��`65W��5l'������Tw����5	E6�8�6�R�f���0�_��'j����5ާ�5�
0�Z��6c�$�.�,7�9�5�p6%L�6��7	;!�u���M}i����@6OL`��
�5P �6�_�V@��QӶd2�6�J�5�=p��G���)6x(ζ~�-���|%-7s�5G�`�V�6�]%�/ �6jF�6ť�E�H�F�J��S�64*����4|v�ܶgKj�ۘ6xL��؊��3��&�6�J�6�>7�x����Ͷ�O	��l�6B��B�@������4�(U7L��I66b����5��f���W7;97��L��37�}Ե��ѵ�W�6�?*5_���T�6��6Lu�5"����\�6]co�h�54�:7w�6F"۴�7�F_�6���66�ߵו��=�'u6���6l��� ���䭘���6 ���G35�Ez6�������5j��5
�77�P�D�����F�y�;4�6�=�h�X�4C���Z��n"�M257���5�l�6ɏL7jd�2e�� ��6��ζ(� ��-b7ޯ!�p��4���5w�56��6$@�6��"�*�6�����5�5{���r6~�5�е�{�4e�1�rQ�62�L�>�V���p�`U�5��7t16 eO6�,�6B56��4��6��6�S����Y����5�kӵ(FA6_�5�N���|�����j�7eO��ק�à6<��5��䶇]���a�^
�5Bn6r����卶� �6�~���Iӵ�sh��	7\�=66.=6kf�/��6_NF�L�VB}6��[ǟ6H�A6�6 -̶��5X5 6L��6P4w�6��;7��7��!��	G�8 �6K
�ԝ�\���w�c��w6�[�6]��6����j4�����	�-�h+��t;5baʶ��U�W7;���6�o����V3�6�u��f�6�D�6V���q�367���P�6[z��<j�56<!6Ȉj�L��� ��3L^5>��6�r����15�@6"�66�5p��5&��6|���t	����&�i@��L�-6�=�3�1�`A�5p=����6P����b����y6�\�6�矶Q�5�%�JfQ5�Ǉ�u�g6z�6E�%5�:�4�����m�����������~��6�=�64%n4�Y{�	_����6�ﳵ�t�֪��|M
�����X06F��6����󎍶a��5�;�5�y�54�=���u��Ӷ�ǂ6au�"�-6"��6�U�5#3D6�h�4���M)G�G1,6 rO2�µX-��r���D�������5G�6�q66����˾�>v�����
�,��5�6��}�+̈6�MP5k��`��ȕ6v	�����Ҷ��óʭ�65:�ͺh6u��D�6�w��d���PԊ3q�7��V��V��0\.�� ���|�5]o&�e�6譔6x��5!x6&`1��V�������6|��5>`6�un��Zڶ���6���6gb�5� &7�E�5Y���Ct�4,+��MZ_��7�i�#��5���5���
�ٵD!�6��y�7ƶ��5�@�5\r�5�㶴�r6A���6
[6A�}6���5��7���H��5���d�ޤ�6�d�6 ,3�7�6�A��N60֣4��ҵ֐�5�6t8��767í6o�*��!���%5����x��6�\6�Q�6P�6$T�6��6��F��_��#�6��õ��-�� ���Zs��I�6�2c6_��5�D�4
�w6c�b6d��6�T���mr������t�6���W�9(�5k{*��@I6d��6�T�6�٘60�����4"�6L4�5`/�3�Ւ�݈6�6��L1׵(x�6h��6�����ܞ�T~��G6��6׆5��5* �5@eQ3�.�5���56@�6e
!�N��5A۶v��, �����b����5x췴(��5Q;�6�u{67��6vGS��W��^4(���3��6������6�35�76��H��NJ���ŵ�-B6��D6���6�صЂ���1�L+`�B�׶	),6����<��5�ŶLrt���2pǐ�'��(���@�Y�6D�e6�Q166)#6p-25���6-9�5�Tk��v�n�;6�Y 6�L6�BZ���364<6�g�5��(�$�H�X��6��6��!6���3!�F�%����4Ym��o۳�g$6�`M�,|6J�)6pG���r���
79��5�ư�-�6����5�eq6,!��T�o�0N�5yi͵��6�GJ�I'Ӷ��5�Ə6衖6
^K�tZ�6�8���,��L:'��a6z.�5�k6TT�?h�c#�6�����v��5�ֆ��0�6FmA6�ؖ��[6@{�3#����Ũ���5Ɨg�>?�50J,6�<�5ȟ"5h�3�3�5� �*F�8a�6�*u6�5$�(���t6}z6�6r���r`6���2��5\���t챵�@�5�������5h+H�]�h����5􇡶M\�5�my��R_��
�6�
�-6p�W�]�S���5JAK6�o�����'����E68+��653H�6bJ+44��ܘ�6��D4���6��	60�Ѵ���Vε���6�v�6!A���4�5#H���m4��~5R+�#�
�l�S6[�5
����;5�<��JD���TE�DS��\��@�#5Z(�5�q��֯����S�?Ѝ��J�4�ƞ��;]6KU�+L��sӵ>�)����6p���i��6E�A���޵tp���L��(Ŷ���5@�̵�����E�[��)�6/�^��{�6Z��r��6Jo��%��+7�~E6�o�6��5��#���6�{��I�6�ܵ��s5�&�5=z�ni�����E�5�D�bҥ���5�k\����5NVV�#�5�	A6�3�4�`�X,�5t,����?�ʰ��F�5��=�6�Z���=�5ԓ��xc����6����S�l5���5� ��
��6p�Z�)�Y6���4ꗣ6*��4�r76ͫ6>`e5��A�g>��l_�F栵���6M��1.�5���6V�쵟Pp�BFe6�;l���Y6�1W6HC{�����V�<i��|�7�6�t�6��*����6���6�g�����t$6�D(7B��������o6⽬����5�Aն?8�6��+7h�5(���#@�������5/��fb6I=e�V��6}U�6���m8���*� ��6�}�6��C7N�z��g�� ��3;���ZG��X��24�6�߸5"��6<��5��i���Pڃ�#97�
�^�@�-��.2� ݡ�(��5��g6�\7L���ڒ�<S�6��ƶav@�`��42^<���6E���I����=ʶ�7g��5?/��2d�U�
�Ĺ\���>6�HC�^4�6\*�N�����\�6l�5H��6�s!6�	�7 I�3ʻ�W\��t���(c��`�5>y~62I+��~����(�ߗ7b��6'g6��6r�����7(t�6래6U��65��5H���y��6�嫶�,�5>�R7rf��a�5Ll�6��|�ybµ�	�6ˬn���q5���5�ǜ��G60�P�,5�-&�s����R6 Ar��Y2���Όj�r �6ou�5����g9�Dr�6�]�6¬��j�%�0�~��907��7���5|a��հӶpM���/7 8���7��#ڷ�.5�Ό��	�6N�,62��6��6a����Z5�"<7�.��vB7����@�4��ж��/����6Q�C���p�6�ь5���4}�,��D��ti������S�6�da���.���߶^�w�r�	6��z6!�5�5X�?7�H���P�6�b����5_c���3)7__7���38216�W�5)\��D�7�.�����<�ɴ}7 7�6��6^���]/�6��~6��6��6	锶�(A���u��7̶rx6&��4�9g��_�7��6��6�N7���B������ζ���X���X7����|��5���ie�j.׶�w�G����g$��ö�O�7�6|��o��6�������6��6�O$�@t��|Q�J��5��(7B��=���銴���4v��6�.�5 �j5e�7�v� J�5�7��5�q07*>��-�5C�)6�y56o���� ��>�6��6���B
�����D�&��6���e�昢��61p�6���6����w6�$p���+6���VU�6��&�ZV��X�6��E�A��6}LX�@-�5�E�5��h�ٴM��Dcs4���6�����5��E�~6Vsq5R�50��-�5@��p^�7h3�G{x���0� �2�!�2�F6/[�68������d3��|��Yε��7��6 ������'5Ə�����6H+��C%7�y-6o�ඐ<�6+9��77�����Ro��T?�[��������5 7s��6�-�6/@�6�x���25�885搤6Hpf5P�65�nN��k��(��>�6@3�30��5��㶔��� �67ۏ��_�5_��6��#�.}��`6����xڎ�����*�6�^07 }����6�+\�h���U	5�g]��PR�U7넧�pq5@�n3 p�0��6�*�6\�5�-��)Ѷ����������6+�
��-	�H)�67#6 ��2�۔6�x|7��5��`���K�5�A�nLg�*bC6�~b���4Tࡶ��5��5��?6x��6p�����5ԛ�5�U��*\�6xO����6'���h�4(뫶�?�6�\6��6��o��
����5�96��e4_��4�fô�����ӵ}+۶Wv�������J�4x\ ��3>��y��}�4�$6�q���"7T�1��a�"K�����^��X*�6�x��b76�����6p��P���nܯ6�8�6wLc6�k<5��6RY��/k����f��(�͵�p6)�$�S�(���E������O�5��5�T�575�}����2��G��5�R�6(�ǵw,�6о�4�!����4H�ӵ��A6�O�6�ڷ�(�6Y��|ۄ6���6�;�5Ԑl��6�ʼ3�5H��״���vk� �Q30�ߵ�A�5��ѵ��5N���E��8?>5n������5Hu��`���W5�9�,�ڶg��$S\�����66|\�5�T5��k6��d6)W�WK�58:������M�;��5!e66�6�!�x���k�����9;���R���5�Z�5���O��X���P5�XP�� ���6~�	�6�M�dݺ5L��5�/ն�[t�t[/6|�|�,̟5`b�4��a��c~6@�P���5ߟ��Ӵ g�;�X6��5��T0�Ԩ�5��.6��=6O@j�4҉��Դŧ26V��f��5)�h����5Q�5�)7�g�����6/�55�6���6/C5,r���!�r�}�b:���4'6�i��_6 �C�l ���
5z�Y��556��n�8 ��I����!6�96XtU4Җ�6K!�6�4Z6���5����عx4�\(6+�7��,3��N��ȶ`�ʹ��6h0�5'+5��267�/�HѴ��<�Jȭ�^]n�oI���:R�(�b���/5��^�d6G�`/�@˴��D6!�h�xȖ5^�5�e�5��5�z�2p�$���4DZK5꽴��f��������_26�õJV�5&����O6��Y6���5���D»5(M�5ܴ8u7�f�*��6�6��5 A���5��k6�N�5$�ε�C6Ѕc5��4��I���^6�(����:�@��5gW_� �ó�xb6)Zɵ�t�4�Q��Ȱ5��6/p���4�5�N4p+e����M��@�`4�є���~6��*6�S�6��5���5u�M��ɴ.���΄�����K55�06-|6�MY�C86�91�,�4�e�5��7p��}���Ƞd5�nҵ�ż5��K6T�۵��#6fM�5`0����R��7��D�޵�-v��j¶�!�6˨��'�ӡ��ڏ��"��6�R�F862�6�(��6tfs�g��5��h޶��@1P4,�#�cnw6?��ga6�����ī��	*��
0� ~D63s5�`6R1�.v3����^���|6���E0n�D��}�6��5$�i��26Ly�6@{65f,���%
7όG�,�y����4��/��6�
5|��X��T15�Vѵ�,5F�^6-��5�l����6�-66�F6F6�C5d�5��6i��vW �t��5�K6֝I�<� 6Ǽu��3�5h6-�M��f�5�E6~dS6��ĶT���|ߝ��v����6�T�� �ó4�60 �6�}⵪��5$���@��6�}6X�X��U��;\�6����
�5�:6��67uI�Ѱh��Q�����d�6@�4�s�4m
�5h���ަ��צe�W#�B�5�-6��R6"����y5Ĩ�5kx�5�"
���5�]ص��r��b����4�h�_5��5(�6pP�H8���4�91���T��`6�)�ϳv�D�o��`6,�3@�5�T�6����ܷ5�����L 7F��� 蒵�6��3����9��:��t���&7B=&6��5f��6���]�
��6��6�Y�K}����6 �U6d��5,Z6S�R5�D�5�!ߵ��5^z�5��66��7q!X5�E=6ɭ���Z���A��Ls�:Gȵݶ�C�6�6n6@d44��y6X���6�Z4�N��;6��@5�}6 �1��-m��E�5`�I��A"6�;�6�\4��ʹp��6��T� �6���Z�5+�	7PV�5x_�5�r���� $�61C�6�
1����5����z,��,���ً��Ť��0�6��5�򢵓��6Յ%�d�}6��
�.%�6*u��+6�m�6��6�k6uB�Æ��7"5�w񶪪�`�5����y26�rٴ�N2�(Y��h�6? �2866L60�5?w96܊��b6�J�����5����Y&��s5������ĵHj�4i�!�98�6~�6^�%6�~�6�=���6Q�{6�7�6����8���������Rx6<��60�;�s6��R6v�&6���%6�
��E�3�7��,���O���^o6p��L!(6�-C5"ޯ�H�5k����64��4��|쀶-Gض�c6(��5ɀ�8�D�����/M��}����6�뵀�/�{#6����5�|7�u��F6 ��&\�5Ē�5ӳ�ؾZ��]j6�'���4pt�6�g	5�{��5�$7&-7:�6��ب6��L*��b��6�k�4�6<Y�4���0 6�(D�7��w6:��6$4�4~Mb��A6��ٶd�5<�6�W���ز���4\�6 T�6�k�Ը�6�A���'6t㣶��6lCw6�>4�C�6Ԑ���ֵJ�5P��Z|R��y�6  �/�� �Z4�V��4&���[�5�h슴�*�5�764�6��6��T6�N˵>���m6X��6g�@6@l�5�	�6㸨5 ��2@��2AE����5E�7N>>�p�׵������5D��4 �������ʹ4p�6�v76H+��{I�υе��g6p��5E&��M�5K+���6+])5M)6�A�5�v��ڝ�x�L6������6*Կ��ֵ$$�5�Zs6p-5�/��()����6���6B��5���5pI5��A�Pg�t���r�M64��63�4���d6pl6[�6
6��z��m��_5u(�L���c6"��6 �2�_�5fE6�(�F�������������6�K��($ֵŖ(�ܬ�5ȴ���$�5T�V�(q=���)6;p6��5W��(I�4�����=68lG���N6@���!g��\�6�^�S�6����н�4�6�蓶��5��r�ߵ�f��=����۴��5(�*5(H���϶Ie7�򞶆�	6)5͝6��s�0��dOy��s�5���6�
��~��0_�؆:���%6[=m��H����ص��5��75��)6d��6��5��j��r36-���&8� �m4"���@�5ޓ=6@l �T����w�5��5@+��S��96ȏ�?3޵.[�5$t˴b2���
68��53�0��6$A�5� �5�!5�b�����P�� O��|W���5`��3rϷ5�i�4���]j�5���T�l5�g&5�g\�������5x��zʵ��6��V�	6�U�Fj6��	6��O6������D�b�4����	ݳ�1�4aG6t�=�د`5=6z�Q�3,~x5R����g�~��54����6)5� �xh�@�?�cf6��o�䴸�;4��5���G�5l�4T}յkV�5`̎��P�3/R���3*�
6�2C5�#�4"�ȵ�@�h'�5ML�50M�5�e��Ҿ�5"\5d%����ʵT�x5����3֒ǵ`��3 �H��PM�|65z�6���f4���4�.5�K�5��$���ȳvbӵ������5r��hь�n��5��*6��!����4���4�Qc�5�4��(5���5P���t�4w������6@C`�!���>�5=�����5�G�5�[�5�34�'�5Z_s���d��,}5�!;4��൦�o5��4}744�5���3�?5C��4��4@��5�ȶ�`��4f$�5`}F�S}��R�5��6��4��5 ���i�4�B6�ǉ��υ4��>5P�Q��2`�e5�0������4���B5>5���4��(5 �95�`�5 9����4@6��˵t"�� ;26��6��B4fp�5"h;5*�6x
�4�����>J5 �o5���b��5�Lʴp��5?R6P�04�v�5��Q5p#V6t�6�8�4H$�57��5��I4��r�ȹy6�K�5�6W��|��5�6�5�n5��?��?���p�5-�r˴�z�5@��2��t����a5<!6@�s5���j��m��C�6dn�4H�O5��5��@5m�6A6���rV5����cI'58Ҧ������f�H�5s���`�>6:j6�Z���~5���4�xܴw����4&���H�50~2��� �ҍ6R��A��5�6�6�5h�赫!6͖�50��5N������ҳ��ֵ<��Ĩ���k56"�6��P����6&cW5�X6`ڼ���-6o�e���+6v�ٵ#qZ6�W��D��3pi�6(9��<��53܈5.'6(�x�5�E6է���5�54V|6�G�4��5 �b2ƾK6��`ߏ��W76ʜ	6G��5j}W���W����5�Tᴀ͊24��h<6*%6��<��6�|�>�26*86��6��(��i0�GD5�7N5�9���@6��C������F�5b"�5h����5��5�܄��DX� �5D��6,�?�^�&���u�T7�5����nW4q����4�O����T���?6:15Ha��H�^�SL|�b�50=K���=� �&2�@b�T��4�6�7��J�?�C�5�e5�Ժ��g
6&߮6H����3��4���� �ʱ�G6�e�4�,�5�:�5h�*6��c5p�55"�6dG��F#�5�!?2��T��r�5m�6���4X���""��е~��5��:�6L44��=62����_P5Y��\��%�4;|ص%�X6ƅ�����6�4� Z�(/Դ�4L�]�#8,6�5��3<���ր��RK�`�ʹ�u�и7�����5����*�5M26 �<�p�&6�_��r%���aM5�ճ��"��;��^�@6�bu4tPT6��}�|����]5�6���6:�u�@�E�y���TϹ5A���a̵�6�D�H�6�"�v>��P��4^�5�JK4*6T6�܃52x�5�Wj�;��5J�5�[6��$5jf�5 �o5Z�M5DЃ5Jώ5���r5�.�5ա#���A5�+5�64���h�5�.ӵ(��6����0e�bmȵ�g��V��2S62�5�� M5�p�5�	$6�X"5X��xQ5�VR�)�8�X�E����-D�D�4��8�3Ŕ������y�16q}�5<�6�o �@�"�J�{5B�X�����'@5B��6�Đ�,���(��5 pV�f��6���4,x�6�O��l'5^��6��ƵϢ���"�}�J6ۀ�<����ε6�X쇶�7�6��E���\��A(5��"��6��7��Z6�����+�6@�44w.�g�6�z26�T�P[�6L(�5�ߞ�ΰi6Oф�j�7��x.5����(5�zF��56
	16"[�,6��y����6���6�.�l�i�Ў6��x��)�6����S�6���5A�4@(p��ӣ4P�5շ�5�Y"���6$N�4�~B�)��A�x��Q6���F�µ�ڴ5�W-6�!����D�z=��H��6�C5�D���6���5�zy���4�Iz6���Ѳ<��|�6e0�5��6�A6p�5߾�6E�
6��i5T��6�o��,�?����uW4�$7F�6�c����4��$�B�!5|F��>�� hE4�O�� g6z�v6��86Jl�D؜�������5.���'��6��5At���6B�5 S;3�O6�a�4��76����?��6^w'��W�5���5���3�Jz6���Y_6o����5�5��+7�o��ɡ��)����4���ܵ(�G6�t�5���6�6��7���5�m7Ӷ6Ry�6���!)�5q� �T@�?�Ͷ�]7,�269+���֣6�<6�ސ��W7�v�6���46�6��۶�/-��Nv�V��6� ̵�'V6�R6�):6zm�6SF��q��5҄r�)6��6�6E���0����� ��6�\���}�6��5���pT�4+|�6B�6Ae��@�6@�5�^�60~5��T�$j37:�(6d�6|:R��-J�t�6̅v�NT6�b5r>6�<`�{�6��6)�5d�W�Y��=��'R�86������Ԉ7{��Pl�=f5$���̋6X5.�5 �2�&Ե�C"6��#7��$6��6����4~6�m�`�h6�1L6�V��0��5�;,7<ܸ��A�6�W��%~�6��5��a6�۳��C̵	�6��6��5�E>6�	O5,(�6��6�˦�0f4�Av5��b�:��?$��ǵ�v5Q�;��֪6����8��n�6V����"
�B���D�X��6 ��2�w�5�q���P6���6`��4�̐�tZ"�,�5�Զ�X�5���~Z���ɶ�H�6�D��yZF7t��������8;6��}6��G6��[�(~ҵ]*7��m�)ߊ5@���{�l6BV.5��.65�l6�M��b=�5�*�6��95N���ؒ=����ȳ�����6�Y�6Ȃ5_�6��5b+����f_W���6��6]o���&�����6003���5t��5���"���W ��F� �5�!���,�6��� e6߶�5Y�������[�&�õ�h=�6-�616��G6���6�/�]B6��6����C76��p�z��6��5¤�ĥ�5$<��D|6a��6��-6�@6��-�졶h沴,N�j(�~+v6T�|H6�P6�儵��6�$�J��6�k7#n�6���6 �&�?91�`��4�F���v���2Ѷ�=.��ٯ5���5 [���"U��Ҷ6��5¦�6�.�4�A7��0��^��t�6!�V��6g6 ~��O+�6�Z6�6'5�愧��ܛ48aε��77��� �>��e6Pd�5�l޵�]n�pDl5�؇� ٶL�u�2�����5 P������̡6��NI7+S���䴵�� �����0�˵D&�6��6�3��l͘�<���BW���X�6k&7�M6�j6��Q6�⼇�:oO�q߶N{ѵ��6o��5��_6�i��G4�5	xR6��.� ��4�K��A��5 ��4L����E������6R˿���5��6á�^������"O��(����R���6�& �������5�k�5p����.��y5Ռ>5B�o��q ����
��Y4(�6و���B�5x_f�vJO54�6?´B�﵀cC1Q�
5B�D��Ҷ~)6�j<5�Ζ4����* i�4b&��o�w�-6��@�p(x�
F���﵀�4֫�6���h�Zk�61!K����67�:�~����Y�(G��XX���6��7�$���]�#��6e\�5s6$�5�d��D%��U���uR6��Q5U��6�G`�^�µ�8�5�ڶ��47h6�g)���4� ������ޜ6�Մ4^Jd����6�r6�8�������Jp6}�35M�u5�9W��2�ѭ���=��A���jR6̌5X��5�,�60�+5A�Mx��YF'6�Y�5 5��Ķ<ס��4��6ˁE��]k�h O6���5�޴����dHK6k�"��6���Ad���3����Hn�41�6����Ӏ�dI6�}6xY��-���6���6撸�ա6�H�3��6��"6���J�L6�ߤ5����5Lpx�|`5�d�6��^�"u6�dֵ�{#�k毵ٸD���c6i�L��	A� K`2��������mG�6�Y۶�j��m^K6�X5��5��B��.68`�4��1���7څ6�s��%�5����Z�K6poy4�2
��8}�i����*�o&�dK 68x�6�z6��05Љ�*��5�A6:R���B�5�N�5�����6�L��Պ��nU6X��4\G$6F��5b��o�Ͷy��5D����{�ȇ6���6Qci6V	5~��5��6-������T���QB�5{�5��5��6�y]�mɶYHK�b�Z6;�ص�Ҏ��Ϲ6ҹ�8y�5|Dl�@��at��J�ֵ<�趄�V6@k���#��9�"�5`fo4�	���e5��5�s��V���?���>�6�6 �4��B6�|�)n���&6�0	6����n�޵G#�5I�Pdh���N6sI�6m6�|�6��۶@k�5�%����,p]5 �4䀃6�8�|�V�8�.=�����5w� 6Hu~������s�@��r���ྶ���66)��P�26z�"���6
�50~���m@���B��w�6��w6�a��:1��g�7�⧶L@
56,�����4�55B��06��7;JD�Q��5�6��j5��"4P���b)����t�6�)T�2��5�\��W]0�S�7�lu�6d��6���6Dg6����H�L�D6�F�5<XB�	�h6&����6L�6�5v%@5�|j�"��6��ɴ��yZ�P�}6lµ5r���:{����$���+6��46�����ߵb�5�a�6��g�{-G6�#85�]����j�l�5LN�6x�x��ʶ��c]��W���7c5�<����i�������`����R6�5+�6��6�|���e4�}:�<��H�M�e�6l�(5l)���6l���*�%�6�Z˶��״���W�B6b�m���(��6�mU�u="5���F�a�6YĨ5]Զ�D6`�}5��6W�6H�	5�B6�}��^N����5��D6�̴����L#%6��
�(8V5�^o5�7����'ȶ�5��Tv��Z^�6t-��u%<�CD�Z˂��>�4������@�:�ȵ�\�6�����X-�JN�5�ͤ6[�p6�ƅ5dʶ��6Ix�V�P�l6�y�5ѩ46��c�i*5�ͱ���6�@��16�L0����z|6��6��t�y����6�X�������#�`�
4�/g6�27�䟵���#���D��*���3�.�@6H�F5���憶����8g6P�Y5s��5��~6L̂�f~���|6e��6�����6lBt����47c(5ԃ�64�M5(7d�W)���$6x�^5���4p��4n��dt�&O�L^���^6��4�������ڐ��RK�x�nzK6P��5 &4����4��_�.�3VZ�N5D�6|e�8�.��O����?6����;� x���E4���Ӯc��b�4U�4Y�6�<ٵ��y��{6*=�5Xm	���@����6��6��#�����6�錴J��6P�մ�����A6�gȵ��K��>�5��������96T�,�Oڮ���D���v��G�q����6&�6�CH4<^[�����.�����q�6�oH�6��)J7�r{���5v\��Й66�����f676�Yd�vÕ6�#	6-�A����6$G��N=��Z6��5��5���3T�6脶�P5؇���O�4��5zi�Zz6H�6Mĕ5A����G�6H�5Fࢶ����/��E�n6w]5 !��R�6��|��z�G\�H�+6��f���H�l�)�U�����5 g�����dD)�c�Ͷz�)���6z��5�Bi5��F6V��:+�����?��h��4�'�6��e�P�5��6
^05�;�� �5����u5�z6����9�5aV�\⊵��z6v�o� ^l�R���-��6]%�0��<�����,54�Z6��B�d�6Q��5�K15�XݵrQ^5�u6��>��E�Pߓ5��W5��l6�qg5͔�8H��.�Ƕ:=]6�';6�����rF���h5�к�����-����#,!6��Ƶ��`�E�~6��4*b��Q�ct�6x��&�5<��߬6���5���5�Q�5$�.5(��6�e*6.K55r!�4�@��<P���^6/�L���Y5��M7�qy60T��ކ��ۉ6���3�3��Kt�E>��z�2����5���U�3�é�E��v��i���d�]5&������xp�V������^��Ӓ4��@�d�;6���6�i�~��5ޔY�z����N0��T���H5�d��<fM5��)�֡���h4�"5�����*,���,����5�hC6kG6Ź5y)ⵉ����6�ܣ�pҴl����]U�b6+��(@�H�.6W]�������f���w�)H25�:��;�6P�+�4H�4q�Y�G�L�����i��2m�,��t�5����1���$g���6ά5�� �6sE���ɶ����%t6seӵZ+5�Ӯ5j� 6p�5��&�K5<�����
96�O6�e��`��X�6ÒI�QDε.;C5 �3x�5�96�"7� �D�jB/6 -Ĳ��P�
������5���G��6�ȴh���م666`��5P7p\3�3�6��ܶ8W���8�i��TDX6��6�#6��(��6���L�6��$6�S72!��7���> 6d��5��5ؔQ�Z���=�ܞ�6�\�6"������5`,�-U5��6�����,�69a6+��6w�4땶��H�G6�'7�ߵ-.����a�n�϶h���e��Jt�6U6 r�BWn5�/��ϼM6��Ȱ��X�B50^t��π5c��6ID��w���N�X�g�z�E5gՋ����nd6�.q6���5���5jON6x�"5 y���Ƶ�Y5
Ό���5C��JO;��0�5�>�8�f���6I�Ƶ�_���6��1���96������T7�'���/�����ڗ���O�5�]U���5	h�5Ѓ����6���6�!��hM%���E6L�5L-O���5�qĶ�
�6Æ��:lƶ-��6��g���,������LU4P�6���5ЈC����5��{60��4����}ʖ�*�U���1��6|�O��n��I��6J��6<nֶ Z޴�r+�����~�6���5T)µbQ�qzE�0��6�Z��B�6������6t��6�+6`Q��5T{����5v+�񪽵֒S�h>�5�Vö>W�5�6������6h�Ŵϟ63CI��4������	z6=G�5�쮳��E6���59��5�#5ڣ"5s�C5���5��6p���r�5^�	6l5��7�7���ߎ6Dm�� �6�7��.6H	�ng� �_�Z��6��5F3�6@/4ө�60�-7l��nv6X/�5�F6ޏ�5#,�5g��6�%��"p�5��5���6��6�P5f�k6��6{�64�5Œ���v�6��Z�g�Ĵ�C!��l��6��5{��4*��6�6�Z4 b�6�$y6�S��S6"�6L�,5�;q�P6�$���o%7������6�FͶ©v5z�7[ʻ5�34<�*���B��҈�6��6l��5$�ܶ.�3�p��6��(�3[�6Xq���"�4f=1��	�5��G��]�/F]��6�s6�����#~����{-66'�6񚷵ZO��6-�`Q���6�Ⱥ��o 5��㶴U�6���g����5|{�RL�4'͘6(_��J�#���Q�g����6���-?�� G���ʶ1	Ƶ��ʵ�yŵͷ�56ʌ63� ��/��#2�2^0�9j-6���J�$��J\-�p:��P$q6��p�6��}5�?��؂�Zc6�6GP�6��6�jZ�;
���P��Hj��� 5t���wб��!v54��6g6_��5�6_v#��k��+��6�+����4g��6+ԑ��T�6c���9���h6����E�6;ֺ6����0R6z�� �/1� ݵM����.�6WO ��ڶ����Mӵ(�6�	��֋N��k����5'B 6��5�o%���j6Y��45|׵D��6<B�� ﲶ�a�6 t�^e���,�!oP5+ l��V67�N����6�������s6ą�� :16����R��5�Q�RC�����5��̱��������F��w�6���^ �5F�t��р�N.%6LBv6F�~5����%6`C3�'��Y�5򽥵40�`��5��O�����B��Z�������5j��5l^6 ��1�)K��x�Ge�$��5�9o6ĉ��fB/5�Ƴ��{65��ϵ	s6��4z\߶��!���0�x�;�\3q4��ϵ�p���� �bӶ���5��4�ﯶ�U6I���n�&@A5�JB�߇��9�6ݍ�@u���3i5t�;��\�54���ט�6��5�`l��.�5T�O�XI�4^�6��[�04-3�Т6�/�4���6�
۶��16�i�(��5�6$&�6_6�5��S���6�m�6���6\������4�v6�-����6&Ƈ���,�7 ��5�Q�6��a6 �o6 �2Z7��X5�D�4z���脄5h>n�\`l��05`5�b��>��8ӵ����y �K�C��fg6�8�,��5_�6Z��6��5���5�*��?6�w���\7� ,�?v�5���5�����T�6>�x�����5���5���4�oj6�~���资(	6&9߶ڳ�})V��={6�2���K63�O�6��5��<�����,���u��6�0��6��6�6Da����뵾�35�+�<��r8�6d��5�O}6v�-�n_z�@�p6�']6����ƈg��C�6����ve��3��B6v�Q�)S6�d����56����K6�"��iN��A�5�"N�����`P�4�/�s�#6�'@6v ˵ S\6X����@�v7��(N�5 �1�1>�6��ĵ*���2�-6#Q�5���@��3h�5�5r��6(�6�aδ�ϸ� ��5�6Ҙ����7��v�l�>����5��5\�\��!�6�]h��S5�4p6���8����h�.O������ �/4T�g5�!-�al6i����9��v6 ��5�>R�ֻ5�ᶴ�6\�4�W6�
�5 �6��5cؚ����q�@����5��״lB�p�u�x�k6���4y��60ȇ��&5@�
4��
6��6)Jֶ�6�!��l*�&�B6���5�� 6�U�5�ٜ6�6 �36�����*��q�5)�
����5��4@b���ɑ�G�:6׳v��'�4��6ԑ7���*�D�5�p��6w�k5(���v�6l.��t����/T�L���\�5v$��'4��5i=�ٴ��&6е@m�@�A�����\t�5R"q��ק��9��[��������Q.<�dԈ�S���l����%�5�ł5>l�5+X������5���5@�q5���0'Ե��S5�H<6� ^�d6FN�4NҸ5d��2@�5{`5���4(���V�)�F��5�CG5 ,����4�>6�=U��&�5�D�@5D�36}5��Ȁ#5������
5�˾5U�k�K�����4�-L6��6�L��6��⺴��E�5@z(3ˆ���O6d�R6��M589�5x��-����5�d�Cx6�{۵n�$6���5�Ś5��]6XI�K���5&@5pLu6��5�=�}=�4��������6{�i����5�D�5p�\4	h�5F��5�঵���4�5ضH׀4 �G��&+��?�5����i���G�������5iP�N�ϵ��U���Q����6��*5~R�4�<�4.�h�eb5�S�x�F47�#�P��5j�T��=���|6����hy�5��t5[�a���;5���ݸM��? �ZM 6㣜��r��W�6��%5�˵fP61/	5�jq5��x5�4��,6����
��� ���[��b6�L*��4b��:z4�/ͳ�t6�hĵ�Z�����._j6��4��u�t;6�*�rsw6��6�ܴ��C�y8>61#��Ȁ���6^y!�3&���E������N6ߗ����x6�˟���9�n6V�4���4�ǎ����4��60O[�<�@6z]J�#�3�,��6�l�5��x/24w
����5��5�c��BFص�s	�N��5���v�#6�p��|`ٴH�>�p��5�����T5vw�5Hk��q�25��5vN5�J5�4_ ��,�5�	��&y�~���eʵ�n;�<9&4�|̵6��!��UE����5.�ٵ��'��ʓ5���8|ճ��Ե��#6���4�`I���5g_�E��vS�4�����\5���4-�$���õbu65��06Bl�6�R���3�4Ѯ�Ȍ[���e���o5h�=6��s���4&�5�M��x+e6�i��Cյt��4N�6k�h�4�6xL�51]�5�����N>6"v�����5��ʵY�H�X�G6��5א��Xa�3�Mٵ'2�X66�Ì��P5�#�εD����A�H�o�&��5n��v�:6�V�J"��B�D�`�6���6�4�5v��ƃQ5���hhb�k�6�n5�+Զ�@oV6ܙ���54�5~�4��5�	�P���f�`G�4��4���_-h�z���L�6n�j6�J���r�=5qG��o´K�B6x�(5��1���S�t<�X�3�XW��T��46^ҥ�-���3c����d�Pb24�L��5�'s�@�5�c]��%�6��5�����5���#o�6��5ۂ�G7a���6�ѵ�c��0�}�2�x��E���)�4hz4�GU5�q�5�Ꜷ�:ش���5�6đ6y� ��I/5��+6�*�|n?6#��6 �B����#������5q�6lك4�U!6�1�؊�4��е�
���m��a��������f6\���*6o �6g9)���5��6�I6�т5����l���"�hb���䕵Z��d��� �y��˵l���u%�U�06��CC6w1C��.�6Kζɘ5.�c�2�5$�5m��5�I�X޸4(�-6j� �H�3@�n4N�`�f]B���k6��a�P�?4"kL5ās6f6Ȭ�4p�괊�4�5Z��'=������0����q�	�4�1��[�5y�k6X��4f=� 9:�`Oֵv#����\6�6l5��Aw��-_���<6��O5@���#5H��5�ֶ�W��8-3�֒�S':6�?O�Y�6�-�5����s�5H��Q;3�z���&q���5���͵5)�4�>
6��;6P�*�[fȵ?��vb�B����ֵ�B���s'�%�R��м��6�
��6(��3�6$6`�4֒��|:5󚴸��5|������B邵2h�5h�ɴ�p�6��o6g�e6��"5,!F�Փj��K��@�5=y�5�ܺ5:D&�ٿ���ȓ4��X6p��46�M��7㵔gh6l#�x��4\b��ϧ5�>�㨍6���!16p�T5�ih� �U�D`6Fw5 L�0�X�}��t�56����P6~48;�4��/6`�ߵhc4dc1��yֵʭ6�I�5��5�08�� r�xC[5��ȴi��5�P�4�[�=�6�������Ը��_�P�Jn�5**뵜z5��,�y���壃��� �귗�kP��:�q�x[6�޸2��?�@�x4Y�85��v5��5n�ԵE�$�lo�5/�5�k�b6ŐW6ѾQ��`;6|}��X6Tɴ��T5D_�*�5�c4���6�Ը�9X6�J5,SF6��<�d���zH6zK6�� �t�R6#��0§���4�	��86���5f�!6}�'�H;��|HV�_���$�%��X��	=��!�6h�i��ܫ�.$l6�A��9�;k�6^�z�C�.6��6XL5����t�t�:�d�}6�~e5�Z�~��_��	�6*ݺ4�u��(H�4�|#6�&�5|u����?�̵V6Qd2�$��5g�3��x�4s�6R=����.�3E�����#���N6�yF��4P ����4(�k����6�U�7y��?��5����,b���6��54�絸�I5(6�5�6t�45��&5BU��Yǀ�O|m6}�?6ǀ6���p뫴\@���(6��߀�6_R�5q����58�5��[�����'�5�S6v�5 ό3�Ŗ4�$%���q�@ꓵ��^5�͑5�D�5�"���V?6��<2�5>J2���U�HP�5���6q���v��	_�����5����5����M�H��3�s!��n��|)��(�5��4��4���5t�����3�	@3F��6��m�H4
�ӵB8�5�6Ъ����ֵ�仵T�׳2�����W�6z�ܶ�B�zu��r��6�96V�^5Ui6����2�6�ߴ�aⵊa8��B
6��,�Kw6;��|]�5;��嫶��5p��3�5��	�*�&�zd'�cI6��6�,o����5�b�T�4g�ȵຄ6'Hw�����}��5��Ҵ	�5ơζ:.Z6-�6(�R���qE��Ke5�֘6�Z6<(76h���ѝ5�'���r^��BX7���6�d6v�w��&W�~��58{�5뛾6���\�60�L�z���	���W5��"��:˵[�)���6�O�6�pX��
�4��-6~�t5Y��6��<�e�40��5��6��X6@*�6��5R�5�Hm���J��X�3d�6ЭӶ |�2�4�6���5#dG6C@�:�,��К�Z��5�V��5d��$�4i�6���z���6FK�68	���T�sIm���B6bBѵi���,6oE6g�Ѷe𔶠�6-ڂ6��ɶh%R��Q�45F��cy͵��7XkE��kH����~Ҷʥ� �1�R�ӵ[�6 Y���ɚ4�^���n�!=�6M�¶:Ǆ5�\ѵ�(��6D��y��w�6��4����� 5lJ��^�vc5��H6�]m6�(�5�o9�<9�4��6���54���1^�6NH��`>�3z���K�]��6<�
7R1��6�5�նz��5��6��R�O��6A�5��Z6-��5<^���6��>~�6v�?6z�Ѷ�`6{�,�0�]6�B����X�Roi���6:ѵ7��wf�585w6�+3��eʶ4ġ���O�����^����j�6�M��Z��6Ãv6���+�F�~�����*��k�K7Z턶�yQ6;|7m#�5ZN�5Dv�5��̶�2���S����6G��v��5��J6�����w6A�?5����ヵ�W���k3|6���g�6������6n���(�~��}6`k���T���6F �JB��|�����?6��4p�^���P5�3�6
�����5��=6���6W.�5�,'6�B۵ �5z���[�5H����ý6ϛ6(�5r��5ж�,�~��6�yP6H͊���ݵ:����6��O����N6>�rP����X|���ue��G��@�ز�P�+��6�Gζ`�h4���6�l�6�J6�~��������ų�Z�5��W��g[�F��5�KI�-��5��
����5��`4�ɞ��XL6��.�ˎ�� ��z�7j���|k�5��]��z/a��8�6�	Ͷ���,�K��%���ح5\#�b��6�
��4'7X�$4l�u5$ �5!��5t�?����6Qn7�����϶ґ��Y4Z#Q���<4�S�6jbܵ�獶ĈX�F�w5v��5�*E��ҋ5N%���;5ƪ�6B�:6u��6 �����5 Vj�]g6B�6��I�N��5@��4�ZE�lW6���5�Ԑ6ҍ�g��6�\h6(Ȅ�?�5��5�y5N���๱�$?�5|鞴���W�+�0<b6H��t?��H�3E�6F�]��&�6�06؉��(Sb6��T6�:����6^�R6�zk�|��5�x���]c7�Ɇ�D��5�z���;�4��#6�|�af7�!6br~��n�!I�p�5x�j5�R�5��6�Sg4
[R6��5w$6��ɶ4��5'$�6���5���8��4@�9��`�6W�t5�� �����x5Z��5b벵{ 5�S6��6.���)�|^��S	;6EY6xݵ�2%���s6M|6�0b6����S-6�$N5�'��Į�6�[6plߴ��� ����M5 0ƴ�͌��4�6��������a6H%T�ī����5��.�d�+6`�n4@�˳�D'����5N�� ���6.�%��m�>g6�;x�	�65�!�5����O6J���̫��@�6��L6P7.6z��$G�6ˢ�<-D��H��3J5t.5�̶��/�,�Եt1�5�؅6��� 𢳘�.7�~�6�a�@�ȳ�~|���6�t���=_����5q�6(y�c��`f ���6�f�603:� ���5)4�5����`$����6.:���C���m 7������l5���O]����6lI;5f1�mL��.i�5!�@�P5��c��6f�7��1�5<۵ �\���F��<B�T\=6~)7436�ڇ���@����6	��F �6��5���(V�5L��6$}B�����̢ȵ[k6�� 7�Y6��Q�Ĝ�6��5
�I�J�
� -6�8���{��
&5'����R�5\(�4l�7�u��Jƒ�;囶���4Y_Զ`�6v�I���4����5�RB��<5,�66vJ�s���n�
7"�ɵ����x>�����R೶`�s��j�N�6��C�(��P�5��5�3��|	k�lT�5�uʴ������u6�t���Z5�rK4[oN�}z��\�)6���4nŵ��6��6����D�@�T�6�?�����6�P�4)82�$��5�ڵ��5�S(6� ����ѭ�5;�7��1�"��Pe^6������5;�5�I!���8��<6������[6�H���6���Hv6�S46І�60���:f��`8�xY�d�6���t����"�4�q5���$�3��x�2X��̡�\�"��5���4��Ҵ��Ŷ+jh6X��Ǹ5��7�N�6h6g�4q�6��5�����*tA7�ԵT`ٶ��h�2O�57̇6@��3�뢶��U6dB���oN6J%l6}�Me���
��A�b�6ڳ��,~���G"6/ŉ6��=����@c��]f�@E�4��6贫4"�"�bq�5������b��a�@Rm36�m�z�4���4��I�@��4$� � �C��b652͛6K̴�Z�5RA�5� �h�86H�6���/ؚ�J��5{�6�p6�cx�b�6��ʶ���9��5/ܶ4�6!����(����6�+&�t45��5!'�5^9&�s��6Hi�523�5���5��[6���5<O�5��+6�j6�����f�a�5o6��ƅ�5�FƵu�5���6�D5a럵��B6|��6�WI5�yE68����Et6�4���� �3gbq5Ba6�m� E6<��5�@�5On�P'-7n����t��k7��5 ��3�5S�Mă����Ho�|S��0����K�3�]���}��z1�6�F��p������6���3D�6��52��̂�6s/���/}5��6.�8���4ơ6��H5h�Ŷ��5� �4�u�p��5N-6P���r6p�ĵ nr�Ԅ6̃��a*T6mK�6qfX5I#��K66�6�R�6.چ5���ہ5v��5�j�5k�ڵ��+5L���п6�R�5���<����5Nu5Dy~6�� ��E5�GR�=zE6S�ɵ�.��C�J6Xv�/���S�bB�K55�4�5De����h5�f5
T6i~�4�sشj,�6��51Y	��H�6���5`�5��5�ؠ�a���RZ��}S�5�IT63�x(���R�6��5���6��*��O��V�� ��	!���C�8�����5Lř6N3W��z6�z�"��5����c558E�5�]���5 #��~&��ε��WF����̵���o�5����ִ�8V6�Xo�2���K�6ĶEI���4C8?�
�n6"]���4�n?5�0���M6�E��?�c��F���7<>�6p�׶��ݳ8f�5GL�6���6����6ʝ�	3j6��06�� ��]5���5<��44�6�϶3Rt6�6P]�5�̺��E���o���Y6�&6���4�U���6(x"4@� 6�c�6�A�����5+6^�G���N��涵@z���n�6���RE�5L�5�P�5�������:�5�'6�� ����5���4�_u��|x5D�5�JH6�����е�r+�=���^x�6F��݉�j��6�k)��ش���ʵ&:;�S��5�H$��gf���56�5R���NW�6�#�5�����v:j���K���	7N���)�V5@L�)���̑���6���H1ӳ��5�d�6@�4�����36-�7O�6�T���^`��L^54�'���76�v����&��@6`y�5ʞĶ��6�#�5��5Ћ��F~6Td7�i6�T�6�6��6���\H6ڬy62nn�:��6�޵�޷��v�4\7�2-�^6���P6Є�5�P~���6��r����/0 7�~�6�&ݵ7��6Lˎ6npg�����J�K5��5���RMb6�o�,�6�؏5&E�U���O<6�\��Dm60[�5˪m6��R62*ᶃ�a4����j�4��5�o6��6$�)5Pu��ep��_���<6J�.�T�5���6N�3�i�v�65L���58յ��h�P�4^^��N9�6т6��5 �04�3��J���6�v�^�S6u}6$aM���5XP��S�6�5��b}4e;6>�6h�5lj�6Lж��Ҷ���6|:�����34�6v梵h�����5(
�5yݶ$��5&���n6w26O�jU?�����l'P6�d�5�����	7]�5���PZ�5��V�V��6H��4�����\6-�A�ag�\}���&�5��6�e�x$�5�����Ͷ���5�6,\56)#�5Ln4�h+67^����w6���8Ĺ6�D`6�g�
W(�W(7l�q�����6ڤ����7�l���Z+5�B���Y7���� �������ĕ���B4����
Σ���s6�"�6T���_�6f}���B���I�v�/7(��5z��5���6 K}6�D�6 )m�>���;	��u06�ø5h�V�h�g����5�z�5U���?�5�260�g6>��4r�5 J�3�6��C���6���5
"J6�G��|Iҵ���6d�q�P�?6O�86��Z�p0�6x�6~|���6`�J4�Q2�>�c���"6LO�5 �6 ��4
�6u�B7<u���7q��5�[M6�Wo5��0���۵g0��E-��.�5��57��6!uZ6�Z�6B��6����`�(��6"��5x�ʶ������J���b��Ab6��7��Z�5��6��6 �m�-+7q�¶�*j���u7�k�҃6ܲN6(����C70����6���p:�6��5v��6<����e����5FPO�(�s5�k�5|�5\6�5�� �XH�5�Zs6���j9�5*��6$\��&�g�&6�4���.�2R"�ܨi�o�!6p矶2;��}������w�6 �����6�v'6�1�h1�6?*�5��`�W���:s7xFG5�I�4j�����m�q�6���7�_P���� �
��ʒ�>4�5���� �6�A��� ��B���<86&w�5Nv6��7i�l𵰙Ĵ�j;��O�� �6Hr��B#�F-�6@඼�o6��I��9�6�[,�`|���q�U�;6��S��x6D5�c6n⦵.�$��6�4b��3��|�a5�al��766|V�6�@�5��6e���w�ʶ�@�6m`]���6��� ��/��:5(��5�%5��	�LZ�5-�6~��6�����R��P�5��_6^e�6�
*6��,� {Գ.�B���)�6�mߵO��6�?��| Y6��F���'�"���F7�6@9�6 ����ض�^c6Ov��ȷ1����6�ǈ�c��6����#6^6o�6~kF6�`��m�6��Y5����)�6����|�j4��� �Q6��5�V�6��5����D�F�k������6!�Q��ռ65p>6�;7�AL6���5��(��, 5?�7�6���05�a0���� V1�?i�������7i��6P���+3�6��+�`ڸ�l��b+(��Ɩ6̝5��۵��5��@�`	�3p ��(�1� ����Ѧ6?pL��z�9K��5�x� �Ȳ��)�"����
�=t�5�~���x50�I5���5��g׶�G���˶6d�`��H�6,T�58'{����5 uٵRԦ��*]6�[05G6h�붾I%�"�5b�p6#5�o67��6��6�ݶ�!���6�nL6`��~�	5�Y��r6��Z���4�����m��l8+5D~q���ܶ�8նP�i5څ�5"��t�7�Z؂���7r�8�����O6tB6���6�ȵ��'���7N��*z;6"�)6���6=S�TT^5����gյG7��뢒6Y������r��5~Q��@���ؾ6��.5�ڶ�5�66���3�H4������6�Wӵݓ`6J�۵vĵkr
�<�6G��5��3����4䪵4�ô���6~��6�	6��/6a}�� ;�5y�e6(�m�0R��V��5�_6"NX��u�5/�5Z{ 5 �!�$�ߵt�M6���� �M�<h�6�*6p��4��Ե��5���py5�q	��&���z��/H����'�&��6c�C6@E�2ݥ[��1��x66ۜ������~4d�ݵ���2R공H�o�ԴB4��R6�Ҷ��K�J�.�柖� R0�k�6����<"/��U�6R26����%b��5��N6��6fg̵�gU��4�޴g����,4�,6@�6$����3"�T�6�6��Q��E��?�6��65�j6�'2�H��6?�����3�ڷ�4v�6��6Q�5����nȎ�v�<�Ə�6ԓ���ǵ`�y6$M�6@��S2�6B��6��6�����`ֶP���<l�5��5hԑ60q\�զ}��o?6lڼ6:f�54�5T󭵃��6j]6������J�h�ʹJ$6��p�5a��`i5�jv����6��Ƕ8�˵a`=64���/7��6��/5ĕ+���U5|6�6���������В�n[��/�6\zN�X�6�G�3P�r5��(�/6b���6��]1�����Hn,5奴/J�6�ߪ5:訶'�5�}�D��~J���@�`g56��6��#�h�5s�]���5�7-5w�δ#�&�|J+��t�'KZ6�y�5�l6NNG68��\�(J�5�'�5B���r\,��!7�Ō5 �6p?Դb���62r�5B�M��?s�A�N���68�Q�2}��͞5���7���6ꄀ�1����ҋ6zHE��X�6NW�$T5e|�5�8�6�U��#��5����6|�6�5�`�6���&�׶I�6`s��\77X.`6L�J55z��Oh��*�X����7�N6|�ʶ���K����k�´K��=s7���5>O|��l�k��W���ʩ6ME7_��7*֢6B��6����&(�5��	7r�����7Zc�6�ȳ���6��o�=$6Z��
��5Η@�$O�6 �9����5�C�6��6�����B�86�eߴ�ˡ�����u��6��5¯D7U�)Lw���m7�G�6�yݵ+�6S��6��6�̉5���6�37�b���Z���k7bԂ7������5�17/�?�D�E��T���55��6��?5w�6 at�Fw�6tJ�6�6�6��rߖ6�����W6(�u7o�
5�y�4��l���xw���FP�|LM��h�*3�5���z�5Y�>�X6�6�<.5$��܌�6���D���~6�g[���6d!Z�� 7��5#;�6$�@7N�����v���6HwI��le3`J35�'�6�m�k˶��W�A5C�2�6��6n�6����PL��R5`d�6�ϵ��f�X���@bU�XJܳ0!��j[7F��.@ʶ��J�5�j7��63+6��*6��6�l87��5�rj��$�*x�-v�0�n�U�6X36�# ������l7@�6�^��Za�6�d�6βC���6&s���4%?q7 n�2c�6�$�6j(7 O23� P�%؁�~Od�G����.6%2��k6ϸ�x�35T�����<����6�g��&-�����6V����[��Z��ya7�E�6����l�6�ǝ���G7PBQ��%�6�ȴ6�Ƕu�7�Z�H�5��6�K����ֶ���7��Ƶ�KD6p��4��S���z5��6l�5'���q67�7dc0�6�6��7}�
7���6�ڶa;�(|�4�Q�5$c=6��껤�@*�6 d�1\s��P��5���5� (7D��6`Ĵ$&5���T����5#�X7�j=���5�$2��.6H˹��`5�~��� |̳>Q3�^�k�|V�5�2.7����F,%�"ؖ�'X� ��5���6����hS�5���N�6�d#��*7n�[�;��6 ڬ6�bh5�c�ύ���W5��� 6�a���Y�6�5ɵR��5ipd�Z�5Ż�6�'5��?��E� A�>XE�Z5L��6b�6A�e�I7�D�S5>q�6L*6ڬ���y5r\6Rr\6��6�ߡ6�x�6h��h=�5x6w�
�A��6~��6���5p�56�w7J�<����V߶ؗ��J�6�*�6A��� �5��6����!�6�@3�����b3�3���76;�6��g��$�G H6PH!7oˍ7��A6C�5 ;4󣃵2�6�A7b<27ళ�(&�5H�:7�k������s��!6����:�7��7��S7���7����R�6Ɠ
6�:n6@5&��	6�� �aݼ��t�5�"�6���7D8�5�}6�Y\7�7ƒ��X6���,�6���6aF������7��}�i�����<��6��m7�o7�B�6

6ޑ7�{~������^�606[<O78Ue���17"���Un7|�~�ь�4�/X��U�5�l(��]���.7�9��>o6���596X��b�6E}76 }6��Ӵ�eJ6cA�6T�ö��F���4��4��K6�t�����5@rF�pL�5���`�
��7X6R��5GC6�_�5�O5��6P�y���6�W�62V�6n'�55g8�9ζ65��-��p@����6��6pʮ6���5���|̉����5���5)��6�0Ӵ!i�54�>����৵�O�6�2���V5�nx�΅5�f�6�<����6Bkﵜ�6k���)�4�5�������6x@F���ܶ{�M5`�6�̶�3��z���ʵ8�74�6v�
�lb϶a!46*b��Z��yp�践@Ib4��6�P�<nC6�!]58�u6�#7w�������MU�z���P4=�T{.��Z�6J|;6��6�ۊ�?�6�Er5;��X��6&�+6��B5�l6��o6��2��K�6�*�5Ԅ��x<��H6Tι��b���A'6SC-���K���n���z5�8S��c6̸�h*F�xY�6D.Y���ﵘ�5<c�5���� �������Q�c�f�TP�6��6&�XJ浉�
6cH6`��5�J��fc6���4؃�5�k66
�@'q4d'n6y��A>62 "��6J�+vY6�(� ����a�6�kw��#m5wV1��'7�i��>�j�p#k6w:6�����5	
x��������L���̶"6Q;���<v�XV����5L��6�'�6�69wm�긧��Q5$��tC86X��y����6�9��邶�K���5b�F6�쏵���5�]���%5j�K6�
6Z��F�=<����85��E� �_5|>��Xȑ4��U�l�{6�W_�P��0�r5��6�Yk� ��[�e�2�6lY�6�e�6!i˶r��5~m���e58n�4����&�@?���̖������Ɲ����(=�5_��͛Ӷ�a�6U_�6Ⱥ��(^�7L�6��������t�6,���!e�K��`�-�m�5�0����X�{����V�5��$5��ȶl�߇��l�5��d��f��4��൸�m6�Ef6�AA����6�6�J_���$�v �b�96�C��d����t:��ϣ�N痵6!��e#�6lKo6���4>'��(�!�&���8�47B��*cF��my�dyT�`'_5tB�5���4�-f4{<͵��55��5,�����E�b6 C5>�6?�$� I-3; 6R��5Hy(�p'
��W�5@�������~(�Rr��+��5V16x���'vy��~��3�?��������ɳ��S5^5xb�0jy�j螴0�w�j�������P��e������5�����6bC�5~8�(��5JŞ���W�#���Oo6���u͵�,�5th�58�t�2��50(E�ED+6�m5�Mo57��5�"q��V���-5���5j�M�DK�5�kʴ�'�5`�i�b��4 &�:d�5�!6��:5��pQ�4�&�5�y$�Pł6������5���5�wѵ�����5Lr���Z�42��4��5J�U6Rӯ5X��5�0s�a�6xw�5��5fX5�� 6
�5Ϥ5?85ظ��9=1�ۼ��5�,5�����5�[6J��5���C��Y�ՠ6�5����� *�֮��x�ٵ����2M�R�Q6���0	��ve�4>�5��
5����n��.�����5�6gH���(�G�4�6��6C��4 �4����q�4�5Nbn5T/�5YQ6i>����54+��6H��5�W4lx6� 4�R6H��5���6!�εS�P��5��5�#&�v�1�9ĵꦓ6�յ3L`6`�j4@�1�:B6�$6��E3P�I5���[n���26��5g��5@�ƳR��6�	6�|���H��5��y6���4��1�g��5�F5���W6)Q693��k�T�4�竵�6�Z6~�d6���yW��P
5���5,ີf<�5�&� ��2Ctߵr�6���5�e�ޟI�� �4g��5Je5�6�MJ5{�_�V� 6,�������������]�۵�t3�"ߵSc4GU	6��k4�-!�X���"��� 	���*5��ɴ�4�P��5p�34�ﾴ����a"��8�4*(�]�5�����#��R7�5�5L�_6K��5� &��jz5��U5O<�5�����7� ҄��E��Z����65[6("�5�H6�|A��<7�P�#6)	��Ԅ�j�� �3��6P��5��	5�Rm��jᵶ�p��n�5�gܵ�<%6�=����66��X��T���5fW��M���H�6U��5�5ȿ�4P�B� ��6L�W����Z5N9Z�+y��z5P�P��� ���ﴓ�G6���5H����6���4��!�����)6=}?5��6r��D����n��Y�d�*5<
5��6w���J��5�o��Uڅ6��>6��������6�K��\j3*K�6�ㄳl(�4oyI6]T�� �A���
�r����6:��5���4(�47�9)6ȏ06':*����6 6�u��㥵0ƒ��6,b&5&n�57�P�W�v�6&�ض���4v���4����6v%6�������:��"��6D�\5��J���ິ3�Җ���x����� ٤6��6Pπ��6��6v864Y�Ԍ��#<66�"��5Qr6/k��*�A�� 7Ϟ�~�̵H5��{�<���B��5*<s���5U�C6�,�ؘ�V�36ᓷ���M���m�޶�5#�I5|Z�5�Y�6�Q�<C�2u��`��/�K7���6qt9�ޞ�5)[6\�6RwԵ��5~Sr����4QL5N�+�0�H�.�f���}�`g"6Xs��c� ���e76M2��g�57%���o6y$���e6�kT4�-��^v�63Z�6|'���l6�=���36؁6�>�4�N�����*=6g�^/A��ɖ43	Y6������6�_��I9�/�ܒv���>6B�5��E������?5����p���Ӝ6u���=�3p~��1�ζ�6��P���O5�56<��~/�6����9�]6��.�����8�7�D:ǵub�,`���k�ƻ56l��6�6!6���H�f��r�5�}W����FJ6��8g��ys��6�P�5����7�_��54���ā��I8�Gr7��ح4��̴"�5�B��G��h�6 ���ê5,5���5 ��<��Bl�TöaI86�57���������t�5�H(�|��6ԭ��D�)���l����A�D��T���'��8|�C���	56���"�/5�~V�x�a6$�.5���5Һ���֪��X��P&x6}����@����4'f�4Bf�5@>�5ޮ60��UµZ�X5H(S6Ȃ6IZ��/�������z66�Զ��D�嬚����N�6���5#�5!76P��4�ʵkZĴ��5��d�w5�Yy6t���/��s�5�am��ɵ�k
6ʭ��b��6 Q��[5�����6�O�4��4��3�2�6P��5�L~�2�b�wG�6�N�6���5��6n6��z��{5���5��W���H6xĂ4�d`6�5tJ��� ��ģ44ȥ6H�i5k�K����a��ى�Lm����6`j6�̥�{3c� ��5JW%5��6��2��Թ5/<o5�����6�#>4SⵢlY��<ѵ�����J �Դj6Y��ݬP��w6?�96�)6�?�5B������4� 4`P���q�6Ҷ`���h�.6�������6���5P>�49�)6���s+.6��(6��zJ�4��W��7����5���5d�Q��-���2�5zE�����|d%������A�(v6˫5:±��*7� C�3�����Ģ���|�&8�5�����{,�6�6'*��(�6[K�6�E�\�x�L��4�PT6�γ���6*1�5⎵��v�0�5N.&6�����-6�� �pO�4�4�5�g��D76����Ā �Z��5�+���E4#�6��N5NN�;6�T6���̸5�S6?8ĵ�^��갵F�(���b6zɵ�9õX��6P�4��1�>M�5p��4��#6DH��ԸԴ������>50V4y�5\�5�L4��j6 L�5n(6	�6���^6�w����d��x��n�5�� ��_5� 
Ĵ��O7�6��4 K���ɶI��Z�R6�8�>�Q�t�I6��	��?�3���5����^�Ե��6�6�6�C[���n�(Z�����|�޵��2�lt&��I�5�ro65S��R�x���~�/6p'��Cv6��=�<}��}�4�H5�|��b�6�M�Ro�5��~6`L������N�b��4�|6M�@��7�� ��᜴�i�$���ص]�����@���ə6ܺ6&��V)3��5x;�N�$6���4<�86\�L����R ���s��=7Lj��G���ޛ�M�s�M��]S6�ی6�'3��r���ն ��4$�7�ǈ�7/��2ⵠG5�����0��)��M�ئ�5 �y6F-6����>5���4� 7�R��Y�֚��D��5]V�a�C�s�5J�.6@��5��
��9�ZR62�5���50��6�SH50k<�:[��F-6HM�4 �V���Z����6�n�5�oնHU���~5��5��sz�5�
I6�Ճ��\��@\^6ʕ	��<�5�Y�6�8� �	6�	�c�����6��B�G�D�b�X�<�$� ��3���en��9�4���5�u赚յe�6iU�6uٜ6D�E6?��*J�4��66X"�5�c��Q�59��6�A66�JJ5"�����9�5� ��ж�pm�� ��xԁ�:2�0$�5�60n��A
� ��21p��� 5Ұ96d�6���/6�:;6s�ĵx�0�h9�5`+Y�*&i��_�6( 60E.5���6@��3�Yi4�瀶 (H2ҡ\6;z���}�6Ԟ�4E��6��16 !��xZ�Gs���u�6��"6�����35Ka�֌���b� $=��Ő6c�6h.58w16��5�>6$|V5cI��.w 79V��6h��B�5�d2�8��5B~�6�o-6RG�6d�Ҷ�cC��cL6 f3���6KX�5JN-���6����N�6@��6*�����D��4�y6��
�.,Ӷ�sd��e����B6p���/�i52�H����4�i�4�54���4���n��]�������ZD���H��G��(ٸ5������6�	4���Jc�5:/�4�B�%�Q�?c:�+孵h9�4�܁�rӿ���ٴW�4�~�4��l5�с5$}�5�*e5���ꀠ6��<���*�n�6��4�f]4��4���6s��6���4���5O�5��4x열�j�6�`�6�F�X
�6�"��Nɵ��k6*�� Y4�
 6p��4<���$ֵRK�6�_��\��4 �Z5�ƴP�����l����A4~6�&������/6>�6X�Դ H�0�ǵ6�6�G��ʶ>6�6�5�*����5��5)-6�_|��'�A%�5M���5�����S=�h}����ö#��5�z�6��4x&85������ Kѳ�*���Pg�h��6|M�5 ^~��n6Z�62u�-�J�g6�t���L5d76Sa 6U�6,gg�`Y���	6k2��^05��{G�5��5 -&����N�}5Kc6�����^��S6�6���4_Z6jm6���6%	�����6h0w5� 44�=�hLd� �%6s��5ƪ�*f6DB6dk'6�������ҋ��OD6KP��3!��w��d
M5p7����5T��3 E��P�ȧܴ��4��ȵ���4(�S5N�5t�:�M�6P���& �S���\�6B�=6�C�5,S\�(86�5
6���"�W�	��5�ӟ5�`��"2��軖4o� 6D_���s)�V��q6f�׵0]4�,�6�5�j@���/�	�H6�L4X{
�
\|�E�5���5�c�Gױ5���>:��&'�n���W�LW�6
Ah��iv�!5_�k6Dy!4�Z;��Yl5#5���{4��u6��65w(%6������a5ȶL�v�ߵn�Q��P���5�0|�,���j�5�;F�A�-��<6�r_�B�W6��c�ƛ���Ť�_��Th36B1���؁�d!ƶ�Ⱦ��1�5:I���+,���5 F��
b6����9�����4S��nNw�H�r�Z�z�]��_7�R��Bs6��B����6�x6�"�5F�x�׶�A��ڿG6@��4}-��ܜ��`�4j�z��6#�!6+�zR�6%Y���J��h�!�S�6 0p�^́�`+��>������6���D35�XE4Z!���D
�׸U�ľ^7���6�Lb6�_�52�6n_��tr�6,V76��(��$�˶��X�@��3�~�6Of	6x��5����4�
����ީ6�况��_�~+���A�6�-7�g�z��6H��5�!
��ê��6<�S5��� '����&���(7��z؆6���h�6�g޵�˶L�7�*��?�v���$7��-7���w�����6�(7��6�e���_�{�(6i������ӂA5h�0��in���M6L8�4��58��5�s���5��4foε�YL�zӊ����5I�1�H	s5N�k��7���N)5T���p�7��N��|�5�/�6��ȶH1/����6`��4l'��k�#�7�6�!5@E2,w�5<65���g��6�ˠ6C6�6>=R�>u?6�e�B~�5�y��6�pZ��ɵ�9�̕�&���87$�L�����e�A�6x��5��j6�li6�]����U�YV������~���:�%�� �0�b¶`��4�V�����b�(6T�O��H�4�FS������6h� ��+\6�|A�8�.6�l;�����*���z5����G����6t>L��F�6���6XI�h�u���,��:2�I&���E�6�D(�Ao��R7�6\5L�76���5@��6�����0V�5�?6Z���6xvڶ4�l6�+����5�*���Ե�Ӭ������7P�4�߾��Y�68`-����2��)�y�}���5��6���� !3̵���6!�6`]3���"�7V�5�=�5�n5Z����ͷ6N�r��r��I�ܥ_�,صߴQ�3����6�@m5�,�}�6XZF��ŵ~Ѷ;7)���A8�6c�F=��5.6؊ɵ��n4\��5��%���趂.d6D��}�o�^Z��E�5��ɶ��{�gB�6ϓo7*}�6I�2���!����ܔ�V+�6j�O�\g���� 7t�B������6���5n��$�ε� �5$䲵2�7��&6 l�6�fC���:6�(�5hi5(5�&�^�������8��XA�d9�����6�@�L�6��5��L���5t=��wx<6���4�6	���ٳ�������
�����6��h6k���66�Tn�l���J�-5��5\�O6��i�KWZ�L|�6�,����4�)6�e�6-?�5�#�5|�7Ԯ5*j�5w-6�U\�8R�6��Q6�t�ո�6���6��Ӵ8�1�+��D8�5{f 7��5P6#�6>�Ѷ@��o��6�+���}�;z6�>3�6��P5N����@L6��x4��q5~u$5��O7���6�u�6|Q�6Pb�:��6̶�۹�rہ��
����6�ό5`�6��0���}��j�70z�6v�����DR�#�"6FM������ߵ�V
6�,!���v6�f5 �嶊��5 0b�h�7�ڴ~y6h��4�k7A(	�	�ʶL\�5��ܶ�"�I��*٘6s�6���4��2w6��Y�r�6�%7D�6r�5�<��D�%7y���`�Q5$�M6��4���4̩�6&O�6h���K�5�� �U�&��	ڶ,�����6ޏ�Nh����%�6����6�>	�������6h7�5L��6��4o�b�D�>5q�v�~���D�]�����|Ԍ5�{�y�6��65� 7�2���V�h�ߵ"�5��6���n��5�`�������NT�KΪ6e�6K5�Ӂ5Z�P� Ge2L�6��U��_[�0K����5X�5��� l02��5T�5��#�ZU�5ڛ�5~�5dTR5G<���5>>�4��%��5�5�Ԫ�^h�� �����a�̈́;��"�6(����5<o5�C��N6�a�����©���L�5��ݴ��.6z�赙_�5���.P����5�g�5�F�4�� 6��F�h����E�6NѵN����5�\�6op�5H{^5����;"39�6��@5;9�����<g6"3r4"�#�]��f�%�x~4��3!Y��{��������%
���'61"����/gu���G�}Q3����o�6M�����5Fv����w���ݳ�~ӳ��N���w5-ڛ�R�l6�!�"�����5����0�5��C����6��2
����z5��5��5���	�q�Ҵ�4��z�KJ�4�d�	�g6����g�5N�4PR;6�N�<2T���5f�5ȸ��SQg5�2q5P6A�$�4L�5b�6T��ʣ��Z�t;���0���r憵]'6&���:���6��60��5dv6���fy�`�Y֞4��γ��50����A�b�>6r���<�|�޶6�T�6"�H��%�R�0� )�� 759�5H:��*��؅5~V?�ϕ��@���F��<� ��
'6j��(�ȵ��
�XW���>5�W�$Ɂ���o�ͭ���C�6[ &���56�`5n�����!��ld6�Q�3ڣ߶�@Q4T�6MH���W��z�5������#5h&#���b6�/+�����E�Ǻ�5b�6���4��5�}�~��5{�Z���%c6J�(6�#��م5ȣK����4@���+ÿ�	�o��>B�����/����5}9����s�K��t�㵩�絜�_6��5X�6�O5��s����5潋�H��4R�/�R��4��5��56���l#l5  ���6�f�DV5��4R���"��b�6h���!k6��z5`t ��6v�5X(e4j/O��i������&�5��:� qp�Y��'���hK�Cq�tr�n��6k�Ŵ@�c��6÷�5n�5Xa�����y���^�5h�l5��6���5���6̭H6���4.�4�pJϵp�4��)6[�5���3�X�2m5��5��I5�/�[��6�c�jO���3�����p� ]6x�W5�v;��)E���t4`>ճ����4����͵R����v��ً� ;G�:ז6P�3�E�5�����6��41kW�萟��VL5�׋���5��<68�6"��52�����95�@��"�5� Q5��k���6����$�47��5��5����606��3�6���5�X06��c��c�М�4� ��M6h�p4�������<@�1�f6��6���4�8�5Vj��?F%��6逵^$Ƶ$j)���5�%���
?��õB��L�=������5���4�*�5���z�5���ng����6x`2�~ E��(6����qt����=l>6��6�%ܵ�k�f'�5�� ���S���#�;�����@���(����况�b�p�'���4<ğ��6E�C��6f6�Ȅ͵0>�����x��(2����a��3)��H�����6
׼���6�5t�6S�Z�5@��� H2F�g5����f,���4�V��5t?�x�6����)U6`��5��6�������4_�׵�i�5@E3j#��.��F/�5�J��pz�@��3�]6�64�Bӵ���5�n�3*<5P"6�v�5�� ��=;�M6�lB4��O5g�:�����,���M6� 5�����咵(ί4��B�.2�5�I�5Q� �Ƣ15v9��W5�w"�r(����6c�6�%�6�9�(�l4dy�4�������?=s�
��4�ӊ����fE6rJ�"fF6�o�5��5��4��1���ሶ���m�<�O��x���]6�l�%6���4��6G�M�4L�6��5�Id��[6(O�ȈS6��56p��5��=��m�3):ŵhQ��c�6�A��@8�U�65[�6�+�4���5��ߵ�hq6|m75B�5���6(,Ӵ_�����3���5�/�5p�6�i��on���J6|xU6邦��<6�6�״�6n&�5H�9��76��L2����¥�6���j�V6�!� O 6�r����5̴�54��X��6\C�4���k��6�Ul6�M���&�T��G76�F�6X��5�*W�u/4�t���ɝ�hX�6tyڵh`+6!⸵�v3�ﶓ��5]�x5���4p�5;D�5��ƴ�!&5�(z�@O8���ص+x6�\6��)5�l�5�c���	5�rD6gd!6VҒ5fp�5�	��>��5@*�5��&6��	�3� 6>�ε,d�5g�;6\��@�6z�D��5�f!6����f6v��5��H��|��Q\�6:��5\�&�������;5Dj���h6�5{����E4�N��'��5��5"u���c5pT��HV�H`���4�Rش8�5�[�6a��6<�5�M�6Z�B��h�5�k6_��6l��6�&6�OG4�/]6���5�-`5f�5G�
��+6�#,���J5�/�6���<�J6`X^����ܡ�|f�5 ��SE��̩6$��5�d�6��06`W=�8�s6ܧ�6�׵��,���h��vڵ���5���-_����6�����?���d.�5t/f6���6�[6&�5`5>4�M6�5�s�6�e6���6\�}6X��6�x��^�6���4j5��ӵ��J�.2�6]v5���5,׫���-6f�N�X�5�h
6�!���K6zŊ���5�L6��5����҄58�5�+���޵W�06@m��m�5J��� ��aq6�I*5^���#%������� ���� 5�C"6�z'�$���UT4 a}��ɕ��������#-5���5Dk�4�w&�7;�5 *3�޵5o�5����~�h3�4 ��2����P�i� )� ��2�/J�6�!5?{�6��5��X�gC��� 6$ì����,�6��6� F5����i�@�(��w6߃�5��۶WQ6r?6@I4{-е5H���ζ��f��.6�gG�4;,��j��I�s� �jv>6"�%6x� 4�oq6%Xh6��F7`z6�01�5�5�,/�6f���˶�7D@�6�D��Hp��5���5�f6�$�6H"�5�ӎ6�7#�nöPN-7_�E���|��5�r�6A�5D��6��5��Rc�5����O�z��R9U�?�5BX5�1�tM5}���Iu6u`�$�5�_��kz���1�6��5-�嶾A?6���6VWٵw��5�&��
�<6b���B�6p	i���5�;�6/r$��r86��U��{
5�<�50ʅ3�Zd5d�6���q�5J���� ��>6���5�y�6R_�6�655���tO����;٤6@Ƕv^6��5�^5l�6���5�X=68[ڵ��鶵��5�6�C�6�]^�$N��&�46`������5�����������+y4!86�H� �"�^�6M�6®A7����0�}�2m¶�⭶hm��Lb6�얶���� ��^v4l��PH6�5��2�8�J6+KH6��?������jI6��v��,�6��h6f�
�P���j�ض<�r6	��6xN<�j�S���K����5�ة6��5��B������r+A��t��5�*㶃�f5,�5ir�6l��5�6����v6��K�ʚh��똶�H5���3p^:��R6B�6�t6����TM�4�������6P}�53��lr�B��٭Ƶ;z�6a
o6�γRF���	7C�$��I굀�]��Z�pB5��5��5���EJ6�����l�\��56���ԙ�5�tN�3*~6��6IU�6h,^6O���-�\6��#�K�6�Ӷ���38|��|X�6Dt�6ΞY�H��5"��9e�6�:7��u��ʋ6�r6�)S6^X�6�	6��5��z�%�6��6�����6>���җ�^��6⮣6�)ǵ�A�6���6�55^�6�@��dĶ���o�+Q����6.4�K�4D�yA�5x僶�=	6x/T��7�钶g�=6�:6Z�� �h�����6ɼ�6��U6OM6g!i���!7V|6�67�0�5ǋ6
u��T��6ڪ+6dԴ�H�.�]��"X����C68Kk68��ȃ9� V!2Ԫ߶��96La>6� ��֩�6�)�ȷ���%W�Z�;6�p56<�4��D�+J��^��7�������;6M�:��6�G����6��50��44�j��G�6�����Ƕ���U*6q'�6B��<����f�P,	6ҟ
623�5$��6p�;61�6�\��&��B��6��H�h�5A���|v�3o�5lm6��赲݋6.�ܶR�6�`6��>�<�.� n����4%|��Z$05�Hm6��d�v����w���@�6�?����(r� �I6��5��6/z16D����l�5��6j`��Fց6�T�6��X��7�5=�@�0I�5�:,7n˜��8�68r �\�6:![�'�ඎ�}_���,��8����ݵ[Ƅ����f���.q���-6�P5��6(65 ����:s7w���
��M��������6�~���:S���Ƕ�t�6<3��GV�q�$���U�%q�c�7��M5 a6���4���60*�4FW6֙6	�5�,6�H5������5Z�>���4�)|5��B-7hS���ˤ���Ƕ!��6���6u7�>v4���>z�J!�s����ֵ��6�̢4RU�6o�6�����ҵ ���5ʶ��d6����X/ �\�6��嶫�59���Y��y��p��I���V߶��}�L�ݶq#�6n��6�7��e��P\����R���6��'���)� ����oӶ������6H*�5��z6�K>�<�m��4��r8���D65���j2��4��g���J���ٶ{��`�7>P)� A��I��.��5.����b��k��>��6� �6ڭC�*&�6�}�6'�5���6ֳ6�s���]ɶ�7����T{����e6�V'��C�6��\�6����8/X�̋�6S^�6�e��0ɴ�J	�`��n�96Ղ6�6�:�'6�!:����6=z��Ņ4щ�6�͕�$Z�.�7p��6����Z"7`���?�5ܜ%6$���4ȫ��]�5j�5��Q�6�i�6Kn�6";�5TTP6��R��6���!���>����6���6,���������6�h7�G�ڱ�6D/�HN6�@5�6����!�$5��d7�f�6p.�U Y��_���c7���!7�N6��F�t�ԶR�ڶ2�ɶF�p��7�8�6+v6�cN��D��t�)�ȵ�m��}d���m6~�+�6�'*�亜5@��6���5:'���>8��U27�y����R4��+�ԱZ6�H�6� �C"���g�:R7��k���`���}�p�4.��6�3N�E�hv�5Ժ�6�;���7�g�51@)���6�����m�7�����$��SʶB>���6/ݩ���7�[�5&|�� �6��*7�֙�>��5�E�6�U5�s8��.9��!��$�d6|k�P��4�j�5���6"�87�8�4��5�R6TA���g�6?S69�k7��7!C 5���5!��r�!7���3�ڴg�ζ�l<7�+!5l����!�];6�q鵄�#6�Ͷ������6`D��B�6��u� g4�冶 ����65ಶ85��T�����4�!���7@sQ6������6���z���"�6�{�6 8���6�����鶰�4P¯������6 ~�����6�y�4g}K6�w7��
�6�*���lz6����'����7�\Y6��6��7� �L��6Y�6��6��6j�6���5������%�=�6Е��\i�W��R��5݆[�yXi�0hY4���6�O6L�� S45��x� 5�!����x<]6ȣ�5�ֵල�Zw��x�5��15P�{5e�H�5Z*�6$�)�4T06��s��6R�O5S���H�R�l����㵵"�5��5����$\46���6L��56n^5��6���0���세��vW68d�d$z�$ʴ! &�V��6�{���g�5>�/6S���d�\���؝��h�+5�C��r��
卵�^�4��j6<�5#�˶+/*���6��F5Pg�4 	��ϳ�&�3,����w�DJU5o�C6H6��;�8x����6�B6*�<6����	�ѵt)��'���)Aa40��5 §�Ncu6R/6��ƶ1�-6����re6�{3�B5H�T�P�4��4`��3��I5�X2� ��3�U=��kH5�.(�rƘ6���6�.R6�5��5�J4$L6)ڍ����v�6Z9εB��5���6@����e(6��6u��z�5�6t+���4�����$�6�������5/��W��`>�3���r�'7���6�5�G`6 �3./�g��v�5��ϵ�ڗ6�t�������z6�y75��6Y��jY��3��Ҷ*�57Z:�6XEҵۙ�5�b~6(T56��w6��5����H�|5�������Ͱ��˶^��5p�4��ɶ�`�6����da���xs�N�e6�R����|6�2�5��ɶ��(�� ����5>d�6Xp{���N6s��5f��6DEp�+@(�pDn6�S��y���w&�$���?5�ڒ����_
� LB6���6$c���B4ԏ��Tu����2�ef5�"���>�jć6������v6~�;�?�(6: 26��-5�}6?� ���5����N��Q`�6kv|��6�s�Wn����6<���Y�W���<j�5�6$T��r�6��6Q�6�.�]�e6��5D�6�C�6`+۳��b��Z6XE����c5�my��T��D�6�{?5`�4�5<���ݵ�5��O��c�6��(��Թ4Ԑ*� ���z/�5P<��'A-����5͗Z6��l��<3��(��
#5�`�|6�Ê5�6N$6\ E�6��ܚ6�Ƶ�6)'�5�n�5f�Y5����Ɂ�6�[���5�0�57���2��Ǒ5�ؗ���`6��K��ε��#���!��&϶����5Q��Ț� B%�����B6���5X�ϵ(�5H
��p���[�I76@+Q3!�4�n3�tI�5�|�65�&���5B�_���:���o��V����6��´�5:5v��g�5���^6�)�6t��54��5�˴�r�5��0�Y����ֺյ� T6�x��@��|�k6�!3�@��5��l6З�4g���d�-lB5������W�-͵��	�����!�3P���L�6��}��$�5�d.6@�Y5���5�6{5Zy�5�ڊ��
?��¶~�6R,��8b��ާ4��+6U �6g(6
�6fv���}��o�5T�6��b���k�깳�$�ص �5V�U��� �Z��a)�����f�5t��M!6T�'�Ct6���!�L��k�E��Ү�>��5t��5�
��ʜ�5(ײ4T�H5}�g5���6�w:5�PU��[6P ���ҵ��5�-�S4�5�<��
1۴��5�86J��b2?�s�44U6$46������50CεF��D66@GB4JR/�Ȳܵ`ĵ
A,6i׸�p�4 V� ����􋴒����q���6&[�~��6�q4�6ȵB�6J���h��5��x����60y8���)�L�<�z�"5�7�6��6��1Y4r���)e���ŵ�s�^�#��5��6�p5���P&�4kP��̯5��6��6 L��&�v�Ot�0Q4g76��ֳ�{6����%�c6a�� �q3��Ѵ�6�ӵ��R5��5��5���5�m�6��6��D�X�e6�ԑ5�������8և�D �4���5��ᵑw�5�t�4T��5�R�\C5��8��5@G4��h��TM5y�$6ηL6(��\��4��"54�4 QB6��)6 �͵�둵�m&���5�p51�X��O����6:&�5K��5����rM�5ݟ���K76@��3�d6<)[�3ɫ5��5C7��t�'6p�Q3��t6;�;5�
60x�4��Q� ���:�xsN6�C����h�*47V6��5 =I5��@�O4t��5(�6��=� p��� 6�y�5�L6�3��K6�5��4@��3�ז3�K5\7�5��]�8��5���,^��6���~�5�H6f�6��i��9�d���6л6�)#6_��6t����*6���51E;���\h��`6�4��Q��58N�p7�5h��r���B6�5a����5��ӵ쟵8J�4 �~�;�5��66�贜XN���5;�6���a�(����3v�����4�m!���"��5>=��?��a50Հ4�~6���4 ��2�L�"����[�5p�4��}536X�5��i6'I�5|9�}�D6����ٵ朥5��U��_�5X1��w���4P�5nUS�״�6Ȉ��zC��`i"��*6gi�5Fb����6�H˵��6Bw�5�(60�� 7"]��P�L�11H�bp��$�f�3�!΀�@*�3��C6�9���<T5W�Q6Ny�չ�6��6p^;4@�*4鮞�r7�6�f��lz�6x�9���5L�X5�O����.��6|2�5����Z�-6��e�@y6���-�D�X6�jҵ3B�5>d5t��5D���l��r�5�~��(֕��ꐵLu�6�[;6~�����6���3�W�@��3 �M��r6�� 6�g6��86�5p�4�#�5B�6`?5�Z;�څ����ε�5��`��Tߗ6O)�$K�5�f�5"B˵mF�5��,�5`r35}��5-�6��4�
���$&6�/�4��42F�5 �$�#�"�V`��x���.��ί���5 �������5���K�5;/H���6�A�������Օ��?����	5�嵦����@�*�6�5��be�F .5�)�6~�6$�_5)����_\6 h0tx�5 �.3��n�t�
�X��
�$��4ڕ5謽4�T��▫�Rk5�E��x�5uk��a�"4rÕ5��6L5nb���lõ0�'6�|6�	�d���f��5`Em�(�Q���Q��&�a��6N�}5 /ԲWo��G:���>�5N|p��M�5�;�5����Nj4'|5 ��2l�5��&� (�2��5)��5�[���n5 �<���k���紐��5M�S5�N�5��5����@5�Î��@U6���p�3��5�Q��0��4ޮ5�jϵ�d��p����@�4�}�4Z�3�`�Pw!5~�������G.��j�5 0��P�ﵺ˴P!�+�&5����{��51��5����5@z���ɵ�hG5ki ��T&��[�-?6��+���5�Z�A���5`u`5�	6l�4����f�5��F��i�6 ��3h?2547&5V�XB66��ֵ��4.�6�6��b6o,�����w��!x�|�d�r��p�U6�X�4�w�5�e����5��5'%Ҵ�9����6 *23p0˴��C5^�.6�g����s�)W�d�I5�WR6�En��C�PĦ4;Uq5�-8�|�=50�4n'�9I�5 xɳ�:�~M6�m�5x��&085ĥE��y���<6�]�4�N�-N!6��X´&B���Z��G��ؠ6�j��;f�4%�5~?f��O��TΆ5(\��p��/��tf赈T�NTS58$-5`�H5x�5@�������
�F�5�+�46K�d���Ȭ�4 �Z��1�5��5(��J���0")� �³�s��ӌ�5�5e�52�6Ğ5|�:� 1l3]�4��.5��j���x��+�4���5�����>ԴN���F���!�NA�5]�6p�60565��8�)6l��5,I��ڷq�X�5�Z���V&4��6v�6l���|k�62�56��q6FRs6�<阵�}µ<:;�/C5%T��R8ж�g�n��5�|6̅���_64��v⬵���]ߵ`F�6	�6S1�5X$5"��5T�6[4.�@4��9)t���5vM�'�ȵnÌ��4)6��7��i���ag6֔I6H}���G�5�k���<5���5|���d,�4 g6��L6C�$6 M��QL�s�"6�~�5��5�� �]��Y6��5~�s4v�˵�p��@'�3����-�i5vIo6#ն���/64�)�@�[��J�,��5��ƴ�ma6i�.�I�v��J>�O�6�`��x��r
�6ͽ��v�6hi ����FX�5P58A@�"2s�7o�5VU6316�l�4.����6B��M�3p�ʴ|[k6����Z�A6�:ܵ��/���50r��㰸���4XE�XN�����51�6Ƕ5nU�5�0���N6�E���5k6��q50"���s7�R�5�y���ݵ�9 6����d6:$�5�f5<:�4�b��-$6��0��Hĵ庵b����S�6
�b�yV�6�6�5Z�5�4��Yo5���P�[6�l$5<�5T�a�0�Ҷ�>�6��5%�6�����ؚ�\�L�� >6�]a5n@ɵޗ�6�xV63��WK�Ĭ6�������)ɶpqy����46�n�5/L����5��U���޴��*�PX!6B��>�t� �.���55��д�I4��X5�R��Ed�&s�LF5lj60I6���5��d6�Qi5tr���S���յ�#���ZW��3��3���]6cB6�M��L=��z6�W6~R����5(R5��s6̇>���D6\������#��x$�@�6��6���8F6|���f6T����6���5����L6����8�5���Ll�5��3�N� Z����:7l����A6DMz6hTO��A5�[�6!�Q�7�-��z�,A��B�6��$5�y	5@*�4��=�`6�H�43+�:@�5p5��H�5���6��>7�2��=QǶ�C�3�JY��������������� 5��H���8�6v%�6����;G ���1�����vƶ\j�6*5u6���`*6�Eݶ�"�6߾M�c��6���5�CL���26�݂6�N��j�7�x(7�s���M�6����ۣ� [6.��6�*��M�"��e���5�f	7`?*��4�aҶ3$7����8Q	6 86�Y�6���� U��|ȶba�5��4���⪟6>|=6X�5r�T?�Y�)�N�7�6ht5"	����M�$ݡ�=�%7�x)7y��a�46r�	�,�6��/���J6���Z�7��34ȩ�4Ձ�!�2���$6��56H!��P#������a7o�5���ag�6*�:6��gg�������5!7��ն�x57�3� ��6��g7�5U,�6��.�rC�:��5�d��6ȘֶO4���n#7�_�5�����!6����G�6H�7}�6�6X�t��#��Y.7�m�6 1!�&W��B��6����$16����T5(�j�t_'6 �-���~�"�27h,/7�T�6zr߶0z�����6�m7CUͶ��6�]���)���/6�rB����DNе>�X6/�����Jww6*��6�H<6'B��6���]c��?�Z�ֵ�k?���6�����K�6N��JL 7������6(�6�!��,�57���6��6ζ DX7�1D��[�5Vj7�l��\�����4�6�o7�2���W��q6//��v(� +��q	7���6��-5>Q�6�#%6^.,��@��L�6|yõr/�5*3�5t�Ѷ�]5�����&��6���6���ػ@�U�q���k�z6Z ���6�5���5>�06�Y�4��Z��������}�6:o6|��5j�6,��6��"�Ls��:^6��p�Kz�4.�"������ꌴ��b62�V6�*m50%5��6�t�M���5\�B���̻6���톓6r�6;���e6��ڵ@��6���7,6��Q�À�6�\>6�� 4�d65`�6<'�6�>�6���6@�n	o6���6�_o�*.�$/�5 �6
D�5ة�5��6�M�5{0	��6,�o�胺69%@6<�4 6��h6��6h4[6p�{4*�G5��6�k����εU�4>6�6�����+%6-ၶ��d���\6O���^i۶\���˂66�}C�>`��� /v6:LM��M���6��6�� ��S6�El6 �+2F\�5U[6�F6��!�>����6Wǌ5�0�6��0�0L�4���&d96P�,63��6��i6!W�6Z����60ӆ6<�6V���]`6�|S66m�6�S���a5� �6����@r3���x�,5��4V����}7�O��>P���684���6�ɀ�rl�6��(6_�!����6]��5D L6�\&�l3�5����G66���4���`�I4�"ٶ��4�5X�4ȃu5�[6�2�6J�4���5��;6\e���Љ5I7���zεm��'�86���5Mo6\�e68����+6PL�6���;�5g�6$�8� ��5�J;�ώ�B�<�>{�5�M06"�ڵ��6��:��ׂ6�7��!���~����4p�C����ʵ6h�5Y}��<4�6��`ڶ!����5��6<|>��O���굎��6��5/l6�j/5����8��Z@�6�sk��_6X͎4��)��"6�iq6�[&��d��f��6)i�5�m'6�D]5jH��65�y����"6Z �6<�ӵ��6��5A�6>6�W�5� G6?⁶�(n6�}�Rh޵��*�_V� T���6\/���Z6	,6V�A6J��6N��k �t��5�F�5�@��,w�涇�x݄�iވ6���Pq���/4��T�䴄��� �k��յ�Y�6�_�B��j#�5|�5.�o2����{6�I�3�꿵�5\'3����5['���w���5 o�ha�5%��5��r����4�k�5b)/� $5�5Ӕ�4c�4�9㵚����266;�!5 ͛�ؙ"6�\6�8ǅ51� ���"6�te6��6����}ܴG�6 ��3�@����6y�"�6H��4�^����5]t�3w5��5�� ��9������x6���5�Q�6�Iu6�	�5#�`6;�=�Z���76��l4I��2���ժ$6�ֳA.���	5��)6\޳5P;k4x���N�6�<��H��4�6�o�5*����mG���9�J\+6���5�ɋ��Z^�p �ⵆ�(�4	 �5cǜ�p~�����5M�#��;���J5�������Y�6<���셆4��60�m�`Mb3`�'��^�jW����6���1���]�l��$��6��յ��w���J����5�@���v��8cöpm��K6�/��C���q�t�)�>5	�|� 6xf61�?��,6,9g5~�6ϟ46ׂ6�O�L�ش���:��5�fӵk�d��5IY5Rw��B����8I6$�t52-S��Ә�\�G�+�5:�j��;&��=.6��C�@��i�X��26|I�4��&5�ŉ6��P�Դ��!6*˻�`��#<��ᒵ�5�6f�����O�o6[�36&�8��v(���5xkx�2�!�"y�xy[��̡4���� �5��F0A6z��0�)�71	��W36P����5����Q���5��֣���b6^��=y�5 �:����8(���0��x2�!��5JLE5�a6$�+���5����?b�xg���5+��h^!4�k��Jpc�k�6Ӂ(6�D�5ʀZ��J��5����f�6�ӵp+'���6�*��3���5��6�S>6'L'�2���Ŷ�'v�?3�����-紶�����ތ����5M��z�6�������8�	6�j���O�0�Ƕ	N]�n�͵�|D������X��-�_ds6��6,!��L�v5J�h����5m�ٵ	����͚�-��ޏ��.��L�5(�36�16hO5~�)6>���m�66� 6
����5/�b�%�6N��N�5@���,�46rG�5<���ř�5�ں���J�#�\�(6�*6����*�5 -"����6/��6�y�5�!�5�O���xL�n^75�o05�^7��n�\�ŵ��M������ ��oG6X����ɵ��� �C3�ԵH̝5�Q3���!6{q-�T�6���6�E65���\��N�86���ђ��T�6Y�9�\�:�0o�6�3`j����G5X��4����1[��'1�𵕳NH)60�;6�X5P�µ�`�6�&�0�7�V�B5ZE!��J�3������2�(��y�"��㵌+S� 8;5�tH6����#�L�؍R��J.��@P�QP��p�A4����Md6w/}50��/Z�5���3��5$���I���/t6��4B[6F�O5��!����$�5�(��[����5T�u6_�m6��*6�!�6�:%5�|���h�5
nP7S'V5k�6I�76��F<w��.�/B�s˩6xa׶�,5��5�ϡ5�5Z��6i��6�O@6@��3f�6v�e74��4���5pُ6����D����ҵ��5�餶Hw��LZ��q�2D_6Y!�!�����y6�{�����5)��T�7�ٽ5�/жm��5z�5��6�r�3��6}SW���w��4h�4~D��&�5�o��u��&+���W/�㍋��x�5P�i��!��v��5���5�=t5�666���U�6b���
64��F�,ɿ5��4�v��]�(��	6�!�6��"�Z�O�C{��̙t��V
5;Ǿ��.C��,\6޺=���O���\5 ��.��5 D'6X�H��k�5:�6��̵Pp5��1���6��5�5��C68D�d��6�<C4��ε�K67�3�>D��7�=�Adk6*D�����6x��4���~l�6�j��.�6�;�zs5�Tp=6�5�5�Od����4d}��d*6E�k6`N��7�5*ㇶLu�4�<5����s�4t�5 VN5r��l��4L��5�j��/=62v�4p�6D��6%Zb�V�X6�Mi���\6�6��N�������b6'
[� �״(N�5�.M�@	4��68�j���`4���6��2�Q�|6d���7��3XX���/���h�4�06�
���´��h5�c�P�ʴ8`��ƸU6��74\R85o�696�)�v~�6��7�|˫�� ����64��5��F�1ӵ`$e�8$[��˙��)�401�v���*`��u��b�6D�f6�3��f�6/�86�w�J�v��������4y^6�?���:6Q�]�� �*6�,�40�K5���5��3��ɵh˴C.�T��Y��5�x�������۱5kʊ6��l6��q6�k6����P��}�5N�ɵ���5{�5�_�*��6_���=6�d�6�K�tK6s�58 5aų�O�t��_�5�e����H��&6 ��29��� �;�)��	�����4�"��J����'>6�ٓ5ڰ�64H��Ե�Uj���ߵ�(�5݌l�_s���+6K�b6{��5h{��-���(<�*����6~�X'p5�e��h��5� �� .6<�5�]�j86lK�5"�%�9�Y�b������@�ȲV�Ͷ�|�63�X��k�5��`�aا5��8���6�Gi4X,�4��@�ىH�h'�M�#6��5_sH6�7&6Q����F���g�(�U��D�5H�4��Y�X�6��$�c��l�4�4�C4"Z����4�����J�j�Ƕ�4W6����>����BZ4ԏ��s-6$�ȵ6௶p��5"����\�1��5�=�5���0u�#�6r��6��6�s6��~�j�e6vQ���i96�D�5��&��,V5dwQ6"G��B6�(絹�s5Gï5��6g�X�7���a6Zχ6�ۈ5
���Ӎ�g^U��Lc6Nb��-����6Q_�
|y�@B���6H4�uZ�6db�5������5)�4ge1���5�R}���ɵ\� 72q��6�EW�~�6J� 6��6 �Dm&���[6~h���n�f>��1�$6����a�*���4�#�6����+���E<-5v#z6<�"6 r1���5��Z����2_��6���5d���K+�`�W6��ɵ���4�V�6�c5���W����06x0���=6U_�4dm�5ad�5��7�;͉��;j6��5$�6�4�(��2}��fȶ�6���4"%5���5~�'��	�W�����N���6��g�h�H���˵`|�~�36@��3��M��6�u�Y~����5TE����4 1F4X��q� 6b��26G]z6�D�5��4Ա�5�0���6n���2:U5�(�5�ހ����6ܟ6��#�T)���ǳ��04у���6��4`}0��5���6�����I6m�6��26vA��r�o������� A(��#�5V2!�<�˶����9��d��$��4�K?�����q�k6Y *�Ḏ6���5`/�Oo�5R��h�5W6 ��o�6��B6���6`� ��Q�������%�7���5��f6��"6̏R5��4������5x��f��6xQJ4������]4ԁ�5�V�+Wȵp�3���7�.�$�ʵ{�� '=�#�H6m��6p�k5ln6)�6�6,�6�,7 ��̗�6	�$A�6�Ɩ��K�����6|^�5B��6��!�N���8j�6)����.p6 9�3�%6ބ6/�����6	 m6�풳x?C�,Rܵ�5�؃���k�-5��J�7ȼص�ѵ�Q��0w��P}�4>�{6دص��u��{��b/��챥6"���B�6�3����4�L6o��5�E6�J6�&�6x�$�v����5���l5t�_5ԩ5,�5Hk�6�}�5`���ڔ�5��5˨�5�|�t��(�Pg��D�S���k5�M 6.��6�X�F�*�0]�5s�5_絞�˶�.d6^����Ӵ��6&6��5	M#����K��|J�5wW�6W�4��86��F4�^���5,x��Ԗд�Q�R�x6!���b�������8%��J�6jV�� �T�xؙ5�|�6�L�8�B6|��6�]6hk-���>���7�ӵ�Q�6������6��5l4�b�Ե��;6��5\v6��~6�OS��5<�(�;���y�X�6R?��<����q6� 굎���!/65���� 6����톶d�v�d��5$#Y5)Rc6`k�3*�4�T���zK�5�'$5n�6L��5,����b��5e�6���5,JA�pu8�h��4��մ$�5���$��6!�15�k�6���3��5]���1��)�6�X5(PG�����Dµ�9�5����⣦6���6��R3Jz�6��,3���6|=6�5��<5�f4���*6��6�f4v�$���6l�R6Ps�����6�0��෤2���&/6'��a��c˵�'n�|�)6k�5(A5�Ņ6�2F��DB��۵5�`�3P��5�56�+~�Ȳ\���s��]��Γ�4~h66�ٿ5^/� 03�(�6&0�6�
յO��6��%��Y/6�������5�4?��O;5���2px6Ӭ�81��=Y�l��5���6�x��4쑵\�;��D�4�વ��26į6,�5�#�-L���3�x0�5���5��23A��5���5�)t��P���͵Ơ�����6L�l� PB4����S���-�5F�5��M�ﶄ6�Q6@�4��*6����ô��5t4�1�L}�0�6FO��[$3�f�5_V}�|cV66o޶>��5�9�5<����=�)H6������6�R����\6���4H�)���5L�����7���f6��n6ώ�6}����`y�fP6_)'6�����v��96O�5$����V�4[�x��y�0�I5P!�5@с��40��Zw�ęd�䎅�&!3���=6C�n5������ ��(6�����N��5�f	�6���ܷ96�-�5m36"J�=�2����4�x�5��¶4�Ե٪5^�J��5�5�4��M5V���!���z��6"&ҵ<G26h��|���,5�Xt���ӵ ���������.6x�6�D)�C�n谶W׳�:"����5d[p5���tkt59�6�u�6��3�JEƶ0��6k����t�4�\x5\�T�HY�5p�4ڷ�5ĿI�uѶ!6U�͵2�6j���t�����5�>6��5�Ȍ5R�6�'m��E�
��2�E6x�K5�xu6�aU5l�6,㗵|����Z-6���5�^�����q��mĻ���4n�~���6����o��v�x=�N8K���Һ"5��6k��5F�;6+9ö�T�e��D����x�J1.6ҙ���*5��36�5��	�A6jd3�L�6譑�1!r5����-Q�5&'�6v	 ���5������5��6�e6x(���)6��5��ٵ���5[#i��b��"�5Э!53 �������5����(�16����kݬ5�(6��n�����Ҷ*�-6_>6��W�ư7���!����H�52ښ�Dw:��%����B6W��-.�@85O�5j݂5�Y���%5̷�$�"5_T��|�d�F�6�44��X)Ǵ!ܒ�
mq5j�H6�&��Q��0^5�����_&����5�A��ߌ6ڴ�6��Ķѯ"����D��j��>�6�G���p5�hj5�5�Ff6m~r5��4��Z��;���5����̒��a��
6�G)6��96�٠5)L�V�6r��6V:�ڊ����;5��4ҁ�5��ϵGT��$
h7�'~��>3���7LjȵOj\6�R%�� ��F0a�b���bX7z ��z�����6���$�6~^��d�?H6uVA�y\�6 ص�8網's5�:�5�7'3G��DW7��6����d� 7QE�6�t,7^���x��5����O�6� >6����R6��6���07@��4NZ7d�K�V�W7�����*͵�7��**�6��X,�2��6hV�7�F�5�#+�o��6I� 6@�[���4��[��.7� �7`̻��5Rm���q6D*�6>�C7�{Ƕ�R���3�~'���n4�A�.9��Ux��0�4��6�ǉ��'r��ΰ6|J6����ꨵ�e����6m�a����Uz7�ɪ5����R�m����5.��޶_�����163�6I��`V�6��7s?��Uq��2Y��e6��O���ĵ�ݻ5�$7�?7z��A:�6.eA6pr�P��3 �U1a�� �\��f�5r6���64U�69(6��c�3��Z�6x���,�6����ռ��ǋ6�/�60|�5 �����:�v�5����""��dմ*�[5Ly6&��6'e�6�;�6P*6=�Ǿ�~��h4�6���6)��6�<�66Q���l�����L36�ֶ��6��5K��Z��6^'õ��=�C��7 ��5���6��Cǩ��u7&F6P�x�H��7#y,7��n���.��=1��s6�j��-�=��\<�6�;�6�0Զ�=�Ґ�N�7(�'���qG6%X����4b϶6 F6���4��7X7�7O��6�6��)_�C#�6���6^�Y���N6�?�6^�b��0�t��6�U6_�6�啶����=5�	67'`�mZ6��6`a��-"�6�[X�(_@��J7�qS6�7V�5�Y�4.�����qb7d�5K�6l�6�59�W��BF6K$Z7��6v���X��d�5����z�\!6*��6Ǽ%6����Ң6��z5�l�� G>���ǵ;!5�NT�;�6�tŵ�u��}�6���8e���6���@�84�A��ݜ�8v52��K��5�M�5M��6�Tŵ��5�����/�q�6̞7Xy�6� 5�����h���}��S�5_��<�6:��5v>��|��5$C,5�$6���59W6b��/���m6�H���b6S�N5�z�xYK5�|�6iF�6�w���q6t��5�W4�ϵ&ğ5Ê&�w*y6K%76��5�vT��е��6q+�6�=p�7���8��>�56�,��m�����5P�T4���Χ�5V۞6̒����4�
�w�5���H��4s0ӵ�w�6Y��˯�6%�6��5��(�ۜ�5Mݐ��h!��_�����K��5����t߇6�6�F�6U��:��l��4P�6�õ�r:����5�.=6h2R��>U6�l��|Z���y5�W6�ˣ5���������|� ��2�cy��[��Gh64���xv�>�����6N
]5����ܵ6}S��6a6)�ɶ��R��.%6�1�61��|�5���4qw�6���5ݨ_6�tV6�]�5�=�5�f�ws��8�f6u<6��j�f���w7:�� ִ��|/6vM6�t�j-6�2����b�5ph�5�_�4��f7'�=����?7���?�;�4 ƹ3zl�5^� �e��6B-5d���V�6�K۵e����7�y{� t4�h�Hu��o+�6�����6�d35�&�6�c6�P�O��o�58�O6j �5ח���86+�Z��9{6Q�$6I�6
����b3��H����6u�6�����4�Y6�x����6��15�V�SC�67)"6V��$�!6j"��t|�5�)�d�ߵ~��51���4��.��Tf�~6�^X�h��6�jT�,�?�l/õl�����7��h6��B�#7��r�`�F6���5�g32=
5z������B�l6*6�g5~隶�C�6�	���0p5*���ո��T�5x h��o�V����Q|�V0.7JhC���5S#�\����z6tk���]����6F�ɵQ�����+7��Q6�n6���5 /�5�65'=˶�Iߴ��+6xRB6�36�-5�ߤ5"�S6���4�xE�&g76�����r�5��̵-�w���%N660�6���5u��o%5��3��ƌ6�/�
}6:�
���34�����B�6�ض�����6bD�5�O��m�Y5 (1,gS5s��6���ޡ���}6���6�;���5����,56N����6g>6�5{4Te�5�u&�|k����6܌.5�
�AbB6dˁ6��h68�?5f�|6���p����
$�0�
��_�6�狶�x��ђ��M최^g���D���`�쉅3��ʶ�P�=�6E
�6�B�^T���Y����5ӕ���߶��6�o�6����K��"˽6���џ����O5N�5aC�5z�v��ޯ5�֕6Hv ����5\�6�0�5VD��2�V��5�4686����D��$��5��[���4�6ly��{�6���n.�h��7���3��ў5͗�5����e��d��ȵl�$��f6[�6�w8��Ė4�-ѶC5�'ߵ�P�4_6X���u��51�6��崮AD�8�84�fֵ4����5����������L���� ,�P5&6�3���=�6��6~M�5&A�5 ��5��6�^�h�41B�6�ﷵ}�6 Hr�, �4 ��4��i5K\¶۽�6��M�V��6��!�����5��ô�o���L�{��H5��'6h��0�&�6����.6KyӶ'[h6� :��ј�y�^;C�U�����5m
����6���6GMq�ЦW�6��_��Q����5 ����[6w���%p5N����qD��L��26`�^5�e��|B������BŔ�5�����Hr����y�ڄ�5�����-6~���\6J�6<4���+�t���@�	�����-6}-6��/��D�� }6�<l���o��9�SM��a��6}y���յ�.�6>�6�m�5���5�T�6{�ӵ�0�΂��jUp�I�5��$5p�=�wC5�>ӵj&k��n���_�5�{5^ʓ���=6�?�5Oq���5��6��6���5�� �@�a�)� �@��3J0�5&l 6`�5��4�~:5�ߵ�c�6|;5�hE�����h��������6����.��4Ʃ�63�n��^_��S>6�W����5n���?�A��*�3�L�4R�5ܳ
6ؠ���b���%5�GֵuX�5@�3�Cm� #����D��i:��X�R�q6�5f�����驇��͵�B%6!$��"T�P�ӵ�J(67����"u��|�5�U��ʡ5+w�6Zw���+6L ���6�s��LM�5�Q^�K������5�x��������6>~6�۵���5�V�6��l�h�X�����t����Ƶ�N(6,�x�$�]�P�����5��5�?ĵb�d6c�)�*&�����5 �K3R��6�ǵ$�A��6a��5Tv5�$�64`6(Z�5����W�5��5����ԁ6Z�����&���5����!�2��P]� �n4�s{6��b5\/�505=�7��B�Ȳ(�PsH���Ե�JI6������5�� �V{6\�5��6��P�`%��̳��j�7C��6EH�J6�p�6�d���:6�6�'�D��5.y�5N��8��5�E����Z61���泶8��5��41L6��w�(%�6﮶(?�4���6�b��r̶�'6 ���=�.c�6Eϔ�zO68Ӝ5<2+�2DZ��P6��e��/J�쿞���=�M�96 +�3̒5k�E�Bb�5���5a�6�g�5������7�WB��Yk��&�6�[5� ҵ��p6TVy5�+��66��5ێ ��7���]���n�4
��5J���|���S���B���|^6��X��4K6v6�K��v���S�6����y2]6jh�����6W����_�5�:�D�F6vd+5��̉�5���5�r65���gF5�A�5K��5h
6>]06`�(���,��w��Ҭ�6����6��D3�s�$i4����r��5�k6�Sε惥6f׌��g��V�浼=������66 g�4�"66�W�\�ζ5k6l��6�N/���A6Ƣ�ЇW6���63�.5�N�6����lU쵄T66@�0�:���tt�5@e�3��)��2q�vh6�k�5�~õ��36Z�^6�X��P6��Ek5)m�J[�4D%�E\�t��4�36�Ķ�26J���NF��1���6&����	 �ײö��6�Y627n�`-d�&���s9�5��+6"7��u:�L5��k6�Qe4S*�A�ֶ��Ҵ�=�H���*6:�5J��5��� �A�^Ź5N;6V��6����U��os�58F���2�Ԁ86Pd����5J��5I�R56��9����/A6�9�@��3VED��x�'�:�$��������x6 �N4�Ҵ�Q����5��6A�5��q��9`��Lz��)Xr6FC�5�Gj��kU�&s*5R��5�ș����5E�(��'+���:��RK6"��6�`e�䃝�@܏6e7��aY�3F�6��8:5u�76�Ɔ6�.�5�5~��6d05 �4��p�4>}���"6C� \5�[n5���5�����^��ϟ�i76j6,���T("4��,��C6�:���8�\@R��\7����#ZN��'T�jT�6M-�z��5�l{�Э�5�:W������6�6�貶�t5>e��ش �g�X6m5�'ش��)6֥�5�Ձ4�������5����˨��:8�n4��)z5-&F��qX5�Q�5��ֵ��6fB�4����J�5z0������$[���9�:�����n5`Pj5��95L{�6�s����6؇�5�;ɶJ��5������w� Kv���6_�g6^��52r/�h�6��ڶ
���P�4�I�� 7҆/��
Ƕ-�6�Ճ6�i�6����7���4p7�ɦ��8恶L��6<��4
�6]U 7��{�F4��-�5�Q�6��]�"�b����6��y6,}��>�M5�5���6��R5W"��̬ڶ��4��a6������iFy5���5 �j5�4y�6����ȼ��5��d05�iz����5�r�6��05��f5�:�6Nw��${���5!a���%U6Pܶ5��������H�6�#6,�״͵��^o868@T3�OV�����D��'k68 6(�>5����������0C��胶�fN6 �4F�{���b�rls6`?������U�4��/����6��� �}�b6@!02^��5�hõ�>�E��g6�t�FG��bm�\�
��g��z�X6�5���6_+6B�|5 ���w��&�6���6^���"ڏ4��5�ǵ(R��.#6p뉶Z!��흋�
��5@_�6��O��6��Ƞ������u�cZw6����T�G�z@7 'Ѳ�A6����6��P06)��ؓ#6�%�5�ɘ�Hf5`ae3Z����(̵�m�޹��6��x��pO�G����86D�����G6t�ڶ�i�6V�����x���I6OS�5~�Q7�)�5�~�5�δ�)5�1"�p��6]"�L{=���X6���6^B%�B9�,2E6���5�ִ޶�������/�6�E6؛G� ��'H6�r�C������R��\��OLö�~5�>��5����p�q5 ���&Q�l�@�Pള��T����v^E6��-��F�� � 4���G5��)�l�L{���z35O޵[��6��06��>���5x^5L��5�AB�oO�AJ5����a�6���5<��0�60�2�����5�������筶Ё��l!���#.4��~5�ʮ5�K��m��^/�_6�M�5Bs6�j��jx��W�P/�3��4�m6vN�6���6o�����c�6��ɴߏ��۵���5����
�����.6ET6�%�!	6���*�6�7�6�Ѿ�&6V��5������)o�5p,ڶ���2��6�W�6���}+6��,�q"������<���f7h@X54�5�hQ�Jv���>�6!�5�*�@����	����5���ɦ��2�����@��5X0���K���6�5SN��5.d�����@\U��}�6�	�6 ����6��5C��6"��4�E��Ô6�xh��6|��z�5��w5_P
7��Z_�pt�6>_*6_f 6R����46�-�4)0Ƕ4@�5���5�&5� G/��_�6��6��V5 ���6�(77�y�6hm�6�)�6�zi��|.6 ͵.�g�@���7R`6eQ}6��r7��'�Ǌӵ���6 ��3n��4�06�1�5TֵH���58��5l�=�K�����6J<6E���X�ϵ/��6�J�6��w���׵\�"�@�̵�č5Q�n�W��6,��tV���$�w��m! ��a��n6t��`^[�\��u�P� 4~��6J
�5�6�\�4{�5=cx6�� y��G
7�Y6�aw6�nP�������6��s6�l�Ŷ��w6�eC��㐶f�V5&m~57���[F3`ߒ4�E$6@���5�Y��`aW��+4��˴����@���ǟ.��8�6���lQ��
��tX6pUR6�ĶQ���Y�5�����!6�#6l��5�ޏ��*6��z6
6:-z5#�5yƴ#+�6�+�6�h��p[6)e#5�o�5χ5�|�6��� �{4�D!7
 �5�Ѡ6��%6*׃��ݳ5���5Xr�5\6�@�5Vey6F�5�|A���4~�%6n�54f�i搶��ӵ�w%���6���5{��5ܒ�6к5Lw�4�C6�ֶ�p;3�[,5���4u��5��u��� �615|癶/#6B�Ǵ0~��+ķ�»m��â��O�6Ļ�*�6"-������5��b4�'i�Tp�@������6���t_�� ���H�5~l6jY�5�kh��|����m�B�U�0��=�5	���  �4��۶������5"A�äd�8X���9r6�7}�Ҧ�X$���?+5"�ߵ9"������F6��o���v6����0}յ �d��I�6�.�֫U�N]���\6t�
5�5�Ľ�ў;6�_	5C޵(ǂ��P�	�5rٵ4�6�'������Ӷ��t�"O86���d�6 �5n+-6��B5�U�5SQ6,����6fĸ�XӴ�F}5���6�����r6y,�a&6�`7��϶@���hd6�}�5 �p4��G�²-�%6�^l������5C�[�Ӈ5\�6�D�6ZĢ��2k5�x�5{Q��$�X��bz$��(�67�ݵI;��̇�5���Z�����ħ/5��-6���T�|�<u�۳�&�A�.M6��w�L��5 w;��X��/�#�;M��������.�6�R�3�H���L�6⇭5$#t�8n�4x�X��v�5,m�6�Ӌ�g�t����5�46<�����<��3���.�3��7>X6Oã5zC�� ��6&m��̌6�{�6
F���6����Z_�� 66:�6X��L��r���K�O6wT�1��6kد�#���%94�A�6 x��p�60]&��S�5O�
�s�㶆�C6�Z�5f�6�յ�������S�B��6� ����6N6ta�2�@�������8�jL5��4�x	R��AD���\��jmµ�<���9� $4*�����5���6��5n�6No� {��J϶o_�-%���ζ#ɉ6��$5 �۳��4� t5��5T�5 �(5A�������i׵ ��3}�ڶؔ6Ud5�A��Te�6��S6{e۵�>R6�a���Hc���6��õ�͎5�F��=�5Ǌ60Z4��5�6��6�u�61]��_��F7q6�M�6ǽ��д�c��3;5&�>5�۴�bZb5���5���5��&�\ʵ^��5�����5�=�DCմ橛4��5�����K�W�1�#�6|�K6�s�5l��C06r��5�z5�5��5�+6�Y\����5��6М2�P�k6�	
6��4(?l��@�5����`��2/�A6��52� �}6��S�c��4X(��U4��
��7OG6�	��{k5����t�4�S35��ôܕO��o74pm�3��I���Q���4������*6�&��ꬶ�p+6�[.�p�;������H�7�674�5B�-61�˶��5�9�5v�����&6zpN5�I�<^5uͩ5k �6`ZY4��\6H�65^xR6�ώ4^��5I�W6�#��	54�76�-��x�9�D?�6Q�����p�72t5��t�E6s�ж�5"��5Y��c�6�d����q5�[��չ
6���5�<5(El5ٶ�u�ꢅ6G��5��Ͷ<�c��R6��7��� �5�P�5�05�06ؙ�6�=7�A=��\��3�6��>��G��m����.���ǵ��6X��(9�6Hl 6��Kg�6\�6�͒���[6��A����(G��z�ړ5��6X��������r6�À6@�3�fR8�ZA�5XI*6p���,���~�|�׵Q\̵��"������p�5�:�6��5�P�6"Z6��)6�4�#��Jz���e4��~6�@ӵ��C6��M�����1��r��p�3��j��F����"_���L5n4�5좵��c���6=>��Ȅ�0�H��F��8���5�6���J������66V?6͏�8��޵0U'5'rѶ��"�͝���)h��t�6\'�5��ڱ���`��f�����7J����΅4�����]6�~�gBN5�S6�n��ua���ʴ3��Ț�̡жL�5Aٜ�^�6<x�J˵�0�5��15��7���6�NE�^J	�J�����4f[�����w6���5��6���F�쵞�+5���6�3y�+�0ۥ�L<��ף6x�15j��
�&K�5,G"6��44С6Z7�5��.�6.�6z�zF5���6����[5�n����W�$7��)��7����zA6���6�*��ҦI6��5l������ޫ6�56��h'H�/~�6U 7�Ú6 �g���g�P�5�I ��r6�:+��
��n���g��6�L۴�� 6I�5�g5�N5���4�<ܵ�U��`�2l�5$�+6 .´�F��6��(��T�5���5�8������,)��A���+���n,��q����6l��Ķ����n�\rl7�2K��ǵں��:�ʶ�"?�(ˤ�o�5�V5�眶T ִ����O� �n�����#��|�h7q��Dϳ��6$��6��6��8�w5�	�5j�����?7�5��[�:��6~!6�2B5`U�5ޞ�6��w5]�5���ݝ5��ж��G6��󶤉�5V�$��!��Fۊ�"{�`V�2  �0��b��b	6@˫3 ��6H��59i64�趌'X5<	¶�3��`6�� Z��Ԙh6Y�E6��\��_5��6&t�����L�z޲�8�3{��j���J�6��6,�B6�eߴ�������6Tۑ6�\�_�T6�6+�6�GD�r�#5�w��zc�5���.1i5m�7����������6е4�/��56���4e��5���"�Y�a$A6�۶�3f6[e���5�-]���6�����y��Z���o��c�2��pHR�p;��sq^�(iϵf.K5��z4u6>t��/ ���5��2��t��2(��xW6��6V�;�h�5@�6���``��I����7�O�6 ���	T6��n�q�_����6��W�5�x�N����N�6@I5ac��V�5aƵs��5���vҋ��H������L��5:�ҵN�-5&�e��}
��'�5b
"��`)�1��5����8h���6��[�C�xߝ��^�4�b5X#��Q��Q ���ĴnV5�3m5�C�59=�5��<�z1ҵ�T�5bt���5p��3���56N6�۶�5RA�c��̆K6�e(6l���N�5[a�_]����/�S63EH�h�S5�Q,���5	� ��	�{%�6�s��u(�6 �3�6��6@
��p�ų�׵��5�Y��Jp�����G���z66�c�J/6(�;5��T�����*����3
5I� �4���59�)���T�56Dm6�Nl��6Q<׵�\5���5T��[�4`�6h��5C^?6�kͳ���)�5 H5P��6|/c��Ү��V
5�]쵁�����(�\&W5�/6"%��ǂ<6 t<�e!	6`��l۵�Jҵ�⢴���� *6 3N�$��l��Q6�ǁ5lV˴�/�4cB��<I�� ���d�5;��]!�c���L��	�6[���/�,蓵���j�5,S���O�4�zD6Vp�5M'm���5����X�5ت�5�Gy���59�۵x�a5�<V��P�J�$6��;4! 6)��5\W<6���m��6 ��1=�B5��47�������/��;쵖��5̱��pxB61n5�F3d)�5S�62��5���4�5N6��^�.5!�H5�UJ4|�[5�VR6������5c�6Vs��Z�l5����d����n���%�, %6���3�~�6�b�5���4�9N�j8�5
76���y<�5���5ʞ�5�O����,4lwX���ӵi7Z6�K�6M��5�LV4V!���b���R�5=�51�/��V�6�=6���5%��6I/���G�4#�=�d��8�е"V}6^����{�S)��{Ĵ��4�M�S�5��h��`���'��*^.5��$5�36�.8�u(�6 A 5�����6��6�v��Wj<�X{�K�ֵ�H76���62�i6�5��{>b5�'4�)�5��"6]�6[[�6W��6�౵���%�6/*]6(�J�`q�^:m6�E6�k���f�)u6e���0�.3u/B�p�,6ۣ�5(���E4Nɒ�}��̘06$0�4��J��5�ͥ5T7��x�54_)��$66�=W6�=`�q� ���z625D�Tܴ����h�ޖ?6h�]����v����*5���4�vM�|U���<�yְ�z>�5�)ڵ{cu5#�"6t�ɶ��5>?��
'���'�=-�5T�5����6�F�����~�ҵvG�,�6���5{���ڎ"6>>�62��5�Q���l��X�5���5豳���P3��'6���ń������v�5�74`���cK6� >6�B�6��%���5�Gk6��>4�j6�D�5�j6>���d,	�(�74��>5z��5Z��5ݳO5hG�6R�5`V�� d��ܧ�o!��ݔ�}j�6��!�V��6�d������t�4����Ga�ίW4�s��a86��b����6�O�!4�5|��'N362Ej�V��gS��譏4����5��4V;�5�Ƹ�� {5�ݵ�ى��}=5� ��`�`S� �55��6�� >��	1#�̻P6�r��4K����5���5��5�&�&�6�86`�ӵ�!l��K�6p|�6{�����5�hȶJa�66<�4Ѽ�5�?6�����5���� 6p��6�eֵ�Ō6��+6�M@�p6P�"�lTöAN���]f6���6%?��h_4� ^65��6E�16��f�"�5F���&�;6w��c�5�B�5���5�ܖ�236��~�T�z6p�6vX�|���@:h5�q�"�E6਌�E�e�~��58�6Yn��2ߠ4B���Lzx4�'�=6� �T#6׶�5����R���06<6`�69����ߵ��õju���*6s�5$���Ը6ڷu��ϲ6L���r���$N64kl6�B�5�o��0�O�0���m.6�.-���06h�!�D4�5���5ԍ>�/5�5�$63�h6�=5���+d~���60����u5�U޵�B5Ǟf6�rr��d��~��� Q59뵄�"�i���i����AS6� �5>�667�5�ޯ5T
76�S�6������4q�6�w��Jg�#��5H"��2i6ԫ	��;@�t�7��E��]V6�)��  �/ �V��l���˝��?W���~5=�5�{�5L+*�l�C������Q�\t5�*M5��v���"5d?�6�M��X/6�J6ρ�5 ?��{���t�ܵ�U>�P�5�tr5c��6��5��X67E�4�'6
�6p&e�Q��5�ߟ��:
�� ^�N���5~䵄۵�`����6�5X6���5�ӕ����56�"�:i�����PVε�ԥ4�4�5��5�\���L/��W�5x`�Q9��%4��
��ś�t�F6�8��q6�}�5F�5na�5f+|���(��65xZ�5&�����b6�75���53I6��5E6���p�� 0>4(�:5����p��4 7гoM 6L`r�\v�5V�5�Ƶ���5��ɵ��y5����j����$5p����+���ɵp�ôu}�5 �ٲ���5.5@z�,J���5ܱ�����c@,6J��v�,6���5�2���UԳ@�3��!�ǽ
6B�(5�n��� 6�Ǚ���%���c����4��4�X���Y5��i6^�C6,˵�(5����toQ6��93��2���v@� ����#5P�S�֚6�ີ
8d5�L�5@�$�|�쵈e��f���K�{pW67���pIv4� 0��m�vEϴ�F6�kt�@��Y�5 �����4Gݵ5���5�xH4"�5� ���3��4����`[6�I���a5��Q5t�5 ���,<5�����^�5��`ų,���nA��z�?ֵH��J%�5 �(4H�[5>�D5V�����5��6Ys�.����7��H��B!�6�����2?�8��6�笵@m´�#̶�k60�6zkE6xtZ��8���h��+��GY�,Y6�J/5��a6~'7B5��+����W�5���6+����x��H�E~��0��5�~���Zg6 @�1����A����>4+)���,�605�pJ6�͋����6:K�X�6ؓ�6d@,3��׵�����6���3U$66�ٵ�x�6`M���,�HD�6e�L6ν��q>Q6��ӵH��
�öI\6�b޵�={���5L�õ�C	6&浰���f��>�5��q��6�Th�R�5X�j���#��L26�ޝ��e������ =6��S6���6�B�����n�V���5ea��p}D4��Y6KH6�<a6Ѐ�4��"6G�6��v6�ŵ M�6�jD67a�5��d6�)�^n5�5�|u6NԵ�뗶\��z��6�06�R�S�Z�f�9�� �6:��#6̤9�`�i4�q��a��5N.���25�P65���4�J��5�M�6	kŶ0Y���A��� ��m��{F����}�-��5�˙5�*6"�5x$G�Jk�5�A�#6~�+_R6*A35^���/�sŢ�0Ц40��4�yK6��6�Eh������f6{�/6�'6DG����5P`5֭6�85,|��GrA��`k�>�㵛K������!�5��6 �W�`x(4T��5⍳�0m�5�ݺ�v���j���ip��s����t6T�N68W7�K6��6^d���S�5xS��\@l6ȿ+7�G��S{6�]�6�\��r������BA�6f]̶ٶ6����8C����68�d5�|w6��5�聶�����
��U��IU����4@!4�;!7 uv4���5<��5��
7�_$��u������Ncl��v�5��Ѷ�$6
ե6�,4�?��ɶ|j}5��-��^7�9y�I&9���+6��a���I���6�S6�V>�������w~����`�!�Q�a��8�4D6���=����56�^�6VA6s������[�7�{?5��n�BcA6a<6�e�Ӏ�6��m6�A6=�X��6�ä6N�5g1ɶ���5�~�)�G6usݶ�%��t�6??�V�7������U6 H�5.S�6��	6w��6~�g�G.�6��I5�&g��H���N���k7� �����5^m�6���6��*6m�x6o�6X7�B� v�~?�5ğ�6�\�p˴����"d�6@;�o�Ͷ1K86P6 �Y���󊇶h[��Y�S6�<6@6�#67l�5m�t�T	-��
�b؀���z6��� j�4��3��1��	����6�L��h���Sɶ�L*��X86_M������F��6H�6��55[x6����v��5�>q5:�R6�h�d�\��϶@Se� %^50��5^�5��ԶHƍ5�z�2j6 6�86`/6܅<���"{�5�')6T��5vR
�w![��"�	T��#G����5d�)5�O4��t��y�W5.����5`J���J6�3���D	6�z6Z6G���S��6)���K^6��5{N6��}6�{A5�ʪ6x���	O� �;pP6�
$6��@M 6�����S�4>u�p3l5Dlq5�%���T5)�l6 �+5��ܶag�6�qs�;سu66�5Tw�5��6�j)6H�)6��]6�6�������Ǵ�v��aѶ������F&����6 ��)�6]7=q#��i5 �,7��}6�!��9�tWW��ږ68I6��6\5��`�6��۳'��e��V6�0p�o��*3 6xsζrS�6�
2�Ȅ�6 	����4���X�6�2�6x�v��-5����<ڶ�Ҟ6v�e�C��PYٵ��7�X��6Z� �R*�5��6,���6Ə��0��\v|5e���+����ɣ6���58s4�쉶>Ӷt�O���^5���66~6��Ǵ��6\W��¨6Z~B6u�K	26�S���1�6�<u5&�/�����;��s�5l�6hn���ĵ��7�K��ܥ��L_�V5J�`SU6£��i�1��P[�6
I�5�0�H��5���B6_uM60^�4Ҙ6t�76��?62�}4�2(5��p5����$�z�5Ny}5#��6Te�?ȴ���5��6����
��6�o/��Ba���ߣ��H?{4\D�5rnE6�=15���5+�16�{��#���N6��ܵ��K�vx�52(��������CD��]���20��:X��j��6���4x�b5pD�f�%��_�4��5Xx6u�b6& <5h�նX;q5@~�3L�6e<��s��K�6 "� ���;_6�٢�,���י�6H�4gz(68<�^�26��4�8�ش�nG63 �Hg��(*�6�+}��6"�%��b��6*�,��w��UBB�l@��;c4b���i�#6��@�2���>}6�T��`������R�:�?�r*����6?��3��$Ys5GJ�h:7��J�B���Ɏ�%�z�f-���+Pk��_��j�5��	5�5*hܵ���5m鵢vT��5�7��Q��H �5�Ğ�L>6_����I5�t6� I6�/75qV�6���5�7�52�5�B����yC��
�p�35=�6�B�5ָ��W�6��4T����s�5���5�s�5�(�5�j7ą�cV�6%ɲ�4�4�q�ض0S�6���P6��36ԃ�5:G�6 �E�2�6�Ŕ.6����"0�~�4�1��P�5�����ា��m�>�6��ʴq����;�4HVS6Ll`5V��f�6{߇���i���}�t;*��mq6PԵ`�!5����;�O���|6�i6@h�hĵ�3�4���y˵X%�ďq����q��b�������,�H�N5��Z6�5�긵�I#� �5�d��B��q@�Ki6�A��!׵,�]������5��N�r6�i6/�{�#��6S�i�|^۴�%�N<�6Sܵ ,3��V6��!6�;J�00
30��34f��4�4 ����n�5>��5��S�j�8�θG6pk:�:�86�A@� �4x��4�\��ǅ�~L��b��o6-=��r�^�����>��H�;6h^����66�o���5n6M)�)�Z��X�0 ���V��TX|���̶k��6����T���o��7��-�2����x�5�
6�kd��L45��#��:�����5���5��{6��4�%|��:5e	��B�7�dV6,[��o��#P5z6R�,6��\6�%���m75Ώ5{�嶘�;�v®5|� 5D��ȈԶ���62e��<�6D,���6��6D�6�d6� (�4B�޳�;H%��6�玵 ���,k6\�o6�����6�6�x��W+�4S��4"�6uܭ��bϳ���6���8��n����+�5�N�5��6��6L����ƃ6|62D��=6���5c�$6��5�ô�+�uWx68C�5H5\��𹓶8�5�W��e��$��4������5R[ �J=b�,�c6�@6����p�6pO@���f�:�o5��6\4��355�5�I��Z��4��������I5��w6�"j4oʵU[�S����Ѥ��ڈ5���5#Pq5 6.ƻ���>�Fs�6��6e6�4
6_�͵x�6��j���p�I$�qP�6#���B6^��5Bif6�b5�F�6�!&�r6��|�5�3���5�M�N�h5�׵�����d��F!L����0L���]3B8�4�Q(5����f��޻�5�W6�����$7($D���6N�F�0ѵ�86��]��j�5D���(��A��5vZZ6���ꁵ��H5�!��1%7�1]6�ݵT�6���5�����d�5J_��J�&�/�b�B6�ލ4ĝ���\52I��ӹ�Z�U5�0G5��45�Y���eóL>&5zT��g�3���4y|�����6���n�̵=����n[����5����D�.�^o���5hk�� {մ�~�5NV�6�%�6y���(^P5pO	5t:v����n>��)��6��5��5u6���6��6H���H"z6[�(�4��.6��,7�x5�6^`6>�+�n��5l䨵b��5*S�݄ 6�>6���5l}��r7�:U�sf6�	6�6����p2�Ƒ����|6l�3���7n�(�&�4>�5�J�5N6T�6dM5���,x�����4�v����86��G�T#6�#6^�A65|d���k6��e���.6�(�@��4�k#���6>�6 �44�2d�Yt��$ٴ侌�3-�5P�!�P62�+6܆Z5�(�5(�5ͺ���6 ��m؍5�t5�q���ȷʵ����0�������`y�n�6�U���	5<IN���6 ߲�7
���5��N6@�5.�x����������+���,6Bz`��U��ҹQ6�m����^6���6g ��M���ns�r��6�y��7K���~b6(�i5a�6�n�6<�76���x-�6�/5k6�bo6�7=�8s����Զ�����$5=bӶ@U;4]D�����54���썶tF�6t�16�$7x�58�ƴ�l1�Y�J��dζ^�߶���X;�v�ƶ4}[6U;/���5��(6z0K6��5yvN�O���5���4]���lYε�)?�<D�5Ŀ�"��6�蔶V��6�?7%���]Z5\��v>7 � �E�������}���g�.�s���5(����*6D	�,����.�5 �㴵^7�@�6@�6����N����5�Ik���=6!©5-9m6������5��@y04��6��6��q?�5�06��˵�i}��ŵD����ѵdl�M"춬�c�(/16�u76T�h�`�4@�h�FZ6���$�j 6�S��:���*6A[5��?p���
��7@6��$L5 �ȳ�a��Z�C5l���Y�B�H6 G1O�W6h ��	6�����6��6XyF�h��6�ج6�⡶H��K0����6�/7�E�4/�>6ȷ����{����5q��6ր�5Η&6W�5� �6sx��v��� *6&��5�65�ޥ���#��������4��5f�i�5C�6�,��H���������6�8���	��0�6�&+��c�3�%�6b]ϵ0h"5��3
4sm��`�5��Ĵ.�ٵ��4��4xҼ��
��x���/6�5�n#�(a��&���_ࢶ1�76t86tK��M}��ϯ5��<6pQ
4T)Ŵ�1�R�4�,��w-63ͯ���g�F���С3��{�6�1��yL�6���	���S�d5 �L�6�:�}�6�^��\�6j����c6�I��Y�6vܴI^ƶt����f�6ړ�f����[��rr=�@x�3�"R4TNa6��̶ȑ�H��|X� �����64����50�6����;o5C��5"}�5zX$�y5
53L���(�6^����m���9�6"��اS5�
�5"��5��*5TA�4~�5�Y����66i�%5�;5Dz�5a���L%6���5�$4�����4�T�4�א�_����c�5 iT�Ls#6X�\5��� Bc5�	�2�5� 5ʑ8���4�S���R�&��5:����v6R��5h��ݽs6p�`40��_1�5@���Q�kJ�5AR���c7��Y�5li5��5f�&�j��5 ����D�<?6͗6�L7v��|��Ƀ+�`��5F\�����h��4��5���4 �̲���ಐ6��,5FMA�L�X�(�_6�߫5����oٻ5�gB���n�l,ʳ��6٘�5غ5��*4�3�5.�ĵ���0#�4�/36���������5h�56�;�Hjb5Ο����C�n�	�j�s6��5_��5���3N�4��36��.��5(ձ5�d5�T�4R@��<g!5$n�5	����$���5!�*5����*'��!״L�86�5�6�ǁ�>�5df�5�_���Q@6@S���#�rߓ�V�F5��
5��N6�A��B`�6Y��R���
�3�s]67��6�^���g\��a�6�},5�t�56��5�6�	!4B�쵞D�47��4}��;&��6^\6�&����������1��57�_�J����\t6�H6���� 5V��ܴ�5i*�EB��iP5��׶:'j���&��%�|��5@�6i���q#���ӵ���|�7��C5NW'�op+�Ȗ�6�������59�6
]�5��y�O��܅�ߚ5T�6#��6b;6�]���p�5x� �"3�5���6�~�5�ȶ6��5ָ��K�B7�����6V�5��_���2�V6�jX���5�6��(�B0-6�1����6�~i��`�6/��5K��6^�N6��J�z�)6����"�6�5
�.�66�_嶰��L�5�V?6Hh�5�,q�J/�@��g^W6�"��R�6.�.7��
7&���;6�[H6�2Zp@����5���\��4���<�R6�d�4�A"������K6J���$��6�:*�����( |����3|��6�C��c�ֵA��6���6�h���w4�h�a�СC6ֆ�5Lw�6VZ5 �$�wuP6����9���5�ܛ5�[5	;b6�p�x�u��9�6��$6|8y�-��5w6h�����15�6��5d�7����5��5���z�6/��6��"�w�z5��6�t6أ�6�����˖6� (�P}"��)6 &�����y?ƴܯе���5x�z6I��xL4��䶓�5򬵶04ȶn+�5�妶v�� T�6�5|�E6P��6�>�@��4�W�`Ir��M�5���6A>ֶa���Kp6L��5y��5�5tފ��F��}T������6����X6A�}5�+ 6�)�m�6�w�DB�f�6��!6,��(�Ķ�ץ6�8a���[�J�,6����\Q� ��Q��(�����5v�� �]��H�΁R6tv@6��4�ш�$�J6&�5�6LYI��9�6*ݵ���40mv���P��4@��4"+�62�4�m]6�<�� ���`�q��2���5�H�6"8�4�",5����c��]�5�쁶�:�6j���U5�S�o�6�U�2��5�33��C 4���M3��i6��_��6�\&�|�D5���
@D6��5(R鵘��4���L�5�3}�I��>|6
�*6Ⱦ���`M��N�$�����5�3[6�o���26�f#� �� ��4��<ɪ�5�������J�1���g'�:��5 �6������´bеL���)5&F���;�6����F��!=`�Bg��L�05؊5 �2*�������%����495�7o5 ���OH�5�<�V�~ ��\|6���6�C`���5h���J��5`c��X-贷�"5�L���,!6��06�J�D0���54���5�q���݆��o?�~|o���6�`�6`�4�|������4DN�5�k�R�,�:����Ծ�6���5�6��]���86��,5�&�5g�5�GM5}��6.]6��0�~Ir��U�6�8t5l��5JP5`�4�ۜ6�ﴰǏ4t��6�)Ŷ ;(��iǶ�; �,
�� Xܴ���:\6 �
�y'ε��5�6��56'������m5��-6@+�w�W�S�4��e��3���c� ���F6��[6�~�5�}6�`�5�@�5;�O6Āĵ������6Ԫc���4CU�5Ώj6�o�5D����cz5�-W5P�4���5���<�F5��%�6��4h�O��}m�TU�5X#���5~�+��yo5�+˵B!e�=�����5��y� �~��>�5 ,��ľ��_6�/����6#����\˵l���ĳ5@v��"�*�B �� ��{6[���7�5�_\�@��4c5�I����4(|�`�V3d�
����(�.�]<�6��5=���`�Z4�.���$��Q6�1���D5&�ᶅz���;�� \�𤜶]��6$颶�E6�̈�9)�6dӻ6w��5q����X��;p��5
�50T#5�Y6�7$��5vx�5U����ZV648p�z�[�$���f��6�s��K�l�ͬ�4�7�6�p��6w���b���zH6޼��`��4���6Er�5�۶4}y���>6x����95���6-q��x¶�R�3���$0ζ%���~m�6A>�WN�6�ö
�?7ߦJ5^-�5
E϶Z0�6�@���V 6Jɵ��:�e�q6�x��]����6(_f�rW5�0��R�5��4��^66.�6p���-~S5@9�3�1G�H�6T>H6���5@��5�4�ϵ����,���`Ye��)#����@c2��m�6�t�6��_6m����@o��gt�"'L6 ����R���5�A�Z�x6l�26D���B� �E5���53��6X��4H�@��2j��`�k�o9��o�6�)�:��L�6|ǒ59�������a� Q�54��6���5� W��}7����*Ӷe]4�'�4T#����[�4��58}�x�ڵ�c��@$4N596W�.7�yɵ����`�5�I<���-��<����5.C6�S^�rUM�BCo6M�7��5�S76���8!� �$�l��j7��.���5�l�6�Zm��͵��͵_�=5:�6��5��.7�h۶�[�5)�<q��&ȹ��&���L�{$��|[E5�w������ ��2p�5 ˀ��W�6ކ�kTS6o*�5ڳ�6���6 *�4î5��6�S��Q%�6暪��<5�o����p6���Υ�5);\�Lᦶ҉�Y�`��7T]�51o5J�U6�^���U�j5��6)>6R��6(|���0������v��G}��Ng��O
�������նN*5"D��P��6��W5�"����6��R���^�Z��5��ܶ>
������]��{��5?4�6B�c���	3���2��P��5���5�K 4�y67еvp�6�f�51��6Z�<6�ǀ��_5�6� ��$��6r�3o�~�*�W �J��l�$6�i�6�q��2�P��魵�U�5�3$5�34�k
6���a�ֵXb,6��6q���t�5��c���"�IJ6R���k�˵}�5��6��յ��6LCz�Ƨ"6r�4�l6;1���:4���K�H�65� �g�����%6�j6��ų�u��+5�$h0�Nj�^�ֱ5r����Y�D?�6�$�5j`/6��96?�����n6�"�62���h:�FP�5�cR��)�68�V�j�'6A7.��67	M��g�5*O�6\�괸N��s�ö ۛ5�Xŵ,A76l��6296�͵������6H�%�}�6�m�� Aa6\�����J*�6HR.5?�5v ��L�G���5Ii6�����[�5n���X6�I60v5�ߚ6��'�h��� V5�&%5/ö�Ξ6�D�6j��EX5Ht6{Ķ�a�&Z�6,�^�:fö�V�*F�5��� &}6�r۵� ���s6�w�����6��63���cY6ж�Δ��@���\�~�^�6�S6�%��Bw���T4To�ξ��\Z�5�I6̘56�������5���5�o96X%n4����� 6^68�5W�60,�4n���І�6n�p6�Z��B��@�H����Ѭ�6������5��5RNص;}����6m̏6�h6*vض���ZԀ�@,
�� �6�No5�v7�;�5]P�^=͵q��6�nߵ}_����g����6�gm�֥5�N5tf��_�6 ����O��86X����B��<�,7瓁�vq	6]b�6 j�p��6�ǅ6�š�7}��ҩ���H��@�����5T�ض"nA�x)%6 �� �t4L���4�V��I�6@
$�D!^6\-������uN62�V���6��6p�u��lA�r��4���4�})6Ys�6lB`5�Bd�`�P4�hL5ঐ6���y�~z�6�u�4gV��\k�61qh6��6�r��lõf��6 �%��``7�֎������5�+G�L�����%7%:�	�6��C�+�6��r���W���^������6,����S6�����P��m��6xW~6x�6/�ɶ�5o��5��iO�5ty'��W�6�=�ڵĵq��6R��6��7hI�5Y� 7}��6��۵B�~�?k���6W3��6q��5B��5���6� (����7��ȵ�M'��_*5xc�3��/����5Ud��649�7p�6Za��e9b�� 6(
еF�]���j��s��EO�4��r���x5Bq��!X�6�#�YhL�A��lm|���7	r�^B���>b6rs%���.�;��6T���
u?6=��y+�6zCT�9��T,�=�5�0�6��6O�6��
,�5���6�x6m9�O�6�y����"���q6Ҫ�64Ԋ5�a��cr�o�4��5 ���^�6�Q6k�����W�����m�f��g6���6�_J4�
D���D��!7��=7������6�O綸l�8"�b��6^&J�b��6��470�5�k��y��,~�6��6ˉ?7��\�iF���̵P�9�i~�p�i46cϴF�6���6c6+4��Rn`6,�4������6�_�6�uT����6F��6h�굨c87�xf���]57
6)�7�C�6Sjõ1:(��
	6��I�
r���P�6�R�6I���p�?���6�	6���LE��ˍ��6<��6�&�/[�5$a@6]9���#ֳ�]w6���6+7���4�/7k#�6EWF6�\�6���6�^��a���ĵ.� ��ƌ7��L6�|6�i,7R|^5�4��7;����e�^}?���7	K6^1��3"63My��B06깛6�ʶ���5bn� ����w�6��5u67���E`���M4_~Զ.o96P�47���H�6u4���6Rh350u�6)�g6��B�Hc$�����Ls�5h1W��v�6C�6 �6(��6����J�6*d�6`Gx5ŉ���6֝7��8�6x��50Bu��u7E��6�u7�!6q���v�6��/50:�4�Y�5^Y��cM�������P�(�t6 �E6 PI�Ƌ5,R7���6��7���6�F��EI�6%�6�V�4�!��a��<���!7��6��6��s���]5��6aɫ6�Y���۵��n�4񏙶1.	5L�O6h�4�mU6#��D�)��]5$Ă6,&5��(�5(�赒�������x�5ɷ��o7W�V�p�$#��j�����6�`5�˩6��T�4c���
�B��6����̒6�f��Q�6�?��=�"�	96:ړ��d���[6��õ��N��'6vO�\�l6i��E�[6��ɵ�1Y�B=��%z���`6�sR5�
7��-�w'v� Bo�!9V��>���f�����Sƶ��16@� �1��5�̼��;7��5ܲ���S:�T��5�sB�A6�Ķ���68p�5��1'���5̤��d�`6�>��ޱ*6�"���Ƒ���m�T�'��|�6��� Al�a9�5_��� V-2�UF�t�$6�ߞ5.�6��6���5Q�/�������v�7*�\ ����!�5�ǆ5�'ض`���n ��s?6 A5�F���gͶƢL5p�4j�F��?��ZV3lض��δ�5>:ܶ�%��w�6�����´b��E��6GG'��Ꮅ.['�@���;��6�z�p]��^�6����5�>W6|�5^��5{F�6�:+6��6X7�4���7ϵ.�'7p�d�В!��?h6z}�5l�N�T5*�)������Q7��G�T<�Hr̴�U�䥶����gY�2>��$�����5��h6�6���6�}x6��U����E3��[ 춉T[�&������c5�t,�������� �����!7��Ķ8�X6-M68Zζ8�4z�V���g�[j7D�'5��6z�'�LT�5=�6`�M����n�������&5�U$���i��E���䅴�Ո6���r6��h��7��RIw5(-��̣���黴��5���4z,��R�6̝=�p'�5l>�6�b��0�k�fd���_6X]*����5�@�4(֮6�͡5�����6����%7pq�5 �$�É�~_��NT�.�K6E~�6	�ȵI�����>��������6�ޅ5 Z�3סQ5�6���엵Fƍ6J��5�+%6�VU��	�4��Ҵv�6�X���4�F�4|�C��\�� Զ�L�5`�6�*�5�صǎŶ��9����6�A����6��L��R��b6T��5�=M���F6���!7{�*���5�O5��R6����0�~�Ŷ�8�5 ��3�]����5�\�5j�.6��ʵ��d6`#޵$����صHg��f�6� ɶ����lÌ�<�|�е
W��z�������,
5L���B嶭
�X��6PtB�<^Q��A����N5 :��pEx5��=6��76��/���1����"�{�Y͗6�ѵ\-�p�w��-6 <��k�/���<6vn���=6�δ6�qV���6@��5(�е��5	�96l�S�����';�5MZd��J6p] �~�6� �4|˶ �z4��44:7tݵBr9�0xn�����	���YP���6���˽��4`���x�Pۼ�,(Ŷ��P6 K��T�nܡ6Z��6�1��{�)�4��5<�Q5~��6��5${ǵ-��6�6j�a���˲8��5`��3�g�6A��6ӑv��V?6b��58嘶`M�4>���
��5�Ƕ$��5���W��HM���
Զ4Ba�D}w�s�5h��{�D6
������� (�4�z��^Ս6}ݵ �U�=���dE��NѼ���6��N6���6��ݵ`7���H�4T��h��3?+�6:�׶��J�Q��li6�����6�Y6���� �@P��Ʀȶ��5$1_6�:��R�p6�R���K��!m�'�\56Om6��[�3�F5Rf�5��� $ٴpr������GW��5z�г��R��6��)6�)�����5��6.C�5��i�*��"�{�%�"��{�5ľ��(G/6rp�6b6��"6s�J5��5�&�5�Զ�� ��s.6�ؐ6S����X�6��1��k46�	F�9�f����5��56����Ҷf�Ȅ�2��5$�5�еd�6<�a5�A�6�#�,2�5Ǖ)�q�öʶĶS��6���4�!�L�hȴ6��7��Ț�3�~��"�E6�µ�L68丶�]68�6��66S`Ҷ-�l6`�-4�(�5T�6Lt���6�G�6p"#6$1�n������6I��5���5���6�9�6��c5o���6xc��V� ���}6 ��3FE����ȶ4@�6�mE�@Eg���5V�ප�65R~��XS"6`�`��@��ʷ6P2�MЁ�� �|k=6�8�V����Ŷ�
�5�k���{��6T�a��@����6�<J����61Y�oö�o6n��$�6W�6 =���ke��?�6�׶5*���h-7"�#�*���R��y6�?71>6�G6���6d*w�d�4�}`5o�6��U6hU6�F6k��J��6 8�3���3(���`˵HU��^��5 ?4��_�.E&�F �5��6�7N�t6�g�5�a�6s��u�s���@�5��(54���1I7��4�0n6̰|�h�����4�"7p&k4n����/15�٠5��1��!�6�`����k��\6җ#�|��6Bݰ��`4Ǳ� VǴ�}�6�X̵{ѐ3yQ������'$��JΠ���(6�3�ZY�����,+26U�M��p�69ө5��v����8�����,�̶��D���}5���5R @6ujE���M��r�5Ny25��ö��F5��S6��4@yܵ��v�xЧ5���!�޵/���S6�$�p��� �3�`���$�q��Iw���#���� ���h]p5����P��5�6��-6�"g3�3��&!"6��5x��5�'�4��܉�6�s��d�m6�{�5X'�4���Rȷ��|�6���j��Tv6�Ԃ���X��7?�6P��6�5iM�5�,K6dX�:&��`��p�5�҆6ݽ47"o/6\��� ��x����Ͷ�<��&�6׮D6 Aٶ�u
���������ֵ����g46�.����7�&��(�w�<j�6Vw4�㍵@��3v?=��sw5�GC��d�5�eB6�kX��Eq6�YT�'j�Pڻ5K}6�!��s�
����\赈��r?��+g���j�5dQ�5_�{���Y6M其�N>��QS6N-��7��5E}~5,���B�6@���6̉�	w�����mb6�G4ZPy6�i�]����
�>,��	V��Cݵ�����b�5z�3�C7�%&�h�6$�7��5O��H*��j:�v�*6g���-6�P5:�¶"�|�G��6���^5��$�6�,!���A6�6�cB������c�0eҵH{�4��T���L����F}�5H>ȳ�+�5�z�� ���`ȵ<H�52%��XM5K��67U�6�
��	r6f�_���h6�d=6���5ࢮ�,���&t��LW�d���3�
7�s�~�����ѵ����.5����6�8�5̞���8�6�+�68�f�e{Q�8��4J����6�TٶjZ7;�F�l05D�5(-����M�"�6��B6��X6��@5��5��7��/��x6���_�G���l6��T�.D����H6H��5�U;7Io�?�7���\�6�;�5^�5!�5`�-6>��5�|��NP5�G��h	���jd��?6?�d6SQ�O���^�7�/�5l�5��6	���YE��q���
6Gc6�b5�,�5�;�5H�0����6��6�6��f����(���v���26���6&~��7��'3 �&���)6*�.��6��
)6N�^�|E�5C ���e7���5���5�. 6d����6�Un���_5Ƌ�6h�c5)qX6�~Q���+���5��,6���2n2�qV�5,�5���N�5(m�6��#�\_�5�b��HU4~ʭ�	m�H����;6��j�r,�5(�������S�Eh 66�/������`�5܆��&��� �g3D��5��6�(6���5�	���.I6`�S�f�����6��ѴEޒ���ҵ�A2����5�G6���HN��2��+߱���ٵm��R�V5 =13�V�뾵��6���1�pc6�.��*�r6��J4�je6 +۴�Q���-�4�����œ5��(v,�T=��õD~Q5���+]�5�e�5*@E����<7��6|�ҵǆ�LG�f�60���(��4���>����/����)4�ʋ�0N��8@��d�FP@5b{��r�5�]5a̬6�96P'�5����N-�<���|�
4/�6�$ ��}6����P�3��.�6����/x� �u6J6�+��6{�B��I�5`�4�⵰�V6�D��c�6I|>6J�_68�H6��u���6̕c6�B�c�N�ٵ#x ��|�6$}��<��m���5(��6,��4'� �'4�N:��i#7�r6�/5"4뎮6�
,����8!@����,��6���&;��`�A4~�#5�Z�=��z����_6�m�5
�ֵ�ĩ�%�4g�Y6���6����ͺ�cH6�@16LA�4�����5�f�55��5Ӿ6�Ķ������~6D�#5������4Bڛ�tWQ6S����u�L
�5�+06J�o6<�[5�D{��f��Xe����I6��������b$��Ui�����k���}�S6@/n4pz��ڬ���%��+6Ə�6t��Fx;6hE����4��	��d5������4������6 .6��A5����?�6}���n��6�hⵑ|�5p7-6έe6�6�����b54 �5�eдP�4`&�0���%����5>6}ザ�-����>������6|W|�۰z6��:�}�ᶀ!66��V6�5�gԶ�2�����6���� 54��z�6��5�U:��H���ⵥ�5�B組�6�v#6��o��Sb����+�5>H	��R!5��K6s�t4n)	6`Zs5��5d�6�Sh�ˤ4��d���%6[_��W4�J�5�7�5���5�.��L�5��5d�]����������5X��5�g��Fu6~'�x�f���6�8�: �>ڵ���l�5�56,���@�4�2��>P�Ԫt��06@wB��ʵ����`�T4r��5C �6X],�@��\�������	�8W�5\ʪ5gH׵O��6n"�@�i��5����5?F�5�38� ����!����5|���D����4Pi�o6��?��@��
^5@�Z6�$�4����X6Ft�kJ�N@62��5�bd�A9R6 �l3��5�Hw6 A�3 t�R+��]��JH쵶�5� ���G6�U��W�4/U6�.ڵ��*���W6}���t��訊���4'��6�����5`7N4S]C��g4����5�6�4��s��=��=*5��6`tz4�KŵZ�� _5"P������l�� ʹ�
���|=5Ļ����5�d��b����3�U6g׳����5�<��k�5�Y�5�l�5~�	��M�5&6��;�`.3lU)�����*�t6�P��\�� �����<6�5�4�K'4��z��:�:��5����t����6 M���6.'B�����P2q5	y��8U6�4�7Y6�(�H7�A�4�����l�5���̈���"6�`�p��5rGa�Ë16��9��{u6@�;����5�-���7���6�������6�5.��66i�@�5�ܺ6x�96� -4*j2��#�����6(����5<�6�rt5�[6r_�6�ϖ5J�$5�I�0F`�xj��t��+~6
6�7�4(�W����5 z�� Z1��y6@۩3�[Ķ�D ��J��3˵��6/J3��˓�f�)68�W6d^Y�,�$���6�c%7*�4���\ !7#�j6�Fq6hpT��2��6��c7.7��̭>6K6	׻69����;�j+!6�	6��H���\�����;�4���4�ޭ�����6�?��N37	뵶m�m�"�G���D��l�6��6��6`S���y�5�.���,6�����}ش ߘ�H_4|�E6�=����5b�L7�6�����T�n����7���6g/�6��+5�,|6��|6E\_6�յ�XW6����<�6p��4�A�d��6S7�5�oR5P6�"������
�64%���fŵ�<͵���4H����5i0�3$r���~[�*�=�f�6�����iU�"�>���X6ִ6��Ƕx�5r�C:�46ޜ��m�5(H̵6(�%ނ6�(�[���=L6���6҉�5@,3@u��`Kw3�	m6��a�J��6zT7��}Q6t��X�5'+뵩�w��b�6�.�5���6�7�蓶b<�A/�54���%�5����f)6�����6<�Ǵ!^�6�|,6��f)65�$����x�4W�'7X��y 6�N�� C����ȑӵ�I*6��5Rk�p��4�%F��r]6�n6nw{5Tp�5*;'6�����!P6ìG6.�.6 ƕ�WS��R����:7O7�4�B\7�����"7��7��6Ќ�6$I+�NwD76�T����t��T63��6�-17>1V�kJ6�E7��`���延1t��  6�g�6��
�a�H͂7���6J7w�7���
�	7N�6pg��He%�{�6`805�H�6�\���_72�6����Ø�>P�  6BC
6ʳ��Q�h6�5�M���3�k<6���6�O�&"=6 ù�℟��lk6�ɣ6�����7�r����S���[�����4^t|�0^յ��-����mY/56��4���\�� fT��V���ŵ^]���I굌x��
�5)WD�.G���=5 ��3ٰ��3��|B5�⪶�k�5��5$[�4@o�@O�qS6�ε�&�6����3��Y>5���6\5Ͷ�ٗ5h@4υ��:��n;ʵ�&R�"d6z0��g�*�J"�6D��a�5��(60�n�8]B�]S�r�5�����5TG^�V=v�>Զ� 6ߥB5h���wc׵�86r���	6�Y6\ֵ
��m���$�$��� 6MƏ��L7LR�˙850�47EZ� u�5bD�3��[��<6�>�(��5p�ƴ u29�5 �(�^��(63o���B6��3�s���t6�)5���5D+W��A�6�� ��-u���6z� ���6�%z�$S6O8�5�)���459	X6����4
O66�ӵ8Zt���86�o�5$��w,�����6^��5H���ɶ�TA64{�B_�5᧶x*B4H/+6�\���q&6��?6�Uw�gh5���b.�&��5T*�5�淵���6���5D%�5�<m��`K�����ufL68j%4&*���t��Ψ��.L6��5���;6�?�6~)�z�M6@#��\8%6��'�z��5̀�11��� �5�*U���)��>6�K�2�6�V�5pO���6�.���+6�\��,�5�+d�].��cn6$���W�6����ʣp5�#d� �2B:�5 �1�� 56BpR��Uz5P�o4B�z�Yʜ5��2�b�O�,�6�����Bյ@����@+06�{���R�cŵ�p뵖pC5�%�5ƦX5콋6ඇ����� #�u�������z�i�0�!��h�4Z&o6�5�5�`�5��5F�5\C5��b6�������6v���|d*5|��5L�����{�5�>���7��5���3����eУ5��ʵz$Z6E�5��P,�4?e5�A�C�B���,��s6�g5i�5أ��d>�5�Z(��R�A㔶B�^5��H6���$��z(���X��B�5曍��6��ٵ��S6Eb����F���P��<�6%o5_��4�7�r���T�5�������4P�ʹ�A��\�+5w�>I�����R���p�5�̵h�I�ܽ�5%�5 �Ͳ��6�����q=6�%�5��4ݕ06 ��2D�5W�(��N�4\�,6�S�5Ď56�R'�DE���ߴ���4،����j6?ʊ�e�F6��W6�6�=6(D�P�@4����ϊ�$��4��6lQ����5�T6�&�D�	5q饶�� ���K�=0�� t�6\3�)�6\��tJ�6(1�>��$�6Pק5|�8��T�6�P6�Bws�`�O��7��0��6�#�6g5v�6�鵵Z`��t�W6��ȳ
��6��96fAD��%��6f����4��	�s���y+���H���6f�M62V'6���6���6��L�6��5���6M�C�T�5Js�5�,'�,]ƴ<���z_6>Ś5Ht?����f �5+U(���t6����H9�? T��p�5�"�6Ҽ�YزJ�5�?l6@&4 *��� 7�p\�
����5�[3c%R5N�����5��6��p���95��k5�� _5��3'�$�V)�5`�6���5`Qr����5�k��q�
6��6E8~��5@��P��5 MP5���6��E5���5P�5��_5J�m6@vҴ�sy6,��P1C6�ڴ$�e5���5�}䵦�� 俴ө5��I6I 61n4N6���87J6n1���)�4�?�4��������-޵�Ƶ���6m�4��Ƕs6���5�q�˷62��5����4����,|�t<��A�'6��k�D���?�µ���4�[�]��k?J5JnW�P�I4-��\��5<� ����5Y@6���5���5K�����6�.���ߓ5�K���U���6���5����TR���F���ʵ�a@�&!�6��5	S5�i�<��5�c7�����6���y`6"�����5h�.6YLԶd�7�m��PQ~4P���C��6�L/6�P�5��h���6|D���7�96'��6i�� /ﶮ��6���:��6Ǐ�6]a��6��2�7��������60㊶8�66Z�U��
�|WD�N�l7�,�<�F7�u�QY6]}7�#����ص[ W6�!66���;�6~_�6��5��AT�6�6\P�5Zi6 ���6>�����6Ru�e��9����� p�55�������E���5�5J��5�ʶ��6ļ�6044�,!��4��5~Tʶ���6x��X��6eD�VhX����f�ε֊�5[ж���$F6�\�53��&�i�ӭ�6���ɗ2��耶���ޭ4��5:+��y͒��j�;B6��?���\�cZc�� n�v����%�5���5#��^ݿ6�v6���r옶`��G5�|d4��6�މ��x�����	5�bA�5�Q@6,���5,���h�4���@�d�-�Ƕ�e6h7�F��/�ٶ a�Zp��4�6d����b_5�t�s�˶f��6RW�6�sS�J�浡�S�7�{5�0#���w}6��6>�16(i�?@��A��6�-J���\����ǵ@����"�_�C)�6"��58��6*m�@��4(i�6�������5�fg��Y,5l��5�]�Q%���6I�7�)a�w����V6�6ȟ6]�c6���>�����76�Ȫ���)�����g���.D.�:��:^���yö�4
�0A��P���
�5��T��3�qܶ�g_�X�y��4'�҈��<.5>~�6��P6Ѷ4[��(zb�|��5��75��ж���
p6m�&��ю5�%Y6ao���i��7���<87�1�6�Ʌ6�m������֕���|�6�۶ T$�α��/�5�2i�������&���6���n�6l&5�'4�D�&6����6:R;�� ��:6�1�6ș����5LP)�zG6 ^5B8W�t�.��� �����z������5��+6ҋr5T⼴Uz6��f5�q\50�4������.C���5Nvn6腖�s[4�B�6 #̳��,�Vn���2���5��B��m�5�,��7�5��ն��Y6t@6���5Ȣ50�4���A6j_�6�1�4 ����5\:�65/�\�S5�p86���5���66�[��(�V��57�����16���5�d"6�v��(+>6ܰ�6��?�(��q6f�_6  �ZM��s5lvC5۱�5����,��n�5;�5P�N����2�f#�+5���50
�ӂ��Mm��R���Q4���6��c� xp����H�;6Sg���;���ig��(��+�7�����`4/�c645�x!.��|�i���:�m�r�U������N��Vy�6@;'5�{�3�1���M6�j5�д�)�6x|�4�Ϡ4*�&6@�6vk�6�0e�zZ � ��K_|6�$�3��:���<�|�3�H��o 4��<�@��4��J�ǖ� ��\@5�0���p�5�a>6���6�v��چJ5D!q��鯵◸�̈́�L@����F�~�59d�5<�g�P[��L5������7��s�`AN��u��?ə�x^L��n��iv�6]�6���4P���l.68bȵe���]6R�'6��n6�3���o����4����ε�A��џ�5ʹ{6J�߶�?��hMR5�`r�&� ��l"�6q5���5�3�6+ʀ�7���'U58���Q��s�5�Rh�,q58Ě���ӵ�瀶0��4$��
�.4��96Pȏ����5�뿵l�?��	ֵd�Z����%6�W��H�&��84�6�이�ݼ5T���_@���A.5���\�E6@��3^��d�� �U3�"�5x�?��"(�pS���tص�@ϵ�ˠ�1D�5��nl5���5l`6Xԝ�y낶2�+5+�(�#ʋ���5��6�����u�>T��!4�M��^U6b�!���ܳn����1���c!�2�ϵ
���<���l��5=(������5r��5��6t�	�r�5��m����3�

��>�5��x�>]�6<n$�V�6�}�5�6��6t:5�o����5��6q'p�P��LW��H�.5�i�6;I��;���!6+�!�7}y������8���50G�5 �1��?��n��5�`����0��4�l�4��Q��6�6&��<�3���6��X4�g�6��?��PҶ�,681��X6��뵢��5Л_�H〶0����6��60:�6�'�,�m5h��5�L����ҵ�V6���5酀6�@�5��03+O6��W��w�53�6�Pm6"�����9�5���!��g(�͙�5X����W���������Ԓ�T-�5 ��3�-L6  h0ko��H76*1~�-፶vg��ʉ���)S�Ⱥj���6�_d6��5�u6Փ�`4���L5RR�$��N�	�xh�5'�촐�B�j�7\
6w�T��6q���$�5?O�5��5��60f6����:+#�~��5�4|,D�F]�4�57��7��s�0���ɼ$6\I�6伐6�M�~��Ϛ�5��ٵ;�����@��3(��5|�ԵL�N��5�����U>��{��>��5����x��6�K��06\�<�4D���#56?�5�o���5Ei�6�wR6��j�w�õ/#R6Ջ�4��6�+W6tdL6�`Z6�zѶ�gC������S��Z=.6��=�;6x�y6�X�5�8��@��5@7J57ӆ�W�7�m4���6�W��5?2.��]ȵk��Ŭ��*�y}�}g5��e� �����K6�|7~0���A5e��֔�6�2��|�4��.5��
�ۦ���6Z|M6l�2�P��5�u�PЏ���6aoζ��K�`<�6��.�HFY5f��5 AA56s�5�h%6`�6�6�;��(��/:�"[&7��^�� ���q�6˙6�C��5��Y�r���-q�6���v�K��g6��5�j�����V�$7��Y6���a�5��>7(\�6�XY����8��6�9;���6Z��{���.b����f5�~��v��4O�6�$�5�Y6�@��M��v��6���6̳϶b7��И�h5ds����7�6��5�е��+6&f6Z�5�1��WLd7�#l6�Y�5����F�6��7�J�6�g�6r�v��@O6wPZ��������4�JQ5��7� 96#��v*�5.�9��Q6���6�I��E��oW�:dD6����S�6rŗ6�I^��� gB�ޏ��sm6_���@��/�R7TO�j�6��j����7��5e��6���I�B����5�T��l�7�`�6񍼶�l[�v�Y6����T4�6X���8���4�G��ԛ6���6"	7�����z6���?^v5��P7@C6Pt/�F^(6.���x�����64M�63�̶�7������h6���b 7D�� �ϴ	���-��9���e��R ��Ge7�t{�F��5"
ʶCmA���6�]7�p��5��Y��X���U�6<�=�V�6v ���� 7����ƴ΢6����UĶ`�W��uʶ@ �5Kr?5X�)�˦7�d�rW�6	1�6��Z6yT8�X�x4q
B��o�4�o7M���y�व�滦����4�,�4��7�L,5×�6����\��%��=�H�/���6J��>3m�L��������ǳ�EA� �25*[�d~��/S�^�U7���Z�6�� ��3\���6�&����ț�6�5(XǶ�t�6T(7 � ��wk�0�ͳ��6�\����6x������cH66�����5��7P�z����)�7���6<96�]�6�|��
���6-����|4�$�Jㇶ��ـĶ�@�ؚ	6)�5Hצ4��ܿ�A�(�u�6'?�6�f�	�|6l��H鱵?��5�s�5e�2��M���S��(qR4�I�5��4j�����6�5��5{���zx"�Kg�5f�P6���05T���V��N&6e�2�x�k��5��m58�:6,����6�����m6C� 6>���y��5�8��ӟ���86�6�����������\���Ƴh�P�hF��l1ȵ����jD6?�53{�5�8�3T�H]u6������H�L��֖��X4���5���� �	�c��5j�����5�6�Y��F�hGY4��k�T�4ļ�5, �3�pb6�v5�.��.�4Ɣ���f5lǙ6�bE5G_��'�6��5#����*R6�v^5w��d�5�g���� 6��5�O25*wM���굊�����;��2x6 ��	5�榵�<������Ҵ�fZ����ʑ5nP�GH��`��5t�5�ް��;��{�}�5i��X6��5��5�k�Tھ��h��_H��ł5w�H��^5��5���6<��0�s�~X��O�u�W�,6��,5f�5�۴4Fk�5����Mx5���5
 �;c�6��G��8�f6�5åM5��5��x߲4\�4��V���
7&�6�������鍯6�_Y��: �p���(�N�z�66������B6F��^��W4 }���`6���6��j5Xx5�L����;H5�p�ߥ�6}u5��z��t�6`����O��6�ȵ۾���ެ5�*54����%S6sLu6��!�/c�ĈŶȴ86E�f��_�6v)b�*Cy5 y495�&��w�5�)X�d����	6by��N���UG5�愶d�k5^
��9皵E��Wp0����_ܛ�$(�4
��5��J�ڙ6�� �����򲛩1�pm�3w����5���,33I.6�{6T�ε��д��	����6p������4��75�0�4��J6��͵66�k:4'���V:�𴎵�Es3Q�7d�B5fRP��?�6��&�6�h�5,��j2��Y��5nN7�j,���ϴ5��6nي6;�6��u�#m��<�K��;7�� 67Gw��J�5��;6����i�6�E����6���5ru鵎��6��,7��K6b��4��&A?�������%�h�6���6�9���̆������3�BL'��Ct5b��5࠵��ȴJ�Y���5�5��ve���@�M���|;����6�����B6�M/7�"`�r���g����>5]/=6�u6�e�6q�)��� �=6XX�5z�5����,�5�f6�]�' 
��V����>�D�m6,-	6��ͳp��XN�5���4\���� 6�g�8x�4�i6VM
6�D�6P�6�0����R3�'۶����w��JA6ݒq6�14Bɵ���6墄6T豵�յ:m�6ݲ�6�V5���pv56Mr6�8P6�ѳ5,�0��~��e�hf5��55��5�f6��Ƶ���6���5�I4���[�5㵶 +G6X��4���7��6�Yf�5@�N6(>4�&� �>(6بk4��x�A�z�6��=�ID����;6�Y�d� 5	�5�=v�~8�57Ե)�5w!6X�|����5e�{��,�PHL�쭵��ٵs�6�����G��?�5Ti��?54c46Uؕ5��)����4��!��ܰ5�Y�M��6���d�v���6��-�Ї��p���t������ԁ95�5&���6Ыɳ�^�57�͵���6P;�6Zv �NM6l=�ĳW���ƶHwX6�Kʵ[,5Pܮ�6z�6 �E6P�65~;6-�6u�4�^U6��@6B(�l������ĕ�i�5/Z��Dj�6
T�6֗6[D�6l��5�p����C6���5�.X�ߚ'� ~t�Q��6H��M\6��5��#6M	�PG�6ԋ�1�����5�8�6���H��6ր�6�a0����5�ĳ6�~ �o�;5�T.5�4*5�T��0	�����Z❵��(�q���(c��6�O����;6'Q6F�F,�~5B��o|5[u66Z�޲��5��6xW�4s�#6b���F)�V!�5�<h4�e��nT���Ŵ���#����5b�56bִ5���5���6T�	�"��&�W6�+>��y@�8O6 i�쟨���6��m����4v�6�����ܵ�۵ �/���48�R�^v��1~�L62l�5�孶��J�J�6��q�p��5R\����3��!6M�,�ވ ���4��Ǵǎ@�L��6�z$6㮎�'�P��5��(6�yµT5��{�{5D�69��� A�^0,6r475k���7�z���u{�?�4�-5�$u6N�ɴ�TB�p�f�<��ta̵�5�F����'��qvQ��	�5@��*<-6'��5�H5_Jյ�$h� `�4X@74��Ĵ��5��̵��4x�5�5D`6�����p�5t6#ꥵ�7�4��O6<(�5�`5;#"��Ź4�����D���B6���5�]����6�@56�`�6ᗪ��O��z���i�����5�a63�)�8�4�Xm6�g"5�pj��d���Dj��C5ґ��CIw5|�
��&���4���D��t��Rq6(-{�}���8�3�8Q2�0�5�rٳ���5R <6�A�5��񳝋a6z�H5��5��˵�7̵�*l��k 6?����?���_�3�d���Mc��86ע6u\��d�5��|4�����5�8o5e�C5C�>6p����H�6��5�+5�w$5�T�5�&���^�a�06�
6bN��Ȭ�6�w��� ����5Pߩ3�F/���5��4���<x5�?X�Xȴx{�0����vƵ�"�5�0�6�Q5@��6�b64�6 ��5mp6Ɉ86���4N�5F�����i���6��6�ց����3iL��ؒW6�?b4 �3���5_����-�[�6IVq��H6�����Ň�1�u6�5�a�65�t��6��5P>��h]#�a�<�8��	�5P��&i�5w6V�ӵ�$��R$�<S7~���%���s����!68P5�U#�tȮ�=�|6}n=6p>��¬6D��nu�T5�1�4���6@Nٳ��(6[�6�5C5��G���k6�-�6x�5�` ���6�K4H�86��A�Ά6Z
��v
76��������*6`/6�՜�^|�5��5>{�a����̴� r� �q0���6<�6���3����e�6 s��յ�7�4���6��,��05N�"��V����A6NW�����6H��6��϶�,C� ���U�6��4���"{t�)!����6��I6�F�6>_n�ɵg5Ƕ@�>�*���H6P�5b��Nb�6�
�h@�4��.�˾�5$�走����z��� 65fX6�h�p1�6y
6R��5�ε�`�3⸵�uQ�2MN����5�)Q6��K6�G��m�6r��6S�l�@��`1T����6�{ѵ���3��6�#6�(�6M}�6V�h6�}4�"���!�5�y���:�6~�6�F�5�� 7©�6`��6��I6CF����׵�V6=� ���	�'w���#����5D��#����6,{6��7�}�5�bW���A�L��5S�m�����%���3
�s>6 q4�H�)�Y;S6�c ��s�6ʽ��,Y� .�j"�6P�O��#D6���_s3u|ɶH��59��5R�'��9��6��J� ^,�����e�4��6��60ؒ��+/��M+��05���5mH��-����ӥO�$��58S�3u�v����5�ށ��w;��#�5_~�5�?�6�V�T�=�W3϶�56��5P]���d�5�"a��&��0!"6D���/G��5Y���6��6k�5֊6�5J�ψ�5Fs�adu6(�4���6N��؉W��w�6X�7�Ϣ6'�T�Zq6����߶�Ϟ6�ǶԄ5G�6 5���6\�A6x�4����5D!6�=�6��4½��6��ε����I�6 ��5�m6��G���p���+52föM��6XG�\ T�z�5�_~�0;�5��5��06 �B�/��pP�6�e��~�6s)?6���6d65��5+�;�"S�� a2�*T6KӲ6��4JE�Q
ζ-?���|��ؘ��<�6p��6l�Ӷ#��������ӵ>õ��W6��:�	o���>7[�$�6����=~�H[�5�62�u� ǒ��a�4.��5W�D6n����+6ꮶFUt6
ϵ���6�JF�(I�K6285���8<	6�i�����5��=6F
���0����4����6q�6��P6d�`6�N5��=3�����6z��n�65#0���� ���Y6�4�6�W6\J�4 ����-�5�f-��:��5.����2>�6��6��I��#6:��6��4^�.�8�� ᴡ	�6[(D���R���5x65�X�;����6"ȉ���1?p6QM��n6��� ��2��5l�����V�5��_4��ʵ�q@�T�D5�I�Jk7�J���d��]�6Z�6�	F�m�5�6w5WY64w��qI6s����5��n6�Qh�m)6�v�5��6�!����lU�6a���:������W5!ނ�E�5�L�R�d���6��.96�/<7�CP5e�K�8�ö0K��H�O6�䀶"^7&]�<��6�:��qz��ȫ�5Į�6=�a���5{�8�蛨���&6p�~5�N6
	����5�$6+��6�2ʶ�s��s�B42�����6�n��#N[6cz�5�}N6��5�d�3Ġ�4�746��i�6w>6z�Y�8�]6n��6��w�xaP�: �����5}�(5̉z5`��e�X6̉���fq�C�
�4۝5枛5�ć���[6~s@�8L�4�m�61V�5�{c6�⧶R�õ~{)�"'���6�6��5����GY�6[J��2�6%��6�7��a6�*x5��<6fK64%6#,6��1���ն ��X��4>�D5U�� g�iW�0��6���^���p�5=�������4`���L��\E����j6��]���5�Հ5'���Ż6Ȕ<6�K���<�5�쳵�}$�t�h��"�5�j�4��.�1�����*����6��ܵ����S�	�յ �_���5�r!��^@�w`��0v�����.�75��/���5`JZ�	�ڵ��5�6'_I5�V�p�w5A%A6&�A6� �5,9��dE�6Z_�6�E$����5L��bS5x�ŵ`爳 (�5�:]6hЄ5�II5�a��r���Ң�1� ���6�yU���4	�6b>6��˶^^<51��0��4�@6�·�@�M��k4�R6.��mx��
��,Po5��z�R70�4\��5�.����0��4�.��f��65^&6�:���Z۴h�5U���w�zm6a�@��m���b_6x�5]=6R�69}�@�3��~�����T���4�J6x����@26��5<'ѵ���4�)5ؕU4F��W9H6nЮ�?r26G 6�-��H�]5�r۶�U��f"�tJ�5��ʵvG�6�,�5.�.5v�q6T�6xD4�@����=5�1�6oq6���5��D%���6�kT6K�6���5h��޽�6b�׶"��6�n���5a7#w5P����;�56��45r�6(��6����ґ��x46���ǩ6�K3�f	1�~K5HD��Z��9��f��4���П6�yz�j�
�(�:5�``��e�Tl�4r�4��1�@��ׂ����5��i�0�}�(�y�T�86�営�z�6�֯��|�� Χ�^&����c5�2���x6ܳ+��ً���5�#�6"7R���}�����D�(��5�sH��L�6Ԧ6I��6�^�����5�-�4>�~6�����P6^��!i�6za�6@��o��V���G;�N5�6��(��5Zđ��a5^I�6�a$6�)�΀+5s6z�6��*5Y�16��6�k�6��|���	���2���5�f)����54��Y�5�Ǣ�����V]5
v�6\Q�6�H6|�58=D6K/�5�u�:�7de*6��5�kʶ�)�|�7$ƒ6���6���4Ӂ6�8�7]5�t�Ѷ&Ͽ6�1�5�:綸2
7��Y67��6D�+59qn���(5��dܕ��i����n��s*�Sg?�ʝ[��F���߸ƶ�jH6�hn6U�����n�w�.o�>�v6VM����5�p�6Y�ߵ�VJ���S6�0ն�꧵fs�6�i�5�9���"�*ę5�C4@*�6s�&6:�5� ��4|6b5�97X95�(J6v����������a�4F=l���|6�$,6�\�z���6��[6u��6�6�-O68	7&�s76�#6��26�I�8�j5���5gV;�`Lo����5���0�Ĵ>��6�ض�3+���55�4P@����66�@60� �PƆ��$	��x����57Z6�x�y��Z�&�5�a6=�����/�v��6$o�F�6WJ���ҵ��.��(6T9<6NG[�뙶��ǴF�7�2�B��5��4����:��V>�5������*6�b5\f84>�6<c7���0�X���i)�6D�%5�[%��+^69�6���6Z�5�c7�5r�E6�6��P]U�����57e�����6(����n�5p��5r�,6O϶-��4XG�6z4�6~7�5r�ʶ��b6:]�6��'���4�1��ޮ6l��6^0E6a�6���6�:��R˴X�l��2�T�4$�$6f� 74�	6�X�5.���	~ϵ��6tF7W 35R���6/�ѵ��2�������?���!����7��4�_�5�]6th<�t�5Kv���Z5X&�4�_k�z{�6bz����T5�6�Z��u#6��϶�L���g*��>�����5J�6�I��2�/6�'�fm�5B�Y���i�6��5$�S�K��64&�5P �56�A�U�,Z2��h���q�p����-ݵ(l����[6�t�cj6���t�j6P�=4 
u�-֒��%6 t�*f��f+��f~4@�x2Z�469��5�[�������ӵ(-6�u��S��5x�b�Ңϵ�Cg�����+�� u6D�6�S��[4(Ƿ3��B5Ɋ5\*62���H5��h��������5�V�4�K-5Y�6 Kc���P��5��"5D	ٵ��U��S�3
~�r9s6$�6�G�CC6[L\�p�������3�	��\��5�
��ӵ�>���^&�ޕ5b5Iw��b�=zd��ы��#���5�c��0�6K����5�Zh�Fү�'Y�5�5�p����2��e�6*�6Dq�5!�8��M'6���5��N3���5*�$5(Kh52u5���451����5<�8c�6�@�50��5��5��&67�*�ι��H�5�h���q�5򂹵�m��B�5�����\�5,����a����tO��Y4ABR5�pT��v,�(�N�%5\_�67����51l�5k�6l'�5�!��Ϻ�6`��4�ă6��`����4k�a� ��]3�B�v\46��4.ڠ6�n�6��m��У40	�C�6��6���*�M�"y�5�x�h��4"~�6�KN5@J4�!66��S5`�4H��� 
�~+6�0.60�Z5d�W��G�6�c��U�)�X��ld;5�z 5L��h+ӵ|x�5�}6@�c5 B�#�6D!�6�&��|��56V���c��V�I�@ �3d��f��40�L5�5��
6`C4��!5t2��f�>o5�B��m���Lõ3�>���@ ]5���@��6���௝45)��T���)�����n�RH��0]V�$��� ���#�5�K���I66���5�"��3>�v��5L!�6b"��+�4P�۴̕ٵ6�_�ZS�6.�6��6~�7���������#����6�~V����4�|U6�]6���6� ��у6p�-6^AF�j\S��	�5�J����x6z�y6_� �[F�6q-7��9�6A��6�����:��6L�&5��v��da���>���T����Y3�	7����#�4R�6˹�6b(�6�7 �� �6^!�6���lkL��ԅ5ܳ׶�G7<�64R=6}����t5E��6��5i��64j�M/�"�,����6�%��'�C�e�&7%�j��2=�0L�5k�6ⱍ��ף4���]:����4�撶@U6�Ơ7�jV��s�h�}�x>մ(` 6`#W62{�4c2x��5�~��XD7l�-6��5�W&��<6$���IڵK�6t�~�4K�YK6p�	��u5����6?j��3��6wx!�qُ6b���B���7M��_��d�c6���	�6�2!��5
�]zm6ǎ�5cUƶ��\��ꍶF��7J�5�Fe�k�6C�E��w�5����������|��6�R+�����Z���qkK5�贳������6 /	6n$�����6�[�68x�6�6���@6��o��
�;��6j6ǰ�쏶��_6^\o6�l¶ ���h<5�X�5AwO�UI?6��j6sW��,v>�"���Q6B׍���>�0虵CD6�ǵ�K53��'*6���5�U� ���
̑6�i�6��r��\��z-�6S���`>4:Z˶K6^�ƶ��6��U6yM�5`H5m� 7%�xP"6/"���'��7�|��ң&4B��6�6'�6n�ݵ�*�6=*�6�D����5�K��bk�����&6`=7Qq���k6[�=6X\�4e�ő5�(��ם��$U�7�5�6O�l6Y�=7�}���Ԣ�?��6G�6�>��K�5X�.5"�6J�5N�
���6+��6jX06ƌ�5��� 6���6�0:�3�:64IY6�~���-�5 �K�` r6������5�I��l�(5���6 �6�Fy50`7h��5��<��t|�e46����1�4��?5�|$�%�V5��e����I�5o�5�MӵÞe���'5Z!E�K��z�k5`A�5�L��CU�4���k�
����$5�'�W��5�Ķ:��4z�p6K�6}��5�&^���5{��c5��75>�I�Ku@5'�4�q5�g��e#A��{5|�5���5���-�64d����5�4��}5�L��i��u|��o�~6�\c3�r*�^��5_|��C�׹�6��35�R���Z6�����^\w6�杵�O��˗6��
6$D���A�6�$�5��.5~$6e��j��40�����^6�"ߵ�M�5w�ĵ2Y�����5�5��(�3-�uzw4�k4ngD5}l�5U೵ph6��W5 y61-F����C��4�5�0�3��6"�C6��=6�V<6�����J5a� �X	�Z��5�a��z�6;�6*�G���m3��5����6� �5Ҵ��z�5�d50�6 2��^���D6~�
6(;K��j6������5"%C6I�{jC6�A ��r>5o6�� P6��;5P7���m��+5
6Z�)�rXݵ@δ	Z=6v��5>�Y���L6���3ѧ5}��6�����"�ĳ`��<4��k�5��6��v�}Q5
Ft�.i`66�cX�zͦ4y�+���)�P��4D?�4�6���5@<�3�]�5Qt7�"�5�&@�py���S6�[����(5��y���6�Я���:5^��5���������W6y2#��/�d��F�*����4"*5o� �=2[o6������ �"4U�+6o*6���8#���r�2��6$�H���D��3��
A��D#���6�=F�eV�5�Ç��7�bB6x�5����> ��`����+�6�v����4��Q�<���.�0p�4~B�5��K<�6�l�o_����5�'����%6��0�R,6 ��50�?3�P3f� E4�����=6�LN��O�5 pq4/�+6-䃶�x�5���nJ063#V�\ö�|�6��5Y�r���=�DH9�����9���de�0�*���6�T��6v���>P6"�6��c��\6̔r6&����������5��6>�1�|��6� b�.�7`���e6��ඝ���RTe6���4P��5°�k��4p����u�ͺ�6�bĵ@�5k2�6=	ⶹl���96�E�4��.w�6Ȑ2���?�ld��@��4[����nz4�?��C86.7�X7�6��4����5�;�l4�dO�6\��6FS��ä�=96�ɍ4��5�K��x�.��vV6x�.5BY������%�4��%60�5p�'�aе�6���@��6�^�6�4������6�\�9�k��d!z����|7p����������6>6"�}�Bq�4%ᵸ�е,
�u�62�=6ҁ6�?���6{Z�6�����µ�:���n7�� 6���T�
6,��6o^L6�s6�|�15�%)��l��v�0��"�5�l=�����jε�8�4�fd6�$�5�F�GO�9�w��[�6���5�檵P��4X�|��f5��׵�G��x_J5�O�5Nls���d�P�o5 ����7��~�7��5��w5*0��`e=���q4
�/5���679�6�4)7��8��X6���6��6��1�n'X6X�]�����@��C6C�5�7M_�6�����
|�\ք��7�6�%���U�D�^�	Ex��0���R62�a��p��*�*�����>�la��{�/�0E7��Ƕ�87,�5D;��i
7|��5�;�6�Ň��۹4��6Y�6Ҹ66i��6�37��5.����5!�$�6a�6��G7�8m��v��-ג��%�J(66]{���,j��R!7��7�Y�5Y�7�ǵ�86�2�6'<��w"5����.k6@�q�j@��#6�u*�N��5�1����:�Z�f��.�^6^�6������@�a�"�*6���3:X��@�6����ߎ5�&V6H�U5���>�x�D�<�5�6a�m����4p�F�O��Xl5�	۶25��.�4NG��v�	���f6z�=6/�3���5�����v�&��5�5�5�pO6�U6m��m5<t�6�T 6��C�M�6 }�5v����6������6w�|�6N�6Ka�`J5��:6�践���4��X���ꝴ1���#6y���Fǝ�!���H�2V~6p�6�'�3�ۈ5f��X�6��x6�D��pO�6֦p���C5pٹ4��n4�l6m���2O3�Q�,�;��$�ҵI�z6Ch>��f����-6T��4ԋ6
۶"vE6:6�4�W��675��4R��6�)��T��6  �0{�a��Z��p!������\��6T߃6�wJ6����������6���5(h6�FP6z)��(��44�6�u2�Xf�6b�6H95p��4y����N�� 5�^>��5(a4�q���M�w�6��U4�F�����6B�kY6��Z6�V�5�@�&@�5v�˵��t5�6 ���M*5����Ԫ6�����̔4f�F�G���>�.6)零9Yܵz16t,�6��õ��o5�Rq5 �4?] 6f<��27��k3u�뵪^���À�R�6tYδ d��^��5�c;��:�6�5:O�6�v05ħD6��5`�r5���5P#��-�6|G:�`߇4��H���5R �5w>�6A���d6D]4�%M5BF�5��6 ,12�;6D�$6�8ݶ�K�6X_ƶbBG5u/ŶbU�S*|6�w.��[~���4��5ZT�6X��6��S�}*�T=���6±#�/�5�W�5��N5 �5l�)����_l��A6��6�5�5v�6X�4�����j� {��f�&�е�K�5�:l��+6�#��ú���b}�l�5���3�X�6�����"5��d6p�����6�ܶ���5(22�TZ�3�5�.6��5X��6D��5��H6�,+6VS�6�3m6zH�6��033<V6��a���{5�p�6� F6�q46!�i�n]>6���&��6Nh6��V����6��5�!�6��6�D�44�&�i6�%ܵ���6�è6x�7{*�5/��p�6�~ٶ�E��?
�ߝȶG,���6pa�5�05�V�p6�5�6�D#6Z�6�c�(�X�4 ���Rgk�p��8��"�6`2m��y�6��sX$7������6�5�^�����6$D��z�|��Ђ���D�6nb62����A�����6[���2��"x5��yU6��6�cɶ�)6�U�v@5ԉu7nJ5������b�n�v6�:l���P�콍6A<6�˳�OD��������5{�R6�Ƶ6��6`LôH^�5�dz���0�L5�&7� �5�ܘ�f����ގ�X�~��l6�̀6a�}6��n6Z���-�x5j��5�<�6����?��6,I��lr���55�_��U�`ť6z����̟��6n@���x06�;�5�S5��I��IԵ3@���L�6��b6���4]�7r��K�5��E�m�6(��5�$�6���6��N�(��6���ޫ��6ꁎ�T��$�=6=�=����5�17�����6�j7�>L�8%�5�絶�e��M������K6g�F�S���ct5P\��:��wj6��6W��9�6H�86 �97��I5 ��_�G�-X���a�b��6�k4����6vMb�pQ�68���@�!�@G��>���i�7�2�6	�6��A6,�|6鍶 H�Ā7�r����`6h��5��!��,6{�6�>�6�c�6��o�=�R7���Ȁ;�;ľ�x��5s7o�v7��6p4���j����-5dˢ���(7P֡5��6��!68��6�3�r�e�Ro�6@JQ�Tn
7pX��Xo�5���6kP���6��TXN5���68*!����5����ǆU����� hѴ!�Y6x�߶� ��f��A6���ԇ��Az��D���砶R��|l��1Vl����B�5�q�5�}�6�]L4��p�_$�6�Y�6�$�5�m�|��5��5���Zu��3r��52�$��Ŀ�Nt�6��6�������!6@�W��~�3 �5�Ԃ�L��6���p0㴮0��tɹ6���6�Ͼ6��6O�:7�J>���5�C�6����ӌ6x�ҵ� �6ք_�7�|6��7�D6��86$��5�d6��6�&�<𵡳���7S6f��ؗ,6�W5��7�e��U5��36S�N5��̶s4���im��)ֵ�,6���`~N6�݂7��5�]Ҷ�=��Zm`��6�`����@7�K��.�R�Hz�5��<ͣ����6&%���O=6\ؘ5<��5.�i6P6�Ҙ�����8&� :d�*;\6 ��0P�T6��0����6�����4BSd����@ނ4�F�5 �q6�����95��� f�x����|�X�y��ֺ6� 5��S5��6�r]��ε,1�\��M-i��:�6#�X��띶��6�d�4v�613�:Y6��8��C��<Dc6�[6U]�6@���b�z6��[5��{5�5:�����A6���� P4 j�4��� �5�N6m��p�j�q^@�ε��R�2bJ���6�7������n�P6\6��Z�$����O��Q6�˄�o3̴8qN68��5 �2L��6/���Y%�D�$����J���=�������Y/6Uh߶֭5$�<����6�b�6�������5���6=��6�B5��~�蚗6�^P��6446.E���47� v��-���{�52�˶<P5�� je��� 6�T��)��6��ֶ�66�,5�d"6.]���4ji*�pT4dH��lk���x��t|6�f4�����61ʶ��6)�5ߨ�6��5��)��Z��Ⱥ�5��ڵxt5�n�5��A6�A]6���30%���5xP�5Gm��j��?��40.#�ѻ�6�<6^PK6��7 �b�~_q��ǯ5m���ص�U���m5�m6^�/6�l�5�L���"��<6riǵ�g�5�x�6������V4�ق5E�5��6ǘ��0��6�3�47:��tf5���44׻�ƨk�,���ԟ�5n�t6�	r�
�)6 �o5��>5��r4{Z�6��5
�?5q1��P:������%�4T�����0��[������|׵H��5���6L�\5Xd�6Z��5t߱5�Ƕ��0�W�f��5��T���5��8�Ȕ~6v;Q6��H���ȶ4��@O
�����,{D�$��5k�p6i��xHZ6Ӏ��S�5E��6���6����y�����5< �W�񵡉�5�0��D!6�y̵/���v�-�o�6�/6N�j�~��5��F��Ə5���6]\n6Hb�4%H�R�6��}4eW75��6��7���6�X�5Ha��8��6XT���	̵\�5Ү��޳6���5!�5�q�62֚������6�1`3wg,��m�5�l4��1���5���� �����¶	1T6
#6D�
�EZ������!6�C86�iO5�;:���_��?���W�5ܔ75>ٵT�õ��A�F���L����4i�W6
�GCi6$i��46$�qZ�ƚ5d�Ӷl��5RK5$g6�D���|Q6�Sm6H��5D5�gk�5j~5l����7�L�:6*�)"l6:�55�� ���c�e�P�8o���6��6z\���+�6�<Q5�_B�(��5�׷�>ĶY?6B�&���0������
�8�4�7`6z競��5s�6~�ص��5؄f���ߵ3�5ୂ6B5��6�k(6���5�8�5�˻4��6�߀6 �65�����49��5�o5�M[�60m���N��Y96��&6p]�6��6���5��R�]+��sME�)�4�25�!�c:c��6�D���c�5�H�����5�wt��6�w�6�&�PD�6�V5�E�5�e�5Q4�_�f�rg�5P�׵�>�JdM5�o�ٸϵP�x5N�c��!��4���,R�5U�5���5�ݜ5��W�B>c6m�%�{���в�\����E����5�'6G5�`ŵ��y�zb�6��	�c��9u�
� ����6+ty6l���4�����5T�05�m�6w�3/5�vP5���6R��5(?6��m���6�:6D�B���-�6Z����4H��E�׵�+6P�5:D5/��@����Եl���!�5��T6*�R�u����`P��R�� 6eAX6��5t�Q��<c6�fh��>����6�ٵ��6��5솫�rX�@�5�-�5��߶��5N�3�8��5��6Â/4����m�5�>6�����ɴ\�����ŵQ[�D����e�6|�6t�Ӹ˴.��5,�N�1�5"ԅ5K�6@�&3>����/�5��[�=��5b�!��h�3��&4X��4fL~���6O*��� 6i�K��^�6��4<\Ķ�KX6X�6>�����mc�5�R6��6��74�~�4h�o66���qJ�4d�h�Lv,5N�h6wz�5Ŀ&6�*5C��6ᑶ�7���6��];��i�d�45B��.Q�J_6쮙�hy��(3��A�4C�6�򅵥�Q6�!F57�o�
>���qx�������5�~.#���j5X�6U�U5��4���5:tP�߯�48�!���a�����,&������ؓ6�h5�z6��յ���.��6��C�6)�x��4�I�5�l�n��5��V4Z�/6xgǴ�{��s퐶&ڼ6�����5�hL��L���]�m�%�6��5�I���}���D4쒥5H��53-�5Qgf6�9i6�J��\Ua�?�ȶ"����u~�r�����T6�Ȋ�tx��O&6�Q��ԅ?6�z��w����#6��e�0c�&I�P�16kz35SUY6|ȧ�:.E���`6��a���O5��"6��I6��o��5��G6AY��;D�4�烶��5��B�Z��5 ��5�V6���5 �42���%Q6s�%���s�p۶�\#R5���6{w+��9���[5H4c6���j7���Y��Z���#Ƶ+��5�^�54{6�!�5�A:6ذQ6�;_��9Y�_%W6�߶�l#�_��;O�a��5�z>���6x�*6��B3�f��@�5��R�R-!5����"�&�6���U����5��5 91�<�0��.�5a*�4���B�Q��V�΅ݵ����8�׵���&~5�6Ɨ6d��� ��2[�6 &��	�5��?�hZ^6���t���&P637�$�6��$
�>��H����b�dp�6��(7P��s��6]���.V4��v��U=���5�7n}5���5���s�$6c�#6�Y#��e�5˫�6�O�h���k�5١���˶�Ƶ5��;6x���^�	6�j��T���7�U�0d�5���b6��� w�2���5�]:4@�۴��4�h�5Z���:ą����5�S�6�&����6���6�7 5�^��b�6��G7��*5��3�N�5@P۵@+�6\�X��Ea6�Y�6,����6x�z+i���N4�\��ꚬ����rh��BD�5��y��\w3$n�,�'5`{���BO��9L6�����jy6朼���5<��4v���v~)7�L6�R�rv�� 7*���0d�5�� #<�Rg�5f�õ0�s������w���H����6�5]6F�6�� � �/55��ֵ�	6���6ㅶ�����6�"���(3�,G���}5$l���[�6ʹѶ�kյ����%��3u϶C�66���6<!�5T�=�t9���1�6���5 �'��_�5�_6�f�5�6M�����&6�Y:��94 ˃6�V�5,�4�5p��=�5le�6߶�6 ]F4ꓡ5���6:2���~��2!�����5��5ك�5압5��6�h�6/�5�(�`���f(6
H�6&p��i�������H��4�/5�w6�Y�5�~����6H��@P�4V=��9?���
]6��Ѷ��˵��;6����:�6X����5@�l��ܵ`-����6#k���7��µ�ܶ�6�V�6w�\6"߶�b6��?6�i�M-�sQ72G8���/��7_�,�5 �6d�����6��(���¶&'6�M�5�.l���u6�q61
C�606��4,�*��a������:r6��0���6@����笵^�=6h�E�f��5��5���6 �t��|��t��V�e��Jm6&y5��G�������6�賶�6}O6��%��I�6�d�5���*O�5>��6���sĶ��۵��5�����6���zl;5뎊�%w�60�Ķ<��5L�"��6 Э3��صF��L�5Dx^�-<6���5�}��)�}����6��6�oS������86N��6��6�J�6�,Դ���5`���?X�j�[6D���4�6;�ѵ]�66]s�6{��6��NLh����5�]t��M��{�k6�<6��46{�'�2-6d�M�7_�%ɳ5��[�J%���Y�:�5�W�6�⮶`U�4N��6�0���#5��k�������	��A���362�6c�0�U䀶�=�6�!�5��5� 7}�+ׅ�G�B6(_����5�����Va6�Pz68��
2�5�'5�p�6�l�6�j���?��Մ�6a.4`GA� ��2�Ӽ2�i�6��ƶ�hE6�e��}7�\���׫6*xi5�S6�?F6����˴6LA6�E5\툶�NB6l���~�
5�t���J��5�e�2uk36��5[�50��6@6,k��-�5@T}�=z���޵rޑ����60�U5�^�4��y��<+�h�����6g��6`��� ��4L��6R�۶���6j�U��6����5�)�����϶�ǀ�J�6��N���V5�˼�Y�6�R�5��\;y�!�6]�g��\�6�>���gN��E��9���E��6_|66W��kZ�6�I���&��Ο��m:��"\6D�5�e��i�ڵ<g�6��!6�0�i�5,˴a�Ŷf�N5��W�ƹG6v��6��k����<9�5�KV��"6o���3�5��6��ϳ~u�5�����{�6���~e�6�����|�6�7�4�K�9S�6o�w��6�#��4�5���5�^6�^T�NB$66Nд��}��˯5���6@C4!�(,Ӵ�� �I](�P�H�"���	)6�8��Yx�4�&6j�p��;G�G����>~6��3�*6i9$��ض��H6�S����B6^��Ri�6R�<6��6hs�6f0~��=��Е���g�6�� 6:�v6���6�35ՙ�5�}ⵯsS64O5 	�68ڵ�:6L b���6` �^�6P෵�Q6ɐ�����6D|��]Ι��Ų��ζ=wF6"��5��⵲`���5�?HA�.#���]<5�!�E�J�^��4��|��?5y����`5zN�6���4
�o6�쟶��쵪	�5:~�آ�5-�B���jO
69�5��f6-`ڴft��>�y6���`+y������6�_�4r����2�����R�6�X6��57���ZrD���@�� ��,��%L�r��6�S㵢MC5�T6+=A����5�5!Wu6�6��,5�J7;k۶�m��<�6@V��{�Pg�4m0�.!�6H�5��6�6˧n6�H6H�6�7dx�мf6��4���6�~�p}7��5�;*30�4��v5� t6>���c��4�5�Z7H�6����.-�se6l�#5:<�,Wʶ��6�z�l���p�::O� _�(e�6RG6\�7�����6rɯ5jP6�≵R�̶�	/��p�R��6M7����5���ܵx5̍���6���2�4�5�,������,�յ`������6�l�6��4���6�����5�b�5;y �������4��4���i���762�T�j��5;,�6q��5`n�Q��5��32�4�=5ÿO��\N�Z�y6#�ζO�16B��5 ����Q5Ru�5���m����4���5��c��(e���>�Uhv6�q*6C��Db6�t?�0���"���#��s~�6�1Q�H�~fQ5�K*�� 6^L\6H�6/I�6W��5[Z�5{���L��t���5��&6b��Dk��=��=k6�5NR�6	�A�T�c58��44��5zrҶ4��4��6c�l� +b������,�60�6�S�5��r6� ��PT���50��Á6%����	�5��&5tF�5�f5��6*���x]@4X���$6d������{�Y6]T���{�5^!��\�~F���~5 �v3�>6&��6'����6������L�<zH�p�5] ��ø�A2B6��ö@�������M�96p���/�K�~���H�V�ٵ�u7�x\�6&�K6�a����ŵ��W�Z�ص +x6���3V?���#@������926 r����v5.�6���r�c�6�w�lyp�*�}��^����6P�D5u�6�?�|i�5�105�T� �6��05�M�5�D6 � ��Q�5�}�68���"&6P/������`Xӵ�L5������O��-��B	5t�D6��F��h6�ȵ��46^���'q�v#|4�(׵h�4�5�"���_�6�z6x�6�{��5|�4��s�d�o4b�-��5���@�2)q�@ "���m�����c�6Q�$6h�����68$y5߼3��R��>��6`S%���"�϶p���`0���M6ʊ5V�;��B468&�5���5p�4��(� 5�#6�����^��5S��&6����<�5��~6�����/k5|��`~ٵ��56;w6�\�5�d���~���k�4ਾ��W�5�Ew5�	�����x��5����\!����6X�K��68���*�K#�5>>���aS5v"%6�!ֶ���5�=5��6@G�54o5��6�f���D��;,5�1��k��5���5��e�|�5`N��K6�6ЊF6����ޘ3^t�6>���tT6>�Ŷ���6 $^2*�-� �j��S.5�8v6!�6�gs��.6p ^�\sŵ�!O��<a�<�o��5��Ǵ���4b���p���RC6�(+6�7�6@^
��&���Z#5�x���k�(%���-�V�3�7�&6��F ڶ:��5hɠ4:���66��X����L5�`5�b��B��4�Ja5|���(�5 �}3�
��%���xmo5@lu3?�6�b�3��O4`���'�����a��u%����׵H�k5 cʴ�]�6\�µv�A6wD�6̭��Ꮵ�t[0�`C��{��In�� ��3Z]�6ꢵP7���5���6R�"��:M��?�`�]��nf���F���"5=�5���6 p�4)��5|>�5���6 &t3���6���6:#96�.�6gF��a�46O��6,J��pY6�(6u���PBӴ�Q6.7�Ȩ�P�|���I��6�4n�Ǉ�f��5 ��5@&S�@}�3�q�6��&�X^��(i���(N54ǵ�����;46����g�5����6�,�D��fﵐ�L�l}6�l�6�J&6�o�zM��ֵ���hu$��p61t'��>�6ꄵ���%���4��B����6����]���k�5�V����5�=z6|w���G5�hϵ�d�ag5�3���dǶ3|�v�56&���<'�B�0���;6P{u5�¿4�6f?(�t�6�1Ҷ@���d�l6Ȟ���<��-���z�5 ��2���6��6���ͳ�5��6�U�5��6�0ʶ@³��50��4,F{��W6E�/������T�6`,����5�_�J�4��]�5�y<6>�6rL���\6̃�*	����b5fn	6�hk6���5�tI6!P5҉e6R��5D󶌿�5 >}4����De�etJ��#�6���G��?��@൑j��?�E�0C%���-6
�'�@H�4�ow6oe6j_e4@�o4��6��62*1���5>�5bs5��5�.%��5R��6�6�� 6�k��$'��6�5�#��	�5�B�6*��5�؅6� ���b���5f�V6J��4���5��O6FP�6��*��z�5Ҍ6d�ص�76Z^
���ѵ?P���ȕ$5�59�Q6l_�4��
6
e&6�iR6��N5��5t6�V�5�Z��P6�-��c)6��5�K$5f�l}6�7��5̂6N�s�&�&�4Gܵ���5Tn�6��s6f~Ƕn�޶/�5�8��,06`0P4�0�HDƴ,R�5��
�ؖ��nc��~�6f�5��l�MLB�0*+��r�܉J5	6�k����4˼7����9��A5�ˠ����6X1ö}��5����Z$յc����5|6���5���5A�6����56��r�6�Ĵ��:�����X65!Q䵌#�5�m6i�nM6��ѵp���y���&q6��5=�)����5v\��6�G�5☑�ܲ۵R-�5d�_��u-6W�G�<�L���s6'p��ٹ���*5cͭ��x�5��5�Ś5M[�5�tg5\ѽ5Ȩ�69�,6W��0��.1�5�6p�[�S�ڵe���v��)<{6�}���a�4�rŶ���5H�5,�f6�۫5ް��õ��X�R��5pN�6�$��r'6�/�5��5@@�5�>���5eU�6Y>�^R��Q;j6�͈6@�\3��)6@;�����2�.�6�q�5�W!�����/�F� ݨ�b�X����5�A�5Q�6:���A
��r���	������K���3�6Y5�59Q6 �-5H�q��P&6���@p����5�v�����k?�6��v6�.�5���5Ҁ��
�S�f�6$��6@ʉ��6y7l5�B6vj6~��6��O���7��G6����&�F6�LU6�ȼ��C6(�4���6�t����5�8������=�6�T6 	=5/ܲ�}����㵤��|$�5�y$�\J�� 5�4<־�Z?~6� ��
c����Դ#w�6�F�4Cl��K^5��5��6~(6�V6ٝ6p򟵒��L3���h7�5���5��S��$���Գ|_�4�G�6���3>��6�b�4'f��Q�@�=��Q�5��K5L������3����Jj�5�u=5J�k6{��P/,��l�5�16��6>c�����4�A6,�W5�A�5�:F��q�5�H6��6���6�c�6�u��e�"6@H�5:Q605�� �����$6�1�Ͼ���D�5��N���Z�5B���z@6�H�6{o�����6���0�*4�ֵ(�X6�T�����6!a?�������N}6�@����6 Fs�J|�5"_ŵ��ڊ6��U6��6n߶5���`��8?6녶�׵�G�6��B4,55�<>�����w96����@�2(�q�$
�������6�=�5Yn�6�M96a��F���%�_��6\4�54h�6ЛZ6�ɶ��5
�f6ή6eB���9���5���j+�b��5�F�4���6?#6\�ŵ�:6��"6�J	6�K������Є�൬6ݨ*7�����4%�5�7n��{�61�u5�o�љ���c7�b4�l�?�����0N�4V6'ئ6���>� �6u���Bu�����6�d�4�˦6��^�l�k�6S{�)���[6�M��05���4@�F40���g7�U�ip#���ٳ¨�
dC6 H��ԬO�PB��U����C��ꐵβ�5�B7~6�9��,5�y�M���Ǵ\���g2���<5��6n�X�VnŶ�=��$S6�ӏ6���"T6�p���779+'��>)5���5Ʋ�5ۊQ�
ŏ5��^G�V�6:����鶥��C�M���
7Qy�5vf�����6�>�6�#�4��6s}�6w��5A5�����t 5�cf5L"�*���/i5P�ε�� ��f#�֕�5���ଏ�X>N6xr����5d���҆�Wf�5�Lж �K3���4�qh��2����u6 ��hnw6s=D���¶���5O�!�{�G6(I#���4��05��3�v�5c�5� �ɜҴl���I��D5�	����ux�68�͵��洖�/6n��6`Մ�D����ғ��OF���6��Ќ��R*U6�!�4��a[���*ε�t޶B��5L�5�����6�X�Ρ�#ɐ6M(K6���5>�	7��4��h6�{�6y�4��j,�RP���%6�%���޸6$��4n��5L����x�66���6��Ƕ�f�立6��\��P6`�$�3j���z�/���6ڝ�5��W7�S��͢k6>Y�\�Q�~��4�o���Z���+6�L���k�6�b���J��/*58$ǵ ��6��6����6�� 5��w6K�6�15� $���5l�㵻�u�����Pɒ5#Z�56U�6���4�H2�Dɀ��O�@?�4Ii4�{	A6�m6ѳ�5��5`\6�k#6��۵gE����6�K6`���4.�6�/p��q6�����6����6tO���7��o�.��$l6ȝ6DX��*��6�������l5�6��c6X%��46'��w���B�3B�7�(����s6&j5N#��)m6}�6n���4���5XQu���86Ko 6�P�6%�඙b�-6{t!���V����5�3��,��6�td2#ZN��6^.N5��&6���6�.�6ޯ���@����ӏG5������Y����46
f� ����!7�f����"�[Ă5�2=���~6^	6P��3�d���06�\\6寥����5:O�����ῆ5j�5H�l��Չ6���5�6f6<;����6ra�6`�7���>�5Zz#��>2���v5���3�5��l�6Na?��C�6=��68��X�5H����58�E�m}Y6:��5�/1�p�0�V��6�����\�6�8-�D�Z��8�4}?C����6lʕ6�>(�`��6Ǉ:��G�6���5�i��6�U�5�k��yj�����d�4b��6�K[6�4&6a�+<6�P�B�5�f6<�(����6x2�4�)6��5��*
6�L���\6X�5?�o=-6��6̕�5�9Q� ��
�,6TU�5�Wh6^�3~��6al��
��|���BY��'64.���&6@bf�	����+��蓶��F6�m�6�ǁ5�W/7}�6\�R4(����Z5��f���i4Xwb6���`�6���C�i��5Բ�3t�����T6�0���&6���5ZP5��n��:1\6����4��6��г9v�����4f ��}��6�s�6�X 6��\6'J�8�0�k~����7���6��O� &�5�7�7�I6#��6P9��K��5��� �	�R�����4�R7���6HԤ40��4~׵	�ϵ�K6���6�68;���p}6��j���{�c�6���5�h�6M.϶9-�5 ��6jU��ǔ5��5���4���6�!6X1~6|��6 닳�a��(֒��j�5
u�nb6�R�5��l501�5i�6�6@f5��M5�*��5�_6j��5�)��xt�6$��4sГ��=��)! 6��6��ض9Ǵ�'F����6z1��ʘ����3,;M6W�5fHF�P6)���ݠ�{xM62b��bj	�`�U�~�X5�G\��F6���j,6;��5��8Ak6���4b���K�7K96���j��Q򘶍;�5�M��!����E4%�A�����4k[7��76�6@�:�� �6��5� ׃�ȩ=54�#�u��6G�_5pl����8����	�5�<�6w+���
V6��ض ��B�]���T6\o�1�h6����m86��Z�H�m6�W��jcz6��S6��6H.�4PvQ5��6�r��S��Ep\��
����ߵY˒�쮏6�Q���
6Kn6��5k�57Pw6P��6��Z6�$k�f�@��4/���&�6c�W6,DM�o�=7�\5���Y�16|}����15����?�<�6R����(6���#�4J*�3�|��f߮��4�6��{6�����T��v���CF7��x������76P�O��9��8��6�as��@���I6FI��j!� J�4ЎD4�M�tB��"���-'�6ȟ�5.�D7Q�7����l-�5�t7`�7�C��m��&68�x�k�06T��[���n.�JVͶ4�����:�čK6�.M��.�5�L6�䇷�3D6v�ڵ���(�V����)@����}4@�6_�"���ض`�5�5o� �3З�6 4񶼏���5w6�� �\��5��_�&	�6[�g6\�5��6ԃW54�w6������6�%6�꛶�/�6խĶ�37�Y����U
)7|�=6 l���������6 ������8l��P6��T5�L6�C���5"NJ6�It��.�6�7� ���i)� �%�-�6~�6d�6�*��<�c���.4�9����62�ѵ|���W�� 7F��Z���)�6g#W���յW��5,3y5J��5d�4�6tT�����ާ�6 P66���\�6|)�5���5 ��?�T6.2�5{�{6q����-���6�/���㶨Ҡ���s�������6dV�6 -�����I�A��$Ѷ̩c7�����=3@��N7�LV��}�5��|7o�p�5j:6ny���I6LŜ�j5�6Xߠ6��pAж��7Z�'7��?�J��6�������_7:ۨ6�ǫ�pq�6$ҵ5����H7�װ6��w�⬯�t>����ж~�.66�;6<�05��6Ŵ3��;�6��m6��^��6��Y��d���0�� ��P�
7�����m��7^q�5�����6��̶���!Z6_���6L�y7tu����i�j
?5ԏ74 �L�)�p���ɹ� 	��f��5�,����6"��5�I�6�N)�6<6��6����0���"6�6�y�>q�6"���}��q�6�V��~���<6kص��5{㠶�a��DK��,����$7�0ж`C�ؖ�?��H^�����?%�(}/6�e�5
V]�8����5EQM5����
I>6(Lܵ��6�0յ���6cg�"ں6�����x��.Bn67�F��,5@H"4)�C�>���Ƶa��Ph�3�Sе/����"j�37���6��7>N6�*��`�6�w5^�H��	�6�G�@�4 �6 9a6b�p6O�S�Ѝ�6OǶh�e6Cw�6*�����6���5���5�N�62#$�BL#6��p���5Z�5,{�5�!5D~ʵ<흶��<�څеI9O6�����]i6��z6��9���܎��(��6� 6b�=�������&5��:6�@�4��ߵ ]�����D�P 34�4�5T�쵔TK�j�K��R��S6�j�FĶ�q��	����U1���5Dd ���h5�6SC�?�<���o��' �@|����6������	�@��6�0��B������ٙ����5X�e��fS6y��5�s��e�86|1>� �<5�]X6�Ȅ���?6��ƶ�&��^P����(��6�iM6�Kv5{�6����HT�� EN6rδ�f޶�%���O6�v���}�6���5j���o�,��2�":m6��˵��L���.5*�u5�@���y5�1���.6���6��������6tt�4�s��1��5�6�Z�b���
�� ��4_006Tf�4w�K6�Wq6��5�]�5��n5�迶̱�}x϶I��6�����0<�Cl@7�h6�]�9k�"7:���gG6�Rb�o�_�n�/�b&a�WHj6--��Qc6����<��`�ǴJҲ� u4l�1��e5d
2���5�е5(I�C� ��⫶/�{6��7J�����f�*����?���6�[�5��
��5����jȸ5���l��5��!5�q���}T3p�O�vH�6`�ִ�I����6��7��\6�rh�5x���'��ܽ5�pش�\$5:g�5R�
6�+558yV��d?�H���кo5��^�F=µ槶c�6��H�
IƵ�����ۨ5�6�w"6H�4���5�@��(� ��iߵ~6(�
ߵ�	�X��hjm�	�6�褶�:�q��0H�6�A\6FX�)F��6�d�iϟ�L?ߵ.�k���ŶV<���>%6[Ӗ��W���ҿ���l6$�4�k�6z�Q�����*c6�8�|��4����8��H6��˵�lx6m>P�z���Vm��.T��7��� t�4�=	��k�5;���p^6�D�M6t��69�5[޶��5���5(�6��6�h���6�Ϋ��~�6ќ�5Q���{�5�b�J�/�Y�6�=���;���W5�s����3�>�6��s5�1�P�+� ��2��>6f����A6t�)�(4V�p46��5�A}6��76Yv4<`���6����M�6�'6�W��a5q�x6ʻ�6P�)��\ 6M�*��`5J���zh6��86��6�;�6Y55��$>5Ԁ
5`��4���4=5B�P�0:�5�>5��S����*��Mv�:Z��H�e6pP��vz���/�5P�j��T�5�E��`?����5x��?4 ��1��=�z�E�l%6tM5L�5�@ص�'*6-O26���ꪨ���5YJ6��6�~봀A�4A�16@Om5�v�$�е��4��6H�a����'��5�.εB�5O��5��2�b]���0\4�b6X�u��k�5_�c�`*��pP�3�x�=�H��t1�P) �:m5UvT���z5FV6����s5��?���|��
h�j�06I�5��S���I������86 JL5�16�M�4�/g�R�����5A�ϵBR�Ց\61o2�n Z5>�5"ׯ5@K�6#U�5P�e54��W;�[_��Iᶼ��5TM3�� 6��5`×2H�6/6)OԵh��4W&�����������V60�5qk���z6��5^1�a?6Y�35}ח5��i6�K�5���5Lݶƍ�5�fu6���~�5ۭ4����,kn�*��5w�6�`�5�慵w��6W�{���$��f�5�(ٴ��7�����ٯ6윘6�u6�?���26n��5p��5�����8ϵ�>-���5?zZ6�|;�늪�VxZ6R��~G�(��4�Î6<淵�-K6������@�մ���g�5x�6+�26b-�	����K6�� õ��7<��H$5��!6�d���k�Z��6ƒ��2&~6�ȵ��ڳXM�6�\&6���6aj���5(6(2��,��ڠ���_I6t{O6����<���9�6�������a����.6�x���MR6$� 6t�^5FP����}��Ӄ�Z�6:��6o6�J^�b��5+B���(6\���.˶ F�3,۠�p`6X�6�S6��յ@6���?�$M6v(�5�NV5W�5Z���DÁ5�m�5e�6c:��b������~����6��ص�?����%7���ET������D6���.^ٶ������ζ��X�5�\5R @6�b�6�o��&���5y'��=��(d��"Yc���6̛�5��2X���S�5�D�6Ɔ<6�p77�,��O:��Z5�~�����&+�9�5ROa6�@��X�5��޵/�6LB�4'�/6��޵5rWo6�$z�/<�6`�,��4T� 5�ޒ6.�1����6��ԶF[�6O>ض�z"78�r�0��4�vp5�������6Z�6�⻶b��6�H�Td�9��6C�6�,O���95|ױ��7�@|61X5���6�,��#6  �nТ�V���ʄF�H�5贶ڑ�����67��5ն��6|Gض����^�6CI_7���6��T{(5�w
�p	�5x�>5��	�P 9�0��9�6��]�2s#6�븶
����a�x�6T�5k�����l5
����6�i
4��O6���6+�@UG5H�B��f��	��UU��m�9-�58O25�Fq5B���ŧﴤ&i�A�5̃��@�pz.6���@��5�K�5�痴9m60gu3���6��5o�4r�&�W���D����V�28S����6��!������샶�=����q6��p7�ت6���R��>��5��������<)��D#��t�07D"׶�o�Ӷ5�k6��嵑�6��p���5�i��ʹ7� �D�Ѷ�56�AT6\ٖ4|8��ը6������\�P�1�d6X�7@�2���`5�]���I5[+�`��5�J\��F>5<��6#�"6T�ö�i��'J�6{�6���7��K6��K�蠆���Y��Q'��?���S�����5V����u6jtͶ��6q5Z
f�!�n6��66����5M�5�NI�o�$6���r�6�m����68��6�0�6�ŋ6�	64��5�����,7���6 �5�3c6p�6�F�>1�6�h7$R�cR�6��,��\ƵV^ �+�6h��6)7�<�j]�5!�6XW'��d�5<ey6�J6!�31K ���5t� 6�䃵����ҿ޴@�Ѵ�6���6��6��6gq6郢�滋�<�׵ԛ͵��C6:H�5ZZ���4��T�϶�f6(R�6F�69��6���n�6\ˎ5�V@�l�����6�
�4�6�%��ϯ��Z�w6 �_��X�5�2�����6R�����3>-�Y*6�϶�;�3F&��P��8����5��K6#5.��5gSٶPҤ��6�6î�h�=6e��t����%6G
�6X<4׻����$�bȞ5B"���R�6fcL6���6�8�5X�ɴ���)4�4k��N��6U�c6OK6z�6�)p�~�59g6��6Ii�5<��6�G���'6l泵NZ�hn�6 >�2
���r��\X��ۀ�bRk5.���K��6c�5��C�Щj68qf4�Z6������S`�h0ڵfK�6<��|A5�K�6�z��$z5�qR6�N�#�6�K%� �5���<5��4 ���@m5���6�W�h�'5W+6��6��6c���v�_ֻ6��c�
�6XaN50�V5c�����j�0U��6C6 iR5��6�uS����4����&����ˬ�Z�X5�"��;�6�-� ��f��69����5(�5\]M56�6��"�6������3�m+5g��xs�����4�^�5X)26,��4��{�\��5���3�5��tl��z 6���5�ix�5�q646dc�� ܵ������DC�l��8.�5�髶�������5'�~6�7��t>4׫*�d x���� !���b95�:�4O"h5��a5hE6�eo���_ִ�0�����pO5p�4����������$� DA��&6��'� .���6 �V4J<���55V6��r�~�������ǵ�Z�5y@h6�V6q����� ��:16-zl6 ܨ3���5�K5{I5�n76��C6���5���*}����95h_6�赞�Y����`M�^�ʵ^`68���輵�1� ;5j�ܵt&5 "u�w=��KɶfK"6��E��6\Gg5G�6��5̋<5A��5жi4(Ƶ\��5�ݟ���`�lǶ�p�4�H84�#X3���;6O�6�\�t6�L26��۵>���_3��n��J��c�+6v�z�ܵ�6�&i�\�?�\n�5 zA5`|4"����4><���*��kȈ����pε�Ƣ5��<���V6;6���(�5�z�6�u�6䛵p	��O��5b=�4��/6��65�$^���$6�Y15$�:��4*6�Gx5Jވ6����4.60�H4H6%��5֜50�5�8� �����յx��6�߲�06�����05�} 6!��4�4R�X66�t�6���5�w��d�5���9'#6� ����d봔�4� ��H�6��50"ʹ�W�|%�R<���G5&T55l��5l�J���~6�7����Ҵ���5�C�57O 6�7�|=9���T�I��~#���i6��6xq�5�#ȶLj�6<�T5@Ͱ6�!�]�k�� �6��Nj
���6\�� �76��ص|�6�ٿ6�/��=n6w�"��)/6�!��r��X4���24����S3)6})7ز��O���q6�?�5��96��k6D]����n�5�����#t�?$�5�〶v�e�<��6�Ϧ�Zp"6|��v�j6#��6`�`��϶�ݞ��*G�Fc��b5M�62�?5�B�Ą5"�D�o�#�~�$�0q����X��튶��I��T�{/�6�K�60��5�7��RMi���6"a�����I4�y�6�Uw��'�4\�6�46��`�H�ȶ>����b����y�A�_6,6[o�4?��5��S�@�ᵴ�����~5��6����~6����[9A�RFN��g޴�G�6�� 5^6p��&�^��]�6#��l��5^ʥ6NH��r�81�6�ܠ3���6[�o�3f�Jص�6P����W�6�͎48���P)�����嵾����h�6�ʅ6%u�%��5�}6��r7 ��2���6�~��g
�f���6����ۊ�5TP�6�(��3^����_i6^w7*��6�*6|�ε�y�4|��{������.���5��+5�Lܵ�Oj��4�	ȵ��P��p�6IX?6��x4غ\6�[�5E��6KlB6������C5 o����u�����DN�6h46�$�����\6?�'�,R!�5��6����Xx5��2��6�β�5��5��6.f�{&���:6�? ��J5�]��75�-ڂ�nU/��u7����66(}�5p/�6����h{6 ,� ^����_7e�:�8�;5k7�ߵh�̥6NwX������B���5� ��V�5 q�>�6�X�6f~2��,��ĵ� !�?��V�5Xw�6D�Q6�r)����}�6t��5�v��0L�6�ɶI'06@�=6�\��rc��i�6����}�dtI�֕��F۵�!�5��4syB�v�s6|@�6X!�`qK�Og��4��<��5l	}�2~�6���Rф���6�B����v4~
��ݴ���5�ꭵ�Z+6�Cx�����l�6�6�Џ5Q[�W
6\1���C6仭5�w*�vm�^�S�6���L�5��*6��¶__�5��W5��F�B�.5 �/2+5�i�6
!��6R��\��6E������Ե7Ӂ��5b�6�]��_}��X���剴�53P�6v2�@!6"���]/�5�^-�)�X���)b6
'6)���/l��[�� �5��49�6���4HY5�	�5��9���B����]��M%5`"D5��µ�h�4�H��ɵ9�,6<7��4�5|z���a�*�`6��*6�BW��<�j��54��4��B{5P�[6�r�������صPe�5
�55>�6�P0��/P5�H�5���dfu4��^�L�y636���Y�40-�4�#�����5"�~�$#��YkڵB���B,6jz�4%�T�؊�5��o��f/6�=C66�`�<*�4��6
��5�&/����a��|6�y�5�\��u��H���F6#�l64��5�^�5	6z����a6X3
�[[6Ŝ﵁Ǆ4��Y�D���q6m`��7�=��R�6�����ĵO�6�/϶�#�4Yʹ5�:��)��6���6�9��r�5$f��=5��k����k~6o�/6oE^6L5���<� ϲ��Ds6��R5�&'�gyL���2��5��>���B����46S�b6!6�Ѐ4eд!o6PP6�c5�����ҶY��50�5��6�Y �i�}6�iV��-B�|[���d������5|�L�/6sGM����5#�&6���5��b3�}�6�%�����5�ޒ6�Ѷ�A"6O�b6���% 5��b2�6��I�4F��`~U3:㟶ʍ�5C�ƶ��õ�3�5�7q7��r�e6��ݵ���� +<5�{i�.�f���J�I@�6�Ԃ5�M�6��c��������q��q�-�0�Z����5��[�`IV4ް�5�.6sqR��M6��5�S�������Ւ�6��5�������4*$���n6^�N6�D6�?D��S��0´\@���q�6�;2���@5��5�O�6�����6
+n5���a14p`����ö��5>�G������<��!����c6���8�6޼��h"��UY�G�5n���ѵ��-5�D�F�#�������/�(�5���Tb�5��(��?��l;�5�ML��)�5	�0��{�5to 5�����Y�6&i�5�����g�����4"�^6M�-��|6�5�5w�6�'�5=S��&V6~<��ux�Tx}���I6�.���ٴ]ު6�t�5�I��HY�5&ks6��6��+6�~6��f5�"���5�o5�G�������援2�6�Hq6���6NN�5�EJ���B�w�6p�޶���x-5g�R�5t�6��^��<�\4��6��L6�&6�1h6�b����6���@N�4�bk�&�D6�ss�P=�'m����d��!��Z"� �5���\��5�]��$`�5v58�Q4���6T%M������6=�6�x~6��ɶ�����n�;����6}�ĵ�535p�p6�6�I����5@e泄ɨ����3(8�5�bL�������-�����@f6Pd�t��6�673@�m�����g���[4䊇5Xi�tq^����O6�o�6Dk���6\���������������6R��6I=}6���B�ɶ�HO6�bQ6�M6ã�6���5@%=���]��w�58��6@� 4<N�TL�� ֥�o㐶�١��t�� *��\��3�Yܬ5��X�5Q%C��^�5��5�Ec�r��*0w58Yd�.�N���7�xĪ4𰵈�5olʵ��m�݆6u%�����6(��6��6~'=� �5���48ȝ������5c��ב��N*6(�95�F�6^�W��<(�Cb���w�A�/6[����*���e��l��
E��nͶK�$��+36Ι�
�$�|�96x)n�T�����7A��zu6d?�F;H��*�6ԫ[6�����i��*��5z�5��V6�t�@�,6݈6|UD5d��5�Ɉ6a�BC�6P����������3�|6i�n���5�\�4�s5Tt���S��(~�Ց�5�ں����6��˶X/��\:6�]q6�̐�t�67���k�.17���u\Ͷ�,6�UT��\A�`��6v�8�'6�ç6���6dT�5��g�C����@G�4��յĪc6/"7�!״ڈ	�=����V7/D�6����.6qYf�0�17H��-O6̠��K�ض"պ6���5 Bd2�	x���-�'6�+��g��u����X��4n��b�-6�~�85Ú6�*��K�z�6^�����\��O�6,�(6R�ֶud6~�6�>W��/:�Yʹ���6\+"�\z�� 0�k���)�h�k�W47v���O��`Ѷ��7��H7�"��K x���F�+�s6E)���,��}����N6�>�6���6���5T��Q�Y6R6��y7���5 N���+����5*D#�~��6h/5�?�4@�T��J�6
�������*+�~/f5ہ�6F�5vN&����6�037u&�b��6
�5�ɥ6ͻ�5��	�ؖ6��4�a6��6��6�U66��6��5p^�6Lh�9ڻ6�0�6X���껶�x�6>�6hb���^�W�642�5ԶL#F6��"��46�K�}��6���4�%a6���	6mbm6}�l�@ό�������V�a�7<�	5�V�5�[�6��5�q �8r7t�����ԭ��|L�5 �M�`X�4Ps_4���5��5�X7	j��$ ]�,Ԣ5~��5�/�4�&�59��6I����A�5��?��>����7��v�60�4��P�����k�6V���d=7>��6W�t��X�4'H��J;5�\޵�]`�d���<��6�bo�$i�V-_���״�I��:����Z4����i�5��&�������-�(��5���6㤵h���]s����4��T�5̣_�D����#��>6VXϵ-�7�(zA�_�յ�w16� 5�Y�QC��k�6U��9�5~�y4\݋�*�5�/5d�����.���Ŵ�z�5Z C��H�5D��4ju5�5�6��?��藴��I6`mm�í���J6'�µQ�5J�r��G���=6�=�5�S�5?��4ά	���9�@�δѽ��6��"�{A6(ဵ(H �D�U6�
�z -�
��p+�5��O� ib4@��4�샶���4��4��4�j!6�����7g�5�v��0�t�B)����5vڟ5��ɵp�W6�Sy5�6��
�m��L#浌�d���,5 o�5b��� �hC�4�ݸ4\g�4�ι5�Oٵ|(/�����5�[�p���Q�����*6�bj���`\5�����[%5
�'��һ5p6 6;�����ؒ!4$l�4�:N4]�d5|8*3d���7��D��e���	 �B&��Էִt\6�I;�TJ6��.��K�6���4�,52�U�LҴ�q�5ڊL��@�4L b��Ԙ5(�Y6J�6��M56���u68,���m5ж�������6��[5s2ص$95%qӵ�n��ā6�8��lZ�5��Y6<A5�����4������;4��"��]����\�"���@�5_<8�ݐ����5�d����}������k�6�N6�v��V��)ڶ!�6Pᷳ��u5*�5 T�ݾM��%��C�H167�E�4�g�uJ3��մ@��8�K�Ng�5
V���L�bV�3zgj��I5�Ϻ�$l�4�#6��#��#��oK�4��E���'(���6���޴���~~{���C�6���ɃL5�m�5��^4
H����V���&�2������3�l������(���]6PA�����Т���Ν��0��5��5��4��޶n0�� �2�Wt��6'�é7��h�4������
�
����6� 6��޶^�(�$�o5�3���6&1�56�6`֟�p:!6�h�6(����ൔ|��P����g5`�4:ڶeH��~@�6���p�׵�����56�6��&6�zd��R�5���4;�ǵ�d7�t��J�2�NSn6��Z6��i��T�����5Q|�67K�5(���#�k�I6
��6�6z�6�+�5��-�]��6�����:6�4H�u�l��t�)�hh�f������5��52/�5\�6m�6^� ��B���6 {�4��p����kL6��R6*}u��A�4�h�*86�ZM�g�W5O�L6j#j6?t��8���65�]�^6`���.��pa�4�x�� mT3�K6t�5����@6íѶ�H�6&�#�����!�6T��6�b� �Ҵ�v6J��N|�����+/����5�@���76(6�6��Ķ`�!��5p�%��8|5���0}�5U[�5H�5��6��N�7��6�=��,A���6p8N6\.�6[u6BN60m��@�3�.�5IN�6���68Bȵ�ڪ5�,������`�6�_͵��96�	�6�7�^ε�g�LW�� �^3�n�5��?�>N6��W6��6���3�\�6+��6�ɶ����m������6 �N�1���RoE7��,�jt���ܱ�J��5\	�5�9J���]�件5 �����5(�Z6\�$7��;��'6�?,6��i6S�@��側��*�-�%D��p6p����s�6���~�	�M�50�l���q��b6��4D9c5��5��3��L�x������5E�5m�����˵�貶�5@��3 vZ�Bu5VD׵.��5V3��l��ސ"�W�4vz�2a���C4�	&5�}��;�6F<���Fʵ�b�5��6����<E6:�5j�5�Ac6�B��j�n5@![3ʠ(6kF:�`C�3�`��ڟ����'�S��g��I���$D����4|�36L�)�;ǚ6d n��ic��'�5���8#�6fW��=E���C��	ܴU��5�h6�!4��f6�ȴ�ڠ�
�5^�5(�6�0�� N��t�16	5��i��t'� �Z����6���6$��Ҕ�RR������H4��`6U�3H����v�3ԙ����"6e��/3Ѧ���i�Ul;5I�50�Q��ȵ�%,�\�ݵb���w�N6�aU5��6,}�5 �˴��	��N����5����`h��;�$޵��C��Љ�\�6�.�3��۵�?��~f6��5bϙ58�O�k��36.��h��76��ܜ�4�&�4��ĵ��wi�o��ǟ�5h�65��P�>K$����q�5�y�`�(����)�6�E�2x��%�:���v�55�$��X���G6P5g��8�ޤ��:�6���:5��c���u��<n���=�,A�4�[��DZ���͵�
;�@L��N�5z<3����!p�5�-�`I� !�4@yP�R��x�ܲ�ߵR�6��6l��54- 6���5���`ˌ4�U��hJ6�M��� J6e������/04�%�p�6�R<5(�ֵ��p��mP6`k�����?~�5�c5}.�6�Av4�_�2����S'6t���<6�����68@25���5�J��$��6�Ӄ�v!��`;,�f���0�66X�n��׉��E�5�G5{J"��EU4�P���X����x�4q�$�Ƭ5��4�!5����$�(YS���C�lGӴ��:���05�;Q�X���4܄#��㍵x7�5ZW����^�!6y�5Oc5���4�\6Z�ȵ 5�>`>�{p5�k�4�Q"5�m�5'<�<�5�/�M���X�����50T84(ɵ��ϵ�[�(8�40��4���4�r��]����3��4�h����3�6�f�	�S;����5��5֕�v�g�8�24tд�K�5��5t��5��A5���x����5n��4.m�6�?��k55��[42�X���V�������\6�%��3VW6X#W��9�o�<b6f�M�T��Y�5 ���I\6`b�4 nN���
5'��6�W��d&����q5n��Y�5�$�p�H���6�h�6�-����7�X4xY5[�6��������Ǥ5�d�4�7,6�(�4�e5[�s5﬏�JJ!7x���T5��60�۵�D�5��6�d�6@B5��95�K64�� �Њ��Q�6J����'N5ӯ���`6�ύ4��N�:m:5��6*d%5���8F���1�6��5���WL�5b��6
I���|�5d���{ZN6�4���36�� 7��%5M�ڵ����ϯ�rJ��0xh4��u����5 �ٳ�a���=6�^���'6'-6������4�4��4�AH4��6�B�5�z�5=�F6�56�����>5�}��):���ps�����ٶ��H����5\���h�6���5|K���6-L�𗌶��i6��1� �x�Äh6V�i5V�6�*F����������6xJ*4E�m�N�6�/۶���5�CL���(+��P�ܵd(޴~b�5�'���6�����^� |�5�u�5f6���4ғS����6����������6��)�c�6 c���5���36Zc$66�嶊>�5��5��;6[�k��(5r�=��p�6]@6l��t+ݵ��J�n���}�5��ε�T�$��6�z5t�~�~���yo�@�5��[6��.���N8_���!����������>6�-����Z6�X�8�6&�ŵE�ڵ�.�5���6_��(6P��6
p6�6�"�����r�N���jJ�3ڵ����6\�T�o��z�j�b��4�K�5^9��h�5L[D5��_5��N��R�6�$�x���N�6ab���5�L��Of϶?5$�0�&������������Y�6��6v7x�6��c��g6��P����4��T4ӝ�5�^u6(�@��&�e$p6o7��� s�5��6�6����W0��l67P��_e6-�׶�����+���Y���6�V�^
�5<��6�%�5�����7�ė��¡�&z7ō5��5��58�*�ۄ�6 `"���6�>�����5/��E�&5���5������2�$=��%W�6�!�<�6�ݵ�M;�d�z6@A����H3)f6�3�i�1� Q}5������=ҕ����5���5n��P��R����_���g��Q�4��!㝶po޲�
B6�I�6U���]����5�	6˯�4K�����u5��5)� �
a��� 6��C�@6~�%�^�6��45!��\�6 ��ܝ�4�y�5~�a6����S�����_����6n<�|݋��u�6V�����.��L6p�j�ӵK@	��	����5
!�6͍ᵾB7������66��x6
~m�(P{44HH�jF6r?�6�7׶��5��7p�촉��4%ԶWB��T �&���j��|1�*���i`��� 6�K�6���`To6 �����554G)5�84 ��1�j�]��5*�,6�Z��ZM6&DG6��,6���5��n�gR$5�x 5�߶�B��4���A�����Xδ��B3�7�g��	m}5��6B���(�?6r�i���?5[�,��u6�i˳�C��x���L�D46����(����.��|7�5^�h�Rh5�$6�g�6�#6>k���$��:��K6)NA6��7��
68���j6�^1��̿43!>7H�7"�d�T�6��6(���q��6�ٵt��[�B�K�>6�5���6��0�4�W���)��5ҵ�o����,��:�#6=P=��Ց�R%�L�5�ݔ5H^�L�A5|�P6��p�6!Ӷ����d�:�����B ��"!4Eϧ4�
�5�N�5�S���w58Y5O�5�h�5x�����5�0�5xƿ5�o��Ե�j|��F�	$6��84�5j{5�Z�\��4�Ǘ5lt�4'W6�!�Z˵�?�4��2^�a5h�5�`_6`�6	6�j��7��6S�E6B<Ե"<^6e������86�'���c5��5�v6�T�� c525�v�IŬ5�F6�ě�4h���L��`�6�¶�_b6��m�܆o��=5�6����$�+5�S���x�*{6`4$��5Ԯ絰4�V5���6pY*�2E�5������5�\�����YM��뀴���5O$�4��+6�Sa�锄�J�6�a6�(��eO6Xǒ2�%G5�ڝ5��t5S�5���5��_5h�ϴ`z
6���4�_5@&�3�a�;�5ￗ�@#��Hr�5�1���O��^�5S��6PW��������5��5�v)��#ʵr6��6���ϟ�5`Z�4��9�p��3	`6'An�֓R���Դ�?�4���5�6�5��5�4m�l`q�𱑵Z 6���4�H�3Cng5�-��a6�5�|^6�0N��O����5rFR6��w��R�5��B���6Ҽ͵��5��c3��U��2\5�e�5���3��76�/�4�yf5��5"�m���+5JR5 �����#���56��5"O�5n#5J�U�M��4g�6@y��z�*�`:�n��\�v5��`50�5?�3�6>Q6��
�4���5���W��4�UE�+�ʵ�ѧ5f}�5�]5��B�����6ynI6��РW�xs��H9W57�53L͵=T�5lf5w�5}�5���4����Y��ɵD6&�4�q��x�4c��5ݺ���R6��.��M�R��4�1c6�4�ͷ5D�5�V54�����R޴�'�5>�E���(5���2��p��Y�6 �5)�040���·4}ge�� ٵ���5 �&4�w\�t��5������:��Z5s(K64��5<3{5U�6��
7��յ$Z�5W77r�6�&�5,�26D��5�_3��E��H���M7|�>�<Y�5��6j�F6`&�������6� �6%ȶ��W������+6�X��0�V5��,�,��6濅6]E�%mQ��7m���Ķ��e6ЎX���6
��e�W�:���S��G��f�<6�J_�x
ɶ�ɴؽ߶��`6��6�<�6�Uʵ3=�W�6�������E�5�ם6WPG�v�S���f/k7?�X6髼��]�5=�^�{���V5����D��5 �4S찶��7������l���5�~7F>k�^z�^x\6:86���!�6r�/7�B�6w���¤�JB�6��5xUV6�)��4�6�m,6�ǉ��O�v!�����74�G6�s���e�n�m5h���O��O��6\	�6˱6p���|�6�
��!�u�S7=Ԕ6�%6S'���Z7P��(�76�7[cѶ]��.��5�&��閵��W4�߇�|[���77��G��?�6��61���d�`6Y�&7�N�6�Ϥ���n���H�E7�|��vA6�_f7Mw˶.��@K-�d�5L.6_ C���׵������	ضq8�����5�g#6�3�5j�6V
���1�5�&\�T|6mI6	k7�~��ܦ5���6�4�"����6�E�j�xZ���V75��_6�A�4�1����/}46 Ʋ�T´�� ��>�5a%6�8�Ⱦ)�4s��G�����^���Z�}�
�4��	o6����+�b��6X9���� 5P��4��Ƕ�N�6�����%7.&�5Vj6�-!�ɚ��U�6H�857��5t/���f�`��d�6 �ڶ ���堡����r:66��pSq�Jp�6>�h7��޶��5R�6y����6�.S54�r6��
6��:a׵񒶘$6���5~mM�F�B7=�6ĜI6[=6��6ᗶ��7� �W[�52��$5��6\.�B@�4�U�5�,6��563�5���L�	6�g4v
��GA6��4Ȳ���d�V�ĵ�ܴ��ȵZ�6�W������B6�B���/�f��4���j�J�sȰ5ݳ���5T�5Hn�3��5>�6��V�H�G40�x�:>Ŵ���5��5D�Q�mv5�8�4��5p�u4 �F�)���c�4�T���ҵ̿E6��R�:6����FS4�``5��6'��]ǵ���5]^���ӵ���5��5ND��y6L����4���[K4�:j�%>����c5L���}5l=6�5�ȳ5f��5�d�i�4���oy	5����t~w5P�5n6P5l84�0͵\.5�-�4��4je5�5tu��rZ5�p����5�0�4+'�5<Y�4�e���3���ڍ��NG�5#�ų��5$ό42bĴ(�O��26���48Wô@�4 O�3p&�%ۨ�
t�5]��4�A�44ҏ5!&�.�(���B5��3�io�5oi�|�q=��#ٴ0���J5V�5�IW4������\5��75�ǵ4�aM�*i�5k�G6�^�4��x5k-�5��س��6��85��v5�å5~����5�����CN��a�~��L�4�.�4DR�4kw����5�I�4�L�565�Ⱦ5��6��ӵ���3B4�6��4Z�:5����5,�5Ɣ�F��4���Gq5�6���.j�5���
l��:@�5��������Z��5|��SR�5�}е���4J�5ȅ������Bz5��4�*6>�5Z�5G_�5[�ҵ��b�5�,δ\�
6 �۵H;�43�6��5�
6VDp5  6�qM�ztʹ�#6&a�5%1���OA6X~U6A��b����9�4,��5�f4�1_�0�O5�=�4A2�5�s4�������5�VU5D���IQ�5S��5\��5\�ӵ��5<(�5�]�5�9��<�˵۠���s5��
4�Fo4�
O6ɖ����5%�5:o!�MYN5���5_6� 7�6J���"ȡ6G:\�T��5��.�H�O���6�Z�P�6N�6����X��
�^�5�	�6����,N	�H�5�7�?��������77�q��4��5�x6�97��д-����5 V6N��5��S���
.
��6�ǵH>�����2��6-�'���S��J���T_5�����*;6έ��� 7F%�r(�5��q����L}��0�4]�n6�����7����mi�5�9L6�'��ܬ!5��5�N�6��ݵ�(#��Ѣ5���6 m�A��}��6���6)�ֶ�'�H>V��*�56陗6T���?6�۶$��5������C6��������MR�w��5H3j����5&c6��u6��6vfe�ò��Ro6o�)�VR�6�X*5���6$�5.�%7\��t�5ǹZ6�����[�6Vc�5<�6�IR6�:6H࿶���5�j�6��д+�5iĵXyǵA�W6\��5T4��`7c��6�%ѵB�ٵ��4>�������[��� 5�63ɶgf�5�� ��W�6��d6H9�6��6�@�*6 �Q� 9
4����Ԃ�*�L/�5ɼ26b�6@�h�U]L�4��5�aF5�/�5�(��|��6�F6�ț4��5����f^�Pյ��z�F(���l��PK5�j~5��60��4�����F7���Z�5�Ӷ@_O�u�3��[�5v�������5��3 ��?�6n�j6PG05PѸ�vi�6��6�1;4�v6N�6�H�5xq����6��Z5l_��ų�6J �J��0CA���䪡�<P��6>C�5�R6 50�6�������60�t6\�6�����}ڵ8����I6���5�-�4J�6|B�5��r��<6(�4����,�4�FB�d�5J��5����<B�h�6�R� Z"5 @���Ee5s�y6����a�-hW6W�6�t��C4�bH���U��6���E�l�6�/5��B6��۵�C6��:���6kIP6S̻���5 6 ���535�"���f�5:�5�5�Op�5�"�`_�3u�)����ʝ5ArJ6ųG�� Y6���4s�ֶ�9�6�	q6���6&��6��7+K�6.��(���&d�I�L�~/t5F�>��j0���p6�#c�Nb�ꬽ5�� 5�ڸ5�C�6�����'7Q M�
�
������e䵑�����\���7��^�g��60~��TNh6�遵
B7PD�,`��.7�/�6�\5
��6�z�$����g6?��6�Wд�Ɗ��`�6e]��m5�ķp�45�Q@5\Ma6>N�6|�k�~I6TZ���|R�6XV�\l�5r��>�4�J�4��4JVǵڛ6;�5�D��f�4�F(�.Vk��?
6�E6��q6��z6��5��%�G���Z�I�6Dg6�6Hs�ܗ�5+�V�:w���on�0��J��6�U�����֔�6���5��8��l��&�7,T�6�
�]i7`�14�~ 7�������С6z_���4��6]���̯��0�	7���6.�5�U"5�Z��ƞ����-6k6���40Ŵ&v�6�6��3�]�6��5 ��3 i{��Xȶ�|�5>�6�����:6�38�g5�6[��6�޹5�+�8 ����5ѝǶX6-�ߵ�@��h7:�&�g��R���'7Y�6f�%6k��6��J�l��6����Pw6�T6��ǵ����R�6V��bE85�L�6ݰ���4�v���G�5�0�6�7˄˶�D6C�G5:����)�6�=�B��6U��6��6,6����;o�\�U�z7᭷6��\,�,��6 ��T��6���5�j�EB6dN�6�Ǖ�(��X�j�=��$�q�`6״���6���pM�57�х��}�5* P�N�X6�=ﶂ5�6mM&��^��dp�`�&��DƶhC5x�5j����w��ک��C�6 �n�����X�5�\���GP���:6���5�5y��d?��B�6+����+߳rs7��4�7i0˶���"7�t�4��E6mc���{6�d�6ο���6nnc�l��jŚ6C?��`&B��N2����%�5GV7F67BS9��,7�\�=6��+6��3>Ӷ��6`Z:�7X>�$&�6w�5�����$�^�6����u!7� �I�l�d��6-�ම Ƶ �64 ö�G� l55�+�6�/�"�����	�r�.7�#V�}��&�q�6 ��H��5��c�
6���5: �����6�}�g��6�8���o6�A6 &7X���?��5�H��z69�7{ж%O[69n��,˴�
6(����i��w7��5�ي6z�5�S�5$3�Dl�&�G���4&�ǵ�n5萁6?V�5HnZ�j	�@`����5 lQ0�/���4�N6��W��c62?,���?6�V���$5Љٴh�����@+u����5.][6�M0�C�ǵ,�6_r��8����$7 �B��&���U�Rø�"�P�I���b�6�1�6r2w���6�e����[�{6DB�����5K���`�4(nR��=��EE�.�5	 �6�õ
F66�V'��,����6Ow�0�����j��u6@��5h����>J6��?��j!���)�'�R6}36̒7����L;��6����N��5Du6
vj���ǶLh�5HJ�6�LF7���5�l�6䵹5��J����PZ)��5*�C��5��5�7	4Qw=��]}��wL�V)46�S�6%C�D�:����jDG�f�Ƕ<qS� >�6t�,� V�3�rD5�u@�R�\63$�n�?�ր@6�7�@���'6V!7/��
�`6N���M��dh�P�C5��-6D�����j6ܘ�6�
6��g�C}�6��ܴ��4ޫ�6Tk�5�{���A�b�6�ضۆ����A6|P� �.6 ��3r�N� kX�,��1j5dm	��>��q���8���ȵh�ش��6z��5��/�	�E65���P0�5���5\{�5��5J�O�^��5^(,6��ĵ�eԵ��8�Z��0�i�x�b�6*6ꛀ6<í6�No���x6ɶ���-���o�5���4<fL�Z�m�p��6d��]5J��P��hM���*L5�U6`ɳ�˘5v������D¶d���̇� "+���4�`7�!ඃ�16����ׂ�C��K@�6����6f��X�ٴG�6�S
7��j���
5���l
��t,\�D�~6��t4��9�| ���6g�����>�oT[��Hk5��-6wSX5��T6Xկ�Tp�l��5&�F6�d5 �c������ �5a5�6�U�5�ި4�Q��G��5R��H��5�t�4$[��jO�,�綐�6���4�d��Ȧ�3�(ʶ���5��
4�2�5`�5�>6@������9?]��U�5��>6aEG6U������5�_6�4k���~�56��͵a��
�6i���7�6�N5�ȵ�r���5��z�Zk�5855�`嵴HY����@�״���58�S����5 \q4!#��������5!�.61���⁵R��6	p��`��6 Um�����X5����`�R�������� 7�<$4��!�^�I���>)�6����25��^A��6�����*� �����ܶ��̵D���ml��x����7
�w�P54�64��5iw�� �3�� 76!�h��w6'$е���6j�6��6M�����0�b݌6��}58l~��4��86IX��y8a6N�õt�5*�6�l�ܽm5?�F�  6���5�I�4�֬3��$��n`6 ��4��8���36~�h�0�ϵ<��5��4�b`���p�� ��5���58��5�ȳ�g�g����6|������(3$�,6�5~�E�;]6E���m�T�H��^�V6�iG��f)5�WI6D0��nU��B��H�ȴ6u�5v%�5Y-�Ho�2 ޵��f6��5�ux543�6��6;�6�B6b�F6�o6���%�����5�ג�N��6��0�y�4��6��o�qVU6���6f�r���|53^ĵ��F6lV6V�l�Ő��=#��>�)6�;�5�6󵆶�g�efW6%�?6��6�O����ʴ��#��6ͮ<6IV�4�<6�2l�Kͪ6���5�q�6�5h5�7���� ���X�5�����5svR5nI>6��6oʅ��]4�W�4��hn6���5�����9���7D5j<�4�H85pJQ���v�z��6�_��F�4K皶���OF6��5�,�5n�ٵ&\����ʵ��6H����]5ӹ6�[�6�p[��6��J6�`ζdG�5�a���L6�W	��F�5�6�5�6eZ⵷O�5�'Q��P����Dx/��N6|/�5���6>I)�&K���T����<�k6.����Z"��z2��}�4�!4z ��������6�])68�F� )0�`fp3'��^F7�[�%6��$6�[�4
$6��5�p�5r��4��ߵb��~8"�o��6��6��1K�d6�k6D�_�q]y6���������ME��=��S�4��6[�:��pn6�+5p���{�����-6��#��5ӓ�6�փ��VD��騵&혵a8�S5�,*�Y��\1 6`�G�p߱���f6�E6�r\6ps��!����Ե�⓵@k<5۞�P�V�I�%�A��R35R!�6b�W6���4��6t��@9%�UI�_�g��玵�PF6��k5�w�5H"e��f��Ļ�4������64���3��06@���@V5�[-6�/k6���5-z��l6�#�6�F�[�5��v6���G "6L����a������50c6L�5����L5���4�g3��Ef4�o���x��@�����綇oP5(�5��}�5⚑�譵*ڼ57��|�H6�5���$�Y�&�۵L��4� 4�b�жփ���(�f�xE���r5  �/@�P�%��6�5@��a�4v�6F��6�ڸ�To��;�@r�3���!̉6�5<$.��Df��,k�+5ge?6 /o����2�,�\6��ڵl;����PS~��[�6"�95:�\6¸B��NT�:_�6�O�6q�6�6�J�5����d1)6?/���f|��36�P%6�5kl5P�3�L�]6��o�N��5��8��8�5�z6�Eس��6����7U����6ĉ6(�5��?5Ys6���M4H���5�W��t�3���5��5�b&6����g�5 �94G�64b�5�׀5>�^�[-͵�Ł�țp�P/g6X�����6֍z6xQ86�Q𵔾�����B�55��6����DF6������5�:b6p�#���16Fr6ܐ�ǽ���6P�4��5+6�F6��6+��5�>��
��5�6F
���͵t��5D<*5���5���4ՠ5 �Q6H��5.�J���"6��o��=㴀H�P\�	� 6�n�5$�5�)I�pN��0<�5�,�5k$�5��5D���K`6�����/6a6��d��0�6F`L6�ﴵ+�4�����'��A5֫�6�%�59$�O5���[�4�	�4��ô��5�킶q��5n�{6���յ�7�EF��];��?6M�5`�5�'����ݵ�����x6P�36�T�P����3���3��b��娵;�
���f���p5���dD��~'V5C��K[�6a9��n36$\�5 O�5�㵰�W4K06��:6ة�x���������N���4Z��5<66��5Z,6��6�
�5�O�39��0�2��5��N5�~�5�"J6"�B5�5�5�5Nl 6��B4l�5&��6)0��HC��
�怶�C�6�Y�+{��Zb68����{��h�u�^�B6�Pk6�V65!��8�����5��5|ʪ��'`6��"6��"6����6_��4��:6�5�*��[��Q�6�2�6*y���w�5kb�pX����5�|-��V_5}S�6Å����̶�M��@:K5W-/�I�J��{ӵ6��0n6gn6"���p�6{K�6�a��"[6Z`�6<Ė5`>���\ǲlъ����!3�6�9C5Ϊǵ�Fi6~�5�"_��̄4��7�ĶR�6x�x��=�����a�	�KP�6^�(��6n5��� �����5T���,��5�X���<f6 02,��5��6�2�k�R�g�v6�n�4����Y7T���s�'�6�ئ5�u���16��5�;n���5K7��6�񃶠�-6�Ӷ}c6fO��k�϶���3x2�5 @55m�A�T$.6�16hE�5�I6��16��̶�!�5 �	2�o&����ƀ���R5��$�7̚�!; �%��5���vKʵszU6��ֵ��Y6(1�5��������@ 6 �ɶm��F�4J޵�nx5�@�vh6S���0\�6�;ɵ�@��!��P�5l�.�56��\44�6TF�6���64
쵀p�3 ��n���:�6� 촜(b��M6�+�5��X6R̎���W�;�n�}�6�1�5�d�;�[5$s�5����Z|����?�� �5�>�/��6�&��x�4<w�5i,6 U�3�q�6RU96X��r)���j�A��0�6�$͵n'�5rQ�6a�`5�5���`6%��6 {�5A������6�~��Bl(6�d63-6��Z���5�y�4��6E��6��A6 �J6q�7�7+� |91_��5�6�6� � �ƶȒ4���5���i5
6���6#�*��r6�k6R�6��ѵ(�B��(�50o�5��5��6�Ҭ�L�����5Hl�`贬��6�E�4�a6�6$�{��{Z�t�7��6�m�5�~��Y2�6�/6~\5�`6\��6E6$6�6垙�@Բ���5�,�6�6e�$6��ʴD�{��k��X�44��4l6`�}�6rZ���ݵ����5�l,6��#6Y�M����me��S�*IZ��{�3H偵M�Y� �P��ę�R��6�>5U�6r����M5,�L� s��َ5i�e�!�F�"WZ6 @L��r�5��4��6���5�}6��R�!C����U�R=���3Nۑ���P����4�.�<�Q�xρ�@�6}�54�-5���4t� .O��@w6����Y6�s���S��(�5��f5 }�2$#26�-W6�vF��G�4w�76v�'�ho�������5��@~5� _���6&�5Hg��b2���յt��4��M6�6�66n�T�Pg��щ�0z&6@��3>�4*�=��;F6B�5����p6=䵆�6��l�����'t6e��5�y���l�5 �@��3O5L�5d�5s6VC��>�5iL6��5~�5���2r��s����06b���V���4\c6�I���5�>�5��C��洂�������M6Ll!56*���r�5�`<�ծ`��2I�`1H��J�5�㶢+��q:��&秶����>36��Z�36�����[�RH,�z�^�ĮY��si���6O��6�#����6��5ƪ6�75��6�6�6�6�4,�2�Ȇ|3��m5�C���U��W���	�5P6r��6F�6�5��4�u[6�O��x�
46)�Ђ9�O�6�,3����5���no�52����Ϡ6�ܦ��v�65C��m�5�� ��Cߵ�5�3r�$6Dy�������N14�WE����������D����5���5�V|5�1-�~|�����`'���5�s,6h$s�Ne���,5׃5JA5A�5����Z����)��P6��5 {43'Y�#d-���5��c6,��6Se��P�6~����F �����#
�� V4����/�t����F�b���~OM�;|��3�l5�����e���K��0�B�g6�~}��vJ6ߵ�5F���Z6�׳������)�"�?�V�����7���5o�5���>��ƭ�6.B�5��`6E�ö>�6f�Y6�k�5Ҧ�
�5j��5��(��B���_�pB̳��6��4y����]6�i6ֳD�`�洜�6 �Y�����,0��?��6@�(y�5�YL�F՝�D�R5 ��3FD6H�´q7����5��(��.綐E�3�O�6<u7 �.��/�V�5ĐR���c6`)�#��5�Y�5X�ζz��5 �i��^�6p��Г����򵫳e69��6h�����p5T�@�N�#�ٶ����d���[6�+�6�|6���5`�v6�Y�5�V�5Ҵ��L�4wȶ(�S4�F5�06�1��tu5��X��4L*6aX��D�ʴy�����4X�96�
���8d5p_�4�P�6ޥ66����#96d;i���62�ض�N�68�5/���6�?(�3`�5�F������ 7���\,�����5�S��J�6�@P6FZY��y�40�A6�8���=�5n�6f�6l�5l���iȵ�����6�9;6x�s4Y�6y#��Ǳ���5�=)6�xS6$�F��4�w�0�@�6���p &�z"G6�6�&�l�62��
6LVh6���6��7����v!P��ٵ$C4�hd6&�s5�l��L�5�|���V�5P$����;� �.��L6�� �6�|�6�14�\�5��5l��5@L6\)Q��߾�*z(�h�ڶ���,��bg5�vQ��O�5���5�j�5 ʮ6�!ζ4]��,7��5(�5�Kd�>��\[p6Ϸ���6=A 6<+���&ʵ��6Ц��p#@�be����]6�q5&h�h�T���x5j�!6�;�H�z6X�� �*6 4��:��
Ƶ;�6�7��X$�Xi5&w&6�x����Y6j�V6�������е_�7���5x��b=����6�)���2$�t�6��m5��6��Z���۴ ����nt����6��6�=�6��6$�4��6�Φ6������r6�؜�Q�3?�6IS�0�H�I��60�E5ď�6!�`�X��6�?�68���S�pH����6�9���WP�pS�j�f6L8�6/g��?<��U:6��$5J|�� e����70cq��j�62꽶�5�2�@�5�45���˗6��L7�{�6FRx����6i�F�E7�	�p1���6���5뱇�$��	�6�:k�8�7���4���Pd4�5,����ֵ;��6{��F]Ķ�%�5F��6�Ԯ6��5�'6l�l6�N��wCݶ^Z��d�X�#t(6/�6Nh�5��04V�5,�6@���/��H6����ΰ#7����|6��6 K7T��R��̈���4���!�6�D�4�!���6H�|6��6��y`��Yt6d�6$�%5R�I����6Z�����6���4�/�-I6�϶=\7R����ٶ �(4���ֱ�*�öL��e7:+�6F�������k��-05j
32�3���qު6�{�������V5��|5If6zm�5v�6F��k�6�O�6Z�� Vp4F���7������7�¾5�� �,��5�7�4V@l6=Z16"��&I�6��f6ö�-84����d�4o
&�ޞ�^��6�]|�RIǶ�k6��/�/�%7��ж��6��3����50�/�l�0���6`�4���5��-��G6�����lq�6�R���M6�X��
����6��6��6B���Y��6*W��f��3��6[c6���64�t6_U��W6̝� �+�t��5h��6��5[m6]7 ��4P�O6N$�¸6|�[5ܓm5�l���m��9�o�����k�๟�`�6��5�5�'�4,�7��Ǘ6�&ʵ(���o��-��6W��5�+�V_7���5�'R7ܯ��jS����57�y��9p�"�@�I�#��~�6x�۴/�6�0�4�s�5��6�<��&�5ԛٵ��x�X�u����5;�B�$� 6�4DK6��=��>���i�6d6�#��uQ�6>�)��$�6 <�6F�P6�64�Ɏ6�����}5��������g6�q����?6\�F27�A6G
��QT�*O��Ӕ����5�D�6P���ڄ��4yn6��6�J�Ls95��6���6��A7̖�6��ж�cc��'�6l��lQ�'R6n�͵���6��k�L�筶�e�6A#7�^6�]�$6y̜6{����ߴ*:O6`s6�H6�\53�ζ��}6>�S�~!�6_��6�I'����e,�H� 6�!����(��l�5,쎶�����5�x<�{��6��l��А61�6�>ڵ��4Z9�5$�n�C0H�����@p����5'v5�~"�����P]��8�L� ���_����)����6$Ú6�x�5p
,4�ii6�඾u��x��5Ђ� �6.06�����w6S0�����6(/�6����ʿ�������^/�����᏶�~����T������6�ո��ĵ�^�6��5z�(6�����`�\�68�S�7�����4�	����z��6���5�u/6x_�5��ֶ,N4��G��4)��۵�8�5�V�6.����Ւ����En�/�7��6������@6%�6=��6��6��9�7%d�>� �n,����[�)F���.5
����W��oX`5�����$�6俐6��c5�����*��G�4�3t6�1���m�6rk����61*�5�����5��v�6�&��=�6�ə�@Ǚ�^��62U6K;���9Ƕ��5�/ٶT��6�(��zF���5<����6Tu۶�n�6c��YS6[<~6/�Z6@�6,6�"���ѵ��*7�綕m6��]�����>޻��
q��qi���6���5PTF�P��6P��58�5F���\�5���4w����Զ�6s��6��5S
�x[q6�f ���t6�iX�,��������) 5�2^6��06�j�5顷5�R^��R6	_�5��6���Vrִ,D�6���6��-����Ԣ�W���7 �Bᆶ09���5�6��75r0��$�5��,������� 4bж��q����4ē��n��h�����6�����4� ζ�F��.�5�~��̊v42���&}h���Դ@��j�v��&n��'$6���H6d�����6(��~G ���u� �w3�Ff��բ6.�6b!��渵p�!�X�?��?6�۱���K6��y�*�5@�ܵ��67R������ �����Z�6��|�⪶J��6���6����4���6���3� �6�BL73|�^��?���5#�5%���S�G������ H
�I�͵�ĭ��55��ڶ��+��)W6F6�Q�6�@p��o�����xqc�D�C���7^ϵ��~��6��P4���6�ȶ6B�50'൰7>�DN�6NQ�3t�6��60r�6��4��5���61�a��f��*S6������2��Võ������6|�+��P�6�ϵ6Ө�5�w)5Q$�5L��4
M���6�K3^!�6���5=[�5K�7�Ƨ�J�b��ɗ���6<�4v�A��%@4�Y���ݶ޵�S�3�96�U94j��5��6�x6�7�.;6l��a,�nS7�P���5چG��7N�`��3�8�G"εB���n@x���6�?�6���5kè6�����w?7��x��ض�6*�	��^=4���� �Dz�5��ǶEL�\����m5�,r�|_)�O��ʽZ�n�5�W��n3���6$�E5�~�6�d���k�6�: 7�����,60���r̀6�޶b�07 @E�dd����4K��6��/�$�5�6�ia��� ��J��Q��(V5
��6H��4���6"��6��D��o	6�]�V�>6p٬5�	z6�o��mc6��޶����
6$��6%<72������6n�ɶ�}@�P��������5T9<�8` ��J!���6�;��~�T5.MS�r��5P��4bT�5$��6�4 i@���5��7�>Ə6��[4KV�����5p�-�PX�6��������6��E���,��jе "!�z ��f�6X�u6�%7� "���嗶'��6ȱ�6�_��A�6��O5����<��4�8�6@�6����6M46�ӶR"�6[�5�}5L�������"E6����(�6�	5�J-��v6��7BA��T���d�Ҵ�)�5:�ն"�5�tI6vm���˽4~��|��'9!6���({C��J�p06���6C���6�U�L)�6��4�q 7XR��g{䵔}��񃵛�{�%�t�O �6|5�6ڳ�%[G6�	��5�5��ɵ�6?T5�W5u�K=�5h�:6���5� ��� #�:$a6t�J6�Ld��5�|6��*6c_5n�j6i�	��浖�Y5��6��г��6衧���5q? 7p譶�(���G�4������Ь�4�_7\�5P�4�� C6Q���G��6<�@6��AY��"5F��6��5��R��Q��t������q�5>6�¶=�$���ĵ��ص+�&6�ֶPtu���d6t�A6�55�d�ta5����3�z6�޵��B޵�C�5�^5)��5�˗���52¯5���6玷����4�Nq6�H�x���֑(6@�)��~�6X�j�Lw6�!61�5&��P��4���5l'��@�6�����5U��neV�h�s5ҳ ���zε���6z�")ض�}�6�ꗶ�l�5ߢz6F2�5��@�� 7��3D&P7�7A5���6`�6��6d�m6/�����J6�r*6L&&��N
7�~7@�Z6�>�6?�]7�}���Dt66�6]����G���Ö����6<��6�5�Ӧ�,u��p)�6pڵ��5��6 ���8�3�j-6���6�
�6�m���S��3U�N��5�-N5y��6���@7��o��K�5ʕ�N�W��6@_$6z�C5|��^AH�!�Q522�5����TC6@�3�ӳ��B�V6�5�΀5�/4��-�ͺ%�2�6
%���Y�Ȭ\4B�	6�5�p6�ф�S����5$�?6�7e�P*g���R�jT6�a5Fr��@�15@�������q��?�vE� �V3�\�5��4p�/�H6̄%6�5�K�!��6Ӏ_6«$��p6`�ɳ0w���K�����b!�l�5_��5aP���WF��N�p�5!�6��kW��6>���w�4 �b3 еý*6﫬5�K62�:����S3�5_�4��y�$�6ܳZ5�ꓵB{���N3
6>C6���5 |�3��A�PH6�õ��5l�f5��)6�7*502�3p��� ٲ3��6��,6H���0�4�t`���5���L� �´�L�4(ED6 ��3���4H��� ��1�e6x�5�f��~l7��7�4=�6,�5���5�'�6(\�4x�g�xW�5�M�3x�����6�18�X_j���4�06��3��6<Q6(�34�6���5�4��T5���5||=6-�4���4p�5�N5��4�:�(X�4�㧵"rU5N���T4B��3jcH6�Ѧ5�A�����M�5���5���$7�5���5�E��摶C��Ow�5SoS6��S5(r�5�^�5�m6(x0���5�y+� ��2�ֵ�5`a���	���{4�Fݴ�G5��؇���j5�x6�8�5��� c�5��50���#���_L5\���A�4K!6�(36�0m�f���c4��6LV�5p����52�m6��5��~5��]� '3��n�¡ӵ �S6HH��ԯ@5x�6���4��(5N�5йR5�:�54�5@%o47��)�g6�}4\�[6&��5��-6�*5�}�����5e����4�b��,]��<�5���������OǴ��G5��4�(Y����5|�4pe]5��8��{�0���µ�G� ��y����5TV:�C��5�"e�tl¶M�"6Bϋ��sĵ(�b6���6$�;�\��8	�6r�$�pG۶D2�6=Ű�q6 �j5�̶<b��F�6XT�A�Ѷ[�Ҷ�86J�F����5�m���fi6���6��k���v5�,��~��>!7
@�5�e+5	�k6�8q���ƴ��6��J�R��6*�6�T��0��4 $/�Jr�t��5�FG6���� l�@�޴vfյڈ�66"�|��6V�ȶJ16e}7�Z� )���D6�/{�y���c�$Z����ضn�$6R�ŵ��ŵT�$7��0��(�6��x6!�%�9���a�P���z3�`�y4o�8��ѵ`4V�6�6D=���5Y?1���*���S5��k6��6_�5|p7�W�6ѷ�l�5DG4ѯ7d6��µ�W�4$���M76�.T��]6V�ݵ�Y 6 U�3g6jN��F�6^�(�D�c6,w�6��z3�G��.��5��(��(��8i�5J��5�n�6J98��c'��Y4j�g6��X5s�4��.6­��P+���36��969��6�@��2�󉫶��^6
x���O�76�6�V6,.�6��f;!6J�6�b���_i7!궕3�ɵ4ٵ��7�g{�A�F6
g�6�b4%H6^�7l�S5����&�5��4�`�5&U!�y���$��6���RO�6��4�'{���5I����6�z(6�LC�F�Ե�\z�(%���S:6��3�66y9�(��5�Bw6���� �W2��;�>�G���4�v76M6��'6��6N�]60T�6�O�5�KY6F��6PrX5�w7�Ri6�7�`>6X�4X����(̵�)�6W�37g	c6��H6<!T6HT��Ж�a�G6"2��A�6�1U6���6�y�6�X%�&ƅ5L�h?���_�62�h��o�6&#�L�=�y_<6h;T5���6�y���W6��V��մ:X���-�6�~6j:���6��7�<6�W&7���6�vm�:�^�$��`�;6���5��V5��5��5ܞ6(s,������l_56h�5���)��5�ĵG�5õ�J6��5�5�?*6��6�)�5L�66^@�g�v6մ�6zD�5 "Ҷy���b6B"6 ��*�6�-6m6�e�6��6��+� �6V&�6n�5W<���R��N�zg�6�:��k�4ұL�n؋6���6
M��X0�5v�6�$1��^$�}��5s��6�~6-P��F���6*Qҵ��6���4�ި64��4��6��D6'iöB�P��^U�p:�4`��4`r���bǶ,�5lI*6�*6s���f�4��6���x0�8uL��ꋵ�$�5�gL��u'6��5��!���[5�e�`!����Q�`�n���4RBy�"����O6T�)�ԸE�����w����n5N��5�7u�n9�5¥��o��6X�鶎�!��ֶ]赮ص�2 ���.� �2��6����s8����+�L�3��t6�׈5�2U�L���6��R�tU�5	K`63���h���i^5��K�6@o�����50�k�b۫�L�3"h���n3� �'�"y��6�o=6���4���PS
�#��6���6\�@�<2]6x�ʵbk6`�a4���OQ6�6��/��V����ʡ6yU�j'Q5Nj����5�6x�C6N6ɵD�?6n�o6�e��y�6\#���x��|Շ6T,��v˥66�<�초��5�6�V�6@�2��p(6tO6ߍ7�@�6|�S����5w��4H�[�0Oi6��U6��Q���e��΂4B���P'��;��<_�5�a��i�����֑f6��˵p˩6̱���𠶠�+�iM6�)'�r�55TW���r�¼^4D�K5J�=�r���n����5��45�a�66tL��u.5�(j��z���4�5FEb6�e�6�Z��{��M'�6~6n��4>d�AB1�^Q�,�����~_��ѵ[򎶵g���]�.,/5�M�5P�,��쥶��\5X߳5���4�� 6\1�5�O�~$�4W����oµ`TT6�i��`�5�@E6�sN�{�p��f�6de�6 +?��o��NU6�-��Cyy6Gߵ:��6`�2��~�{:p6�
94��.5���5D�"6�a��w�����5��ٵ�k�5'$�5|FH��5�6��lGS5D<n6�$�5~��64QܵH۳�����L埵���5�0�5�Գk�76%��5����36���ںҵ�Q �焔4)-!�4�S5�ѷ5@q��r͵��d6���X��5x�4�g6۩@�̈́6X�/5�����jF6��6bG����5���5��H�
�!6ƛ���)6~�6�6�ስ�>4˙��m���^債�+A6�?�5K6A�46��X���>��86��5^�\6��5�l��J��:#f5�S��?�?5<
���̜5m?:6�ar�����5�d6|炵`?6��	�<rH��"�5������Ĳ���6�����5��24[V{5q(8�C�6�)|�H,�3�3,↶"{5.�46�u��7�4z.���(�}%6�DR�h�)6�.�6�<6��񵀆m4L��^#�4��-�5an$�w����e��V6�,5�zC�h�'5*�4�߾��a6j��ؓ}��Q6��x4��{�?O�5�r�r� 6D�'4�I��s�y���4ގ��V��56��4 �7�7���1M6���55rF���	�J�Ƶ�j5�)6��5ȠٴJ?6MYs�Q#6�k����6�Q�([:�X+7JO�OfF6�6b:�I�6�68c�5T%5�ס�+v�3��Ѡ��6��<&�50��5�Y&6,@Z4��6nt��M�5h�Q5�h(6;͌5��5?�b6<���" 7Tk'6��x�ކ�5|�|�>�
�����ttгw5�q5 �����5�z��T+�o��������&�Nj�~6^�D6��a���6垳���6�&)6�ׅ�&i4�T7�a�HsN5]�6�6*�5��ص ��4�P6���6B��IǢ6#�5���5�zq5֧6]{�5��5L�Ŷ5�|6��5�r���	3�� �6��۵�%5T���4x�5幺5��ʵf|6F���@j�3�e��1P6������	u05���6@�5�P�5�T��(�6�走( ��n�53�6 �@���5�[4�Xӵ���5���4��5��4ط��T��4�0����5�� 6 �5�m'�,�x��c6 �6T+�5��Ѳ@y浑�����#5X��5!���v�5�϶��;�i���W#5�h�<4��s���s�u0N5�b��H2��T��� �^��6h�j��(W���7���Q�������H6tH[4h\Y�6�5Ұ�G�{�ĥ`5h�5�og��&$6 '$� �Z6�Y�6�5Z��6�p�5�bڵ���4�s|6>O�5lSl6<��5�<6l<�6M)46P�49�ɶh�J6�`�5h�����p�Ԯ?����E5X(W��#86T�.5Ht�5oV����6��6���6Ր��t˵���5��	7*�y6�!�5��6�݀4@�>���5@!�4��+��6�?8�`0�c�h����nN6)T�6��6�e����6��6*�6�0�5�}4��G��q5�
�0���ȂP�T���ȶ��b6 V�����f��6�r��4�^N�\�6�۠6G�y6#����o��~�64�۶���ܩ6�3������^�5��W6В6�(�6��8�����d�
��6�k�O4$��5z�66 '6�,ȶ?����6�
�5,��6Hs�ZS4����/*j6�4݋[6"�5`�S3��6�v�5��2A6Pq	6�n��'S�Q��x�5��5O^6!I/7x㤵�\�6+W��5<��05"��4�O5��*5ԑ�x��5��7�`%�6�J�6�lr���+74(鶒q���K�3�.׶xS��F��_����8�D��5EµǶ{6�06�u�5i��YCD��i\����C�5jB�������Դ��>��K64Y�4�7�Ҷ���5�^6+�ȵ���3�>V������'��� 6�u:��U{52�D�7FE�k|V�ͽ!6�6b�7����g��"5��&���'7ȳz�e�6u�p6j����o4@[����4���y��7o�N��p}��ꖪ�<��5� �6l4ʝi�`9�4@�����Ѵx�U��¶n�I��6����to6�C�6��"��6�>68�����ö��N���2���{6��6����J�`��4��40�r�rn�6���h7f��I��ސ�^ 6���\�78�6�Y!��T%6ۣc6��������5����""6�߳~�E ��4�6iI6��O�Т!5/�z��M����p��4fg�D�
�&�i�����5��|a,5��;6U���Ͷ�K����w6�ܵ�wR�X/�5�i	3&6��֒67�0�2�)54���5�ܻ���̜+�Yъ6��6џ�x��w��63����J76&�)���t���bPѶxP�5Ȟ�4���6K�6�}�5�OB�5Ҷ��6`�6��|57u�6"�6в�4Ʃ¶�7,�T4/���x@����578B�N^�5�H�����74�N�x6+ʵ�Z���"y�����W�<k�4ü�5WQ70�Y5(�Դ�6=�%6q��d�µ�J�������7�����2�u�¶x�"53)05�7C@��t���5`Ҷ�������ˀ��ϳ�� {6:�T��I���k�n���`�6��?�(]59�ŶIr�6TͶ/��4Ć�Ҹ5���5�i6��5��4��(��Ͷ;P���IN6�򡶍�.�G�5K7Xw15 �e���5а�6\�}6/p�2(�6�O�6Ȕ+�J�5�t$�r��5�z����4X�4�ܙ����_ڵޅ�3�'���*��K�����6)^�hX�6�\T�4�����.�6x��4���� ܒ�R@v6�C^��%���
�v5�6��5���>�56x�9�!�&6��=5��o�ݯU6d�s6l8r�06y�ƶD5���
�g�c6 �k3�В6X�42��4��6l�����յ�#�;�D�p�T� �e���4�!�gy��s{5�or�e��m|(6*p�6 ��5a(���6嶇���2����p}n��a�/��6 �:�=6�ǵt����[������}�7}��63������60� 78.��g4P�-6���3p��4Ԧ�4��6� �1�۝ⵦZ86�&ڴ
��*Ж5�D5>�6ڑ���Te� 66&��5��_�s�5��B���54��pz4{�B�0\a��L�68ӊ��X�������o63�6���4o��3�A6F����R���-�6u��������ib�QP�5��6�w��/Z66�6�k6�2����w�X`Q6�;6>#�5�H5߈p6U��rwH��56,��5���4���5�c5�dH6�U4�e�t�6�K6
nP�4����fJ��o�5藐6�m��'�6�2�5ĊZ�^�Z�?�
}6S�X�ʃg5rW�6|�|�<���*6(�̶�,36@�ɴ d2��Y6��n�Z��62Ӆ6�p�@u}5�{�h}�5�L��W���ζi�K6(���je5h��5(g�5 _W�u6�6.360�q�P�K��8׵�K�6�cA���6��նD풴� %5���*��\��50��6��<��>����-����6�M�5��?�C���	�b�X�}ٌ5�З���D���G6ڪz��c777���:/6Ԥ�N�5������r�g6��6��W��6U��%��6@��䶠�J���6�Z%�v -�dZ�6�_�6|��.!�6^X����:�3���H����_6X@f�?O�5�On5�J|6��µ�@>4,���T\?6���Y�����<�J6������h5G$q6~��"l^��""6b;���Ao�<��Dx�5T*µ���5n�$��襁s�M6�ѡ�f:��6��\69n���Ŷ8�~�n\���$�ce7h����6h�?6[�*6BA��F8��k�v�nѶ@d���1s6d�h�9}��ȵtk�69}6"*���6}7��Dj�*��6�QM6j��{Ć6�8a4P<�48F6��v��5x�5�����q�4ߋ5L��3��6!�r6�\�,��5>��5�g�5��5���5�y�|�Ӷ���) 7�����N���=�5�ϖ6��54�C6̦�)7�<Y*6�6^�d��6�.4 c=6h�3�h����4�c�56^����[5Ų4½� 
5�p��V��5�d5|~f�DJ�p/5�e�5�H����5�2մ�:�5?�6�B 6m�;��6�4���I�6<���y�\6��~�J�����t6-�$�6�p6 ���i	6�т5.�t5_Hf����5��׵(#�4ξ�6Nr�5������1�5D�Z�����ε�k�5�Ma�\n���#���6����d5�%�5�����rm�06X��5T 5 ����S�~ۣ����6�]�����4x/�5v�}6�Z�6�x6��ݶ�j���0��7Ե~;c7�'��0��E���G����5p\N6�)6�-|6%/u��$�4��16�9i6���5P�����46
k54�ܵ�~6��m5X���07��	��{�e�G5�kȵd"b5�l�6��>����5�� 5�>:�n�6��\5X�4�&�5��g��S��7���r�5ߐ�5)ǔ5��N4'�6B��6.Z6m�6�PY����57|�5��6B�B6��N��w�5<1���1�6���5.~�x������4ܯ,7�9�s.6LVS6�v��槊����5G4<O����4��5X�05��C6��6�9ʶ�r��=�T6@�@2��6�~ֳQ�K6��ŵ[緵�ǐ6`�p�0�5�y��O�26<*��8�a5q_56�!���`�4�a�6�
�5���6M%�6�΍5���5c'��Č�����>��6���RT6���UN��:IX5�߬�$�	6⹪6�Q6�U�6����.Ѹ���16�W+��B���6�HL58�N6�͢�Jc�6$���~54Գ5A^76W�5H�A�|�s4�X�z�6�mR5���(zb5
���=w����5�!�4߄r�k��5�n���3�T�4��5�%5ȇ��^r����5,6�ν6�3�ٺ��V��h/(��ړ5���6d�*6���,f��*6B� ��4.6���5����5�p�5rGr�GO<���6�a�6W�L+�qo׵�����|6h?�5�h<5��������5�Ӄ5.�5�p�5���A��5����B� �8�40�2������ɩd5��|4��ӵ\�ݶ�7@��6�Z*5 �a��h
2�+�6�c6����J��6P��5��G�q�E6��G�y��5j>7W�5� �6�{6t����V��_�����5y����c��̇6�ri��6E��W�qC26�����5Ŷ�GM5Hk���Z[T6��6إ�6~+������!|�5,H#6S�D6j����4~���u�4V�Z5�,A�U����z��,�T6 `4���6���0=v5�Ti5;��6��6R�/6f�����s,�}�7x� �;C�6q	�5���5ޅA5G���6��5� 82�����M�6�X6�9��܌�h�ŵ�z 7�7�6O�50~���|�$9������Y����]��5U��6�����ضZ���)�6��Զ����k;���>5�16a�����(5S�)7@��5���5��p6��`��4�l�6n%�6@�ϴZ7�� �6�g5���6d��6�u7���-7��r6���6HT�6�f�5h�T��rε���5DS4��Ŋ62�6�6�P�J��6��6���1�[5��5V�6�Ҵv����64_�4�^��Ȩ'5&^ض���5|y��.�4�y���6�Q��6S�.5j6ֶ���5(��5w�ε��"����E�6�e5�3�6db6�y6�Ab�ԁ15,>׵ �����V6�
����� =�gS@�-�b5n�J5����⮋5��6N#�5�f���ji�>�l6d�5�eD6̂����ϴ�Z�*�6�����95+�����5y¶��h�4jv�5h�.5�m�jc"����6���6��:O5�$�5�|*�w���L6d����m�6ڋ����5Kd/��;5��4��5�6���:5�y2����5�J6��>6bC�����+2�0R1��zܵ�>z���5���R6WB��4����F5����\��\�[@5��537�g�$��A����'4$�����6��w�ڞi�h�g��6E��v?$5 򐶭C�6Dc����e�d5��6Y��5�<嶔K��j-�|��㧵 瑳�ԑ6>�������(�{�96�9���~6Ou=5�*6d��6��p54���*m���y��ޟ���S4��5p44-5��'���6	u�6P=5�m6���5?W6������H�5�ɵ��96�:5��6�pE5�<6,��2R�6��;6Ra6H�6F�@6n�25�Xo��
�m�D6�=�4��5�b��j�5Έ`6p�g�
X�5j~��Ȕ3B^���Ć5����T�Y�C�����5�v�6�Z�5�4�6��5Sԣ58�G5{X76\�z�Id4�&:6#��6 i޴�����EG�ԭ˶��&qA6In6l25U6B~�6 F^6�nm3��b5���a=63L�z�5�q,�0F5P�R�ehg6��	5��6��L�l_6��Z6�6[�P�����µr�6l��N� 6	w���Q��5� ����`� ����#����H&6'L�o8h�D)'�o�5$��YA5���4�t�5� ����5\�N5@�(3�^O5�	�4������6�7�5l;�9���~�h4���4а��g�� ؈����5o��49I	6�p�5�	�5�&4��p�5�R��ہ6{��5-�=�=��5�V�$�#6�j6���Q�=5��9��څ�*� ��a��r��5B6�?,�)�4�����n���h��~w6�M �6�Y�(���ʵNA26�<}5>����%q5S~�fp�5r�K6
u�5���5�6 �L6�ar6��Ķ�Y���gD6@a�+ʏ�({��Cp�5��4�O���r�5��&�D�C6Xf�B�}���`6,��ε��7�6`�C���5��J6��H�>�&6��F��ų����k63�ʵ���4_��6Fѵ1"��PJ�5�n��$�\5\�E6��6U����c�4��4>�3S�5`�62a�5d�96 �S�m��5Ͳ!�TA�50��3���2\���55�<��5B���5ߚ���<6���� �9���r6�kѵfw�#PL�L�wN���4 6�>� &^��ܵ��6�g��_[��2޵w}��9��5*4k5��$3��	6�4��?�5�
h�"�ݵ�����5���5�`��2x�4�9ѵ�*/�rv�6Fs>6��5��ҵ��4��
5�250����3@*�p��4I����c���U���劶� 6F�5`�d3�斵���cB�0Q�6�@�5�����5uq��B�,P
6h) �� 5��5/���W}�����/�6_�"���� �ܴ�I�	�
6B���ސ�LE�6~65�5�0�2pR6E��W\��%�5N��6��5�i�u��:�6��5H�'��s��YL�V=�6��`6b�5��5V]�����\s6@|������b6�~�5�Z�4ٯ3v5]6��5��6��5��h6�(�4�K6Ev��@��5�H�6�q6�26�r6�����'6�<-6��Ե���|a5I�6x!�5��`�5LJ�5JZ�5(�6h�Ѷ$Jk5Ѵ�6DV�":51��6��ִ��76*(�5��6r����'6�:괬����9(62�z5�wF�a7V�2�;6�x���,��6��X�4T:����4��5��K��(�6`�{�~f�5Ea���Zb�5w�L�D��|�6T�����::6��?6�V��L�6c�϶0�6P���È�(6�6+��p��5�&5P�7U�}6��7���R5��|�6Y��6t����l�5�����.��f�6WΕ5 ύ0�r��)�6���˗W6���4	����i�
#7#�@6������6/��Dk�h:}�����t3cu6ZضB<Ķ��Ҷ��$5Hu6���4���5p��S>76�ws��]�6�o6��5w�;6���Ȉ�� �`�P����|'����5�C�5����h�0b쵎��5dV�5[�6������6�]6N�������R��G6�w6Cu@��{��_7�v���6.�Ŷ�� �ڵ[��5RD6PT��0�5:H���O6~56����w�4�^7��55'�I��6�;6B9��x���=�5H��-�6�Z���yY��8���6��Ͷ@�6�XյX5���6��w��h��W�r_.6[	b6b���v�m��5f�6ZX;�=�,�ۙ5��	7��4P�� �7��06!+�6��6�6�1�6w��Z��Q-�5��6��'7�%F5�� 6��6�y�����Љ	48Ԏ4+�޶0�!7bm+6ޚö�YF6&Sf65cc6�(w7�����
#�:pԶ^���2$�6؄
5�WS6��5h�"5jF�5D}~�C��5��R���\�]�6ơ�@�#6�!�6�j��z� 7�]���;d6�Z�6
��6�f��dPص5�6ě8�,I����S��$M7��f64G97BU7�W�6�t��F6�,��9��6= b7���6a6"���l�R��51�W��� �@�4�ρ��=7t���P7`3�д��5�6"Vp� s�5_ݸ���W��7 +�����6�pf����,������� 6�V7۬�����6�:|5���5^��5���6��6�֕6$Eʹ@sQ4��5$��6ꂴ��6�9��"8:5�4� �xv�5�d�6|õr��5*�5>��5x�T5���x��4�q6�16n�q�������6^$��)@�5\&�0��5 A#���3^6��6��6*Ŷ�7��ȗ6(Kn�uo��Pr�5��#6hz���Y56�8:�"xW6.mP��\�ȃ�����5K���e�5@A벸���-_6�S�H�t���)5��굚�\5 b�4<��4���. 6b<��#��9�O5|��5+*60�6_Ҷ���7�6k��������5bർ��5t���B]�{�s	�*�f5@?Q�\��B@&6-i5�s�h|�R��4�i���IX�`6��,ϣ��6��)6R\��7P���A������	5Xh���6o^�5��4l4�4[/S��i�5�'���5�@���T��d��4�@��>Y�5e@�h�/6���5nɵ ؛�7�?��0�5���2vA����j�i6r&������j׵�Y62y6<����5���4������������@k6��µ�Cf6�2�5�-���
�*�A6�¶���5�K�6��	�T	�5��48?����4)��6���5�IC4�Z�54X��ţ�f�G�(l�6�ݲ4-��N�$�V�4��q���ϴ�Đ�h	�@R� �H5r'5�Yb58�	6�~5pF5e�<��3���y@6l�������@+����40�R�,���?6e�	�@u���?���5�KK��''6�7�V�|51i9�0ގ4&��5�I������K76@\�3�2s6�MX�"6ȵs"6ŏ�62�m�ۓ��h��4<6>���;���5��'���[�
��6�c��|*ڵ@�2����{cɵ���`�b��X��&�5/Dy���3�9ʵVB 6����tM�����μ���g��	N��I@6>�µ�Z��E%5��(��kg5+�$6���6&�|��/�53U����5���-6��s�����M>�6Do���\6�a�4�1����6�qr4�Ӷ�,:�����h�5?�1�:�I���p�`T6�~q5�h]2��06x����5�ѵ�Ӄ�|ѵ1�:����5$k��:��n5 }�"�5��@���(5��6�E��^*�5�ġ5:|P���Y6{�6��µ@��P�N��5���6l�U�p#68�S�0�4�N��� ����������6~Ħ�k�PU�4�}��F!6{�����W6Q�� X�4�G5:S�5 ]�5Lm`��m95@���>|:6�6(��5_1ƴ�xV4ޭ*��<5U�䶜Q�6�Z�4�,��G����W4���5�
�����ʄ��Y��T3x�5K9�6��K�86G2�+��܂N5P/s��X7��^�5�q�5�㯵��c��wO�6ñ'6�d7�0�潫5c75��3��W6$����<66C�5ȶ�"F6����
4�ܝ5�96$.�����5�>��Ƚ��0�5���4b�6d:C���`3�lƵ�P�5u�5�ݵ3\�5:�66V��w3b�O��6��Ǵ
�5�h)�vɇ�B�������.���-��봡��5_����е�6�/��l��5��&նe%5}-1���_�\���Q�P6�W�6����њ6`�׳���5�^]5��7�u��~�6�t*6#���hsе2좵&aw�׈�������L5��5י6������j�6�%�6MXJ�v�f��5�8�,Q�5��n4�u�6�^���k}��"���y�5X���60��չ�dJ�55(��@��7�A����7$6�Sc6:�6���V�6(kW���6*BE��4���h�5B�i6\�)��S��C6����>�XƵp���rd��4_�68��4��&��\�6�D�5��6���2��I�b�	6�}��P�5b\}���6I�*��dN�P}6ys�5as�6�F*�`�6�jD�<�F5I{36Ӂ��6v:$6��x��)�6$�5��@�>��5 _��46Po�4� 6o��5���n��[u6���t�6�_�3M��pa�6�R��6���6������!�����X�05h5�)p���[7D��L��5G��6^�r�@�/�`�����4j�7Ц�3�V�r!96���6��5��6T�5�WY6��	�|��c�6Xm�5hĠ�h�\�p����5ɒ���&J6�i[��k<50*�5�7y�����<�2�d��5���5�W�6���6c�۶������7d�6ޗѶ��&�lM6jc86�N1��v��(G�5��Y��&]��6ج[�xK6��5�z�6�9#�0�Z���t���"��O�6�Е�O���&·�֗0��Q�6��R6<f�4�t�6<e}�h��5B�˵@�^��L-��[#6���3�(5`����_:�!�$����6�x��$I��^����4&�66ă6Z!1�'Ѷ�g7E�����N������`���]�o��5bQ6��5l�64$����6�?�6px�5��7t�p���W6�� 60���Je�6<��6*�ζs6�o �\�#6F?67��57��9��i^���� ���^�D����N�B�6j=���07��6N�6�6�E�6���b�����@�P(� Q|4!N4�ؓ�NC6�����5��� }I�t3�g}d6j%ܶ2[]5{B���q87��ڶ�����]���?/5<�Q6n��6�v�1$�6�E�5 �[5��6E��D#ݶ�&�����6c!Ŷ�v�5ls6j����J���6��K�������V����Z�]6�hT���@? 5��˶�6k6G�6��^�\���֛�6Tjζ���6x
7����_�Y�Z�d���[5�N�64Ý�&��5�a۵$^�k��5i���I����q5��5HA�6y����I�D�z�H����$��`��`K<��u�����Y�,6���n�6��5^�5�Z�5(z�5�.��N��Og�~����
�r'���[26^�57%6�y��l@�6�.���~�b�R��ѶD�6 �5�H5|}6��5�]>5n��Ό���3��q�������R6����0��n����L�5�5���Ϫ��Q-�<��6���5��ɵ*�p����5l^���<��µ �2��̶���5�4��5#ᵖtH6��6�h6 �S�㦭�&�Ҷ�j6 �/65�Ѷż�&�6K�?6���6u^�6�ӵL��g�5Ů6��37(���6�Ĳ�jY�5����L16���5{��6G{,6��6e��wԳ�Pթ4�\�5�Ӿ6�{58�-�t4�2�6�N�4����2�[��nյ���2Ĵ�60񱶥e�5�S���-�9�6�sg�0��4� �6O�l�6�~�6����6q�:6�86��Q6p��4P���4T%~6p7� � 7��H5��6�� 6ک<�\�5�Пl�ԁ�6E�6f�:6�5,����|�XDڴ�/5�R�6,�'�T�6�;߶�-�5�}62g�����5�5�s�5�ٵ�[���Kϴ�a;5�Sc��i�6��n5��6ˌg6�.5�r6NG�6@�C4���5��5���5���4��o��É4�y���>���K6����7kҡ6d�m�-�'6�K,5Wל6��50Ӷ�Z�9�25�xĵ�sH6d5>6(�s5�8��6`"5���4W$���W5D��5���5IO�Hޓ�v�����24$*H6�(3��!�5�w?��sH�&:�6�Y�5h�55@��6�\5���6��� @J/���	�6��Z�,����d�\��yF6�E�5Ƽ0�6&�74f�H���g6�tL5E��5�����-��dy���v���4"˴`�4�и�����-���s���%45 o|��ח�is���%`� Yc�\)m��o�5t�h�_�>6j�����s���B�>Q���m5�d��I�5m@^6�����ߵ(�дr�g6vf���5��k�/M6׵�5�6�L�4Ʒ�6��6�ض�6r�3�x|����h� -��(��i5�5�6H��3Ow?��]�6�ݶ/����dS�@�?3S0M7��� Jb���7��6/�b6�T��ۧ6V�7[��ߵ�E�����3;Ɲ6zC�²�6y���Ƶ)��j�7\o��q���wr7m686H}5��ֶ��5F��J����6�����jTʵ����]�/}�6H��6}`�6V�Ѷ�ϐ�E�6GX6�����j���66���8�c� 7y��6R�z6��7Ƌ06�#i5��@�Hk��K65�=7
+i�)�$rD��8ԵwB���@6x�A6��6�j��s�3�,��S�7	�B�4��6�M�5��X�bJ�60;�4��p���*4��7��x�)�������>57�F��=7Ȩ6��/7ʶ��Ͷ0͖��岶*��5��6bS�6R�(ߗ���D?6tH��y�s�	����E�'7�:�5�YU��T�6��7e�&����Q��7Lw6K��A��67�R��~�J޶;՗6�:1��g�����7�zn�]B�6p��s�$�^����|h5�
�4�ж��6f�7�6����`��N��6p�c��@��3��60/����e,76��25b�Ҷ�����j�67T����5�M�5P��P6,���v���y҄6� ^���&��/�2���6 w`�,�7���5�7l�j6x�6�L6|7}2�����B�)7���6�Ÿ��p��v�&7��u6�8I4@'ζ$i����m��6�r׵=�X6|��5��9�B�M4 �H5�U����	�6��6ؼ'��Ѷ|�v6{����6��D6�S�wx�6V�4��U���7x=ڵM)���_w5N�W��rGZ��5��9l���p�l"y6�k��'�5�
��%r�z���,�L�Pѳ:�"�����5)66��>6x�o����4����;d�<����0�O�S����߶�hmɵ�ζ�fy�er
6_6��"i�5n�.6��l5��6Z:7�Đ5.��5�6��ܴ�}s�i;�ԝ0��E�@���DT'��[�7!�?7ja�6�L�6�z��H�067l68���j}7x��N�µ��'��v��L�67�q6�F6���4��C5�G�5WŃ6���6��4��P[�6Tρ6�.����5���Z��6&��6M��6^�X�5���6r�66`�ŵ3����2�5':˶�GѴ3F�6@,�5�����c�����
���
�6oE�6�15��!�s��6�o����z^	��S46����qy�	�{l��ׄ�(�6��I�K�/�x5�6�ĸ����b�o���6���5F#6$�ö��{��C5��ζi�µ�5�5
7�6��S�h�5^P趀+�5�6!���t6ޅ���n¶h
�/�)5�Ե�bc6��6۠��,�I5�(5�Q �T��`��6�Ǝ5�a��2-6ė5a��R��5�t6�iֵ$Y�6X٦�K���`��dn�5 RI�K*;���,[���	���ش������/62;�6T�S6�Ͷ8�U6*L
���3�MXA6&ط�%�66*��~�œ�6B���$K6��6,H7a�6�5l�趜�d6q�v����6�f�5��l�zo�6e� �2ɶ��@�nu�5Z>{6���6r����������7�uW�6���6`��Զ�4)�6������K6��6���6z�5�MT��v�6���ו�4��5���6�5N��5"r����j�储6�j�5?�A6lE�6�P�5���5*،6���6L�� ��9ή6���5�d-6m`�6@Xa61�b6�z5\��7�M�5	#7�5�i��5V��8E�(����5�٘�&6U��9���Y4��6w�̵�������5�|I5���3Z9�58�R������>6b��4H�5�26�>25�&5JY����ŵ���&Vj6"?n����6��5(e�5 @65ns6�qf��+r4鰺5k���Ή�5�?��J�����5R�F���3@�<6lf5'���\����T�*�7���Z�,7�w⵴�(� �H3��=5-���Ȯ�6g*7� tZ��y$6ڼ�6>;;��Dj���"��w�6�EN6W�W���5�	Y6ܼU��j7���6�ʶ'j�5�{p6U�7�6�В6
��5�����ƶ�A6���6��6�Z7Ⱥ��e�ӵ7n ��J�6�+��?�6D��5p3t4G�"�_���P�#7���6����������Â���(&6�D�.�(���h6�k7�U5�ً6,�;��­6�ȍ6��S7P��4�^u���5�����p6l7���o�櫠5@o�Dw6�2C���M6LG�3��6@�J4,��5�{̶�pI6/$�60�}52�6�q�*臨�O��x�w5�6�4������6�#6�R����96H����u5����R��4!��Z�H7��-5�866�7�l��x��4���6@M�V����B���˶9ֶ��?�d2�6�/�6)�ٵ���;�ֹ�6�˴b&6Pr����`�@n��֛�6d;�6��R��ڔ���&���'�*��6I۶D�5�N6PX�k{ 7��s�����c��@�4�m�66���D��S4~Zڶ63	7����H�6�T�4�K�6��O6��+6��w�t�1����6�즶�Ց�u9V�������$�U�L�Mb��v�6��I��S�6.��6��6b9�6e	i��P� ��5�5��4��86j�Ŷ ��o�5^
�6j@�6ҷ�U�6�/�6�}���6L5|�	�h�r6��[��r@��64?�6�y7$��������r�y6� $�9!�_��5�[��L̳4 ��4۵�}�6b�#�2��6���4r��;�$7}b�6X�'6(
@5b)ʹ��%6��p�VT���Ts�d@�6>�Q5;Փ5��*7,f&6҃6���6��
7����v7�ﶶɇ��U��-5~�L7�g�6�C����B��5 ˠ�xw�(��6�n�6�j�6��	�7Ő�6�=�4��?���=6�
�6�َ6՘f6��C��v�6H7�6�C��	��A	6 ]6�1�H��5Ȣ*�gx\���7 ��3�.%7a��5��ɶ=Xs��j�5�a��A��6j�!5�O����6�t�6��^���,�V5��6�����{3�,�6�����M�6�4�5�S��'7�r6lL�����@t��o��6��=��:�5���5��Ƕ/��6�b��Π��,�|5`>̶H��r��B[��E^6t���פ6wj����5�!&6�����t�Px�ȵ"6�� �8Ҿ��� 7�e���<5��W��>�(6}.�6;�6���Զ"�~6���4蠓��ɮ5�@�6v�t�������.�6��5���4��6& -7�X6�n6 ��6�b���n5�K�6�5���8E��V7pI5��5Ի�7�o��䊓�L��5V�u��!B�,�B�<6zӪ6�Y�6�V����6o���K�c��]6U�8��w������v6e��6+D����d�5?7G��PM���R�6�5a��5$.P6;%6T����Dt�6�=F6i8��v�46����4���=}6�W/6�`%7�����٘��5�5�'42�5�˄6�T��A�6��?�F�#�6��6r��� c,5��'7ﺵ6�Ͷ�5���5B�6HԶ�w��rj��5���o�6ܶ_r�6��)5��m48x{��7�	\��t�6�W��Ķ!;����7���6�<��:�6�y���d�6�6iǂ6�P'6��]�np�6�Zg5���6H�Ŵ���ш6��5Ӓ,6�#�6��6X��4��5˯�6]�Y�7ތ��ث���:6��G6ȍ7}Ȅ6���{x6,;�5L�~5��d�ie�5�5�5E�3h�ֵ5o6���6����@_u2|�0��ŵ	xn6t��5��*5&�z6�2�4ܶ6�{�5G�6b��5.�>�v��5�46z�߶J��������Ȭٴ첌6��ٶ#����A�����6��4���Y~6;ζon��x�5�Z���n�6����4�x�z;7]�6��6*�$�h�G�B�$6�fG5j�68����C6Ei��D�6�N��z��;x��0���g�6����^5	��"6��6��52`���~V4'��6�x1�x;N��K����5<h%��鄳�KO6����t�6�bճI�=6�ao5�c�����ꈶpfO6p��4F�F�Y�6�������5�77���f`4� &�5��i6���c+�6�(�5���������K6�͵pI_����5��5��o�=86hB��T+\�z]�K/�5��(�����
6�o�6oO4�d4��6�3<4f˼�+���T�4H
����6R�p6u��6�o_���e���M2�4(�>�tw�5��+6Rp �t?ֵ^��4�TA6F�l�]"�5,���c����<6rڎ��屴�D27@�G66��6���6J��6�6�p�@�M0&� �V��	�5|D���孶pt�wf7�XC6Z�>6�I�r�{6:EжG���:D�6(U�6p��6�5|b:�T?46�B�5(�6\m�4L��6`
Ѵ�;{���5���Z��4g�¶n�.6�~4�����17�<䴎h36�6ش���5��K��oj60"�5�(�7�<{5��(��e4����,l75&�6��3��P�6���j�6��B5��6��\��5֟�6`h�4�6QP5��J6@"/�s�6L�����7�
��^g�6;�J��C7���6��f�
��6ZF<���6@{��96T���8��LX�(I=��J_��7e�4��޶'�7�H��Е�D9
6�O�5h��6���5��*��臶	ܤ63��6��Զ%&6��;6���*9P6Z%����H����)�H]�4pT�b���>*�������6,�¶M��4�6�$�3�,��y2���W6�4`�6\��۳5m'� ~�3?�����@5���5Z�&6�?����6ؗ�4q� 7d>��G8����5\,65ۆ��pf6T�"��J5w��f�^5�ӝ4�8�3h�$���&3S 68�촇/�����Z���Z6�k�4�8�,��4�=6��s܄6&
�6(�1�AZ6�5f|�5n�q6�I����"NF6b�H���)6F�6�_�4n�F6F��4 8,��p+6E�'6,C �pf�2x��4�	6T�5�/A6Vٽ6�n�P���|N6ԣҵx#�G�6�����������5{��5dZ7v��R�[035Ⱥk�,��5J�)��5����J��͵j�5��n��C�5 �g�[��6([���\6��	�5gS5�-K�Cş6!Ks6<�:5-�F66:���o�5��5���6 U5��S5@�)3���38�4-V6�S6 �Z3P~40��5�,6��+5I6�ĵ�N�5�z�5&C 5�h[6&���΃5bq4��5�}j��a�� ��6P������4H}~���75]th��w���f3�}i6��Z6��.�^ۺ����3Z4"i�5��5�E�5H�6�pK6��4��;6�y�t�A��Q�5.ڰ���P6�x���A�N4�5sT����5t���~�t���5|CU6���5�o�5�/��4�� �����<��A�5T��d=�l=<�P�C��j�|򅵊6�C��P)���56$�ȶ�6�5D�:�0�����6jj���U��"�x5 3/4��6�y���5�?V6�j5���4���4�K
6��5��Y�׵�_H4����lj����3�mS6�H�5��(6Ri���0O6���h�#�DF5��6�H'65Hs6M��59�*6.7�6t�6��4��5�7 6�{�6 �4��4��ִ(4���6`������`i�5�ߗ�-�X��T�5ǋn6��6̊R��jW���ڵ��X6�a�5��5�6/�q6���5*���^6�_K�xz�5`����T6��5"ȝ5;[䶀�Z6��7Z[6�,a��66��6t�L7��N��u�5�^<7�q��i�O6�0j6L�5!C7���H�-��5�6����x�Ĵ�7 �<6C�"��������6�j�6��&��
7l4F6|�6`!/4��.7��*7���6_�7��y��l	�5H�a6��Ķ�n06��i�����Y+7�L�6��7 ��3�6)6 ��5%U�6�]��R��0��6��$6˪�hxi5��6�R�6�7LM1�t�������M���	�4�5��26���6P"d5�v�58����6n76�7���(���|��6�f���]R��w���7��L7P������7���6��?6����A���5Hy��x	�69����68��
��6���"�#6�ih��R��
[�6p�y5P��5���6X�ٵ��F���aH6�'!�M&n7��"�D��}�7�(� ���v74򲵕�Ŷ@6�3
7g6�ɲ�X6�}
7ɶ�ݶ�×6ӂY6Xan5vD���}�5�7���6�֒�zqZ��r��7���W6�/�6v ��cA#6?6϶�C��zf@��zѶ4N6e��6��5�!AK�$]&�4�6���$&��[	6o�&�$8���6<6x���c/6��A����61��6�.�J��ܵ� ?�/�6���
�4�zN6ID�n'A6���6h�55�Ƅ�`(����7����M7�[�6�%�h�55u�6���4�F56ԯ����<�����I� <��)7.��T�����6S�z�Q���#6L]7�UM7VN�#
 7LN���Q%7���nkN6ld�5L-I6j�C6�#w7Ⱥ5�.<5�/�6�2�6����]7��˶)�<�¡6�qF�%�669�6R���G�5�v�@�������;�&7@����T�!7�F�5�4�ً۶��&��z6�.�7ob�60쇶��u7ـ���#s6fß6�0�Ȁ:5��2� n�3ֹ�6��J���+6]�5�p�X&õ��5(-N4I���T�6 !6y���y�i��5W*6��5��=�ۯ����6@I�4�^���#p6�U�6j�L6
|o6�O7�Ē��766�O����\i6�M�5ps��b[B�O=��nW5��϶��5���D6 �_5�X�X6oT�H��4
@6x�U6�ǧ6r犵���i�p��z�5�Of6l��5�_�6��5�?6��L�%@7�l�5H�Ƶ�禶1�)�̨�6�l(6��K5_G7��4�L#6"Q��86�Y6�ɤ��;6\ ��7���x��r6$��6�;v5N\��At����^�5��� =�4@�	�Z�Y6�*��`��܋A6H�4�D��x:6t��4����3<}4]VQ6���3�Y�Zq6>��6l����e�|{����h6h�35 �R�즉6�<O��D(6\᏶X��5���2?5���۶nu6U_g6�����6��Y6�鵨���`?6j�ٌ�T��5¶XZ��e�5�W��?ŴD׺5 PC��|��Z�6�Y���ж��5��3�`�6On6`vV4��6���3d�~6�J�6`#�6���5 �Ѵ��5��0�1[�����4B����Q4rt�5<W�5��ܶ��W5Й�3�)���6�6�%�5��4y�"6'�6��6ѫ���5*����~�6Y酶@I46��D��6�"��]���8�l5��f��+��p��6���6ȅ���\6���4r�̵ӊj6�vF6�p���6mV�5�w���՛6=���d�96}Jƶf9����5�段���4N���xƅ66t��l����y6�O9��_��@h4/����8�5]�6�#�6���6(�S5���꠶��n����� ��x���k6pXg���4d_y�˭4�	��t"�}�4�ު��r����Ѐ96����{5ސ�5ѥ���6��O�"z���~�K����'��o9����5x�4��6�����2�����4�~k��T�6֕�� t2.[��J��8h����x/�8��5d/e6��|5�.��X ��T	b�}�?�q7v�%5H�����D�Th�/�6�?6>ٵz�6��ε���� ��2^3����P6�F���T�S�^I�s�7=���m�`�ʴ/����W���!.�� ����5E��5�\����U4`�I4@�6�!����3�
e��0K6^f���>*6|��4�/6�k�6PV1�\C~� ^�=y�6�6���Ԉ�w^;6���H���ܴM��_5d�|4�kT65�o�����5.�B]/�zF6n�u���a��b�'���5g�6�h6�Ӂ����5�,�r�,�e�5d
ĵOZR����5�����\6�Ϥ�z�"7Y|6���6н 5,2���96Z���L)
76�6�p����4�ps6fDP��5㵓r�6�<��S5�6lŌ5�15]W�6f��T��a��M<�`��6Op6�W��`6'�6�;���ӌ5�7�7����!�^5ڶP�74����6��Q���6��Q36�1���K��ٶ�&#�7�4Y���bu�5X�!���t<�	�6�^�ʧ�t*i6�.m�%e68&8��HZ6��G�.S'7y낶
ش>�5[�̶�����U��}����p˰����p� 6T�P��;O6��8��!M6g���c�K6�4��S���x��|T�6?�W������G�M�T��B6\�F6xrõ��y6W@��  \��V��̀�GDU��V6A�ȶn{�6^�ܵ����h/6�Y���R�6���6
-86� ���7'7V�2�6ҙ�5J ʵp�4,�66�,�5I�~�(q�B��ē�6�y�6v��aQ�5�U5x��5��G�\n�6==1�µ����I6�D,6X�u6�[7����
6�+�Rb7;�R6 ~2��%6���<�l��6�۵���6�`|6X;�5��6�hܵZ�6JU65��5`��4	(Q6��g6����Ng�@?��W6��� m�5�Z$5n��\�5x]g�O��o��6�:o�&�b%�5r;6��j�xv�b��6�J��O16�2O������Dj5Q���[�����5�d�5_Ƞ��N�R�5@� 3��[�XX����5�g��̨�؟�8��>'��4뵸�*�Nƀ6>K���L�5:������6&n�5��4O��5���6꣤�֜6DH4(�'��#A6��l52'64D5�� ��g)6@��5�^�4�P����6Le5���R4�����b��5���5$��4�K�4 8��Zĵ��]���ֵT�5v�4�~������+R���4x��4���34�g6,[ ���}6ƴ&�ڮ�62�������
B��>5@ص���yi�]�6DK6�ѝ�����G��s��6�H�f��5#Id�Ra'6*cZ�����LA&� �@5.�5�R�6x������r/55�������5��5�m�5@E�4_鋵?G-6���4ɺR��/�4y�6�r��X�^��7۵>c6�v�6R@�5�6i����2�>O5��}�kIQ6�U�*�Z��j�6�b#��816 �M6�BV6bw�5��
6a��6bq��-c������gC6�y6�Wߵ,�v�6���.(���-���F��r�5Л4���5�h��z�6`�����)6�ނ�i6�<�6�\��,G��@��D��6�؊�fd5ZV6&-������L6��_5�c���@�5hMd5�j?6fI�5"��6�6�dƎ�n���M�(���&J�5 ��^���ʵq�7,��5|��x ��hrm�S�6�s5X�6̈�B�'6#��P��4J��5S*�Ĉ!6��_6l�5��,�	3��g.5j�16(��4Dr?��62�s�6 �o4*-˴�옶ڑ�L#��l9��yU��-.����G�^6+�6���Ͼ5�܎���X� ��4�����������;��w6�{�� �p2O�5g2�5�ѳ���5�*���,�T�68�	�b��41�J6�m5����.�7�yp�&�'5�ܘ5&��5p�洏4Y5ډf�$��5�_�5Ǐ�5�y��O9��8���?5p)�4����#{�6]@�a����!6���2�G�$ܪ��r�5�=5�-G�^;}��7]��w�6��v46�4�<!7F��� c'6tM�v+f4D�5��G���6r�X���T5J>�n�˵�]ߵ�n�6C^j������+6P�6� T5�%�4������'���U6Ź�6./96��6�_�3�}]���5��o5`�6�$�o5�o�5�P��`ڴ@���w��8��M����nm��\C�6�&��rE���X�4-�Ӵ�/��1�=6^��5�>��r �5���c��fI��drn����6u�	���e6w�Q����@�(6��66��7 �D#6����#��6}�6�uR�v	{��Å6\�/4 �Y6o4��)62>�5��8MD�58b5��J5��o6�wٵC����f5>�-6W��6.���p�4�1L53w�6�/5Z`�b�$�Pj�4��56�fl6Z�O���~�L%5��t5vw�5�%6���5p�Y��ڪ� ���L�6�s�5�!��4Y�4L*Ƕ�\S�FO����2�|׵9v6O!l�2�s�dW+6�v�� B=56k�6d4[5�C�5cش��J����6�� �����ؼ�5�𾵸l|����6�$D���S4N��5v��6B"-6p�5���3B�63��Q]I646�e6!Ɖ5J��@�;���E6�D(5˂5��6x')6��u5�Wĵ��6��5�:4xU�5��j��7�5�c�6��5p��5ơ6	�5�J���6x�D6�g��#�l�^6|?5�g6Z���HK58�4p(C6�&ܵ0^�5��K��6 `�1�0�5��6��_��+�5�c?��ܖ���8��>5�iݴ��5��6�b6�v`5Jh�6@606�A4�g�6�&e��?����_�t�g�dT��Z��q/��6�y6�}��^k�4��-3���6�]�4D[6�N!����5ՆߵZ\��+�3����������Ƕ�e_5�H�6S�fj(�p�ҳ��6�qE6��!� $���5+s�4�{���F��񢶎R���=�6�����y��5ƭ�5k�P6{R6*v׶��#5�����Ե6�t��PE���z6��˵	�65�'5�ޝ6[ۡ�����p�Ͷ�aL�I7\���b�5"���2�5׽-�Bl���!p5k)6)G7�5�+�� 5%376�|�6�57ŉ�x)����Ƶ?��4=�ǵ;/f5[1�}�5)���N6@6Qk���Ɵ����5���4A-6I�G6��25]�X��͛6�Ԣ4��6���5r�e�/�|�����6��5���O�`6�8���Z��v�6l�N��Q*6�L6��_�24F5H��5�7�Kq5P�6�5<��5G8r��[5���4A��6.�h�j�.��d�
6Q�5D�6�U6�׬�E��5y��5F��6ͫu�V�5Skص�׵:XA4ޞ6�V�5�%Ŷ����
��v �
�6����#5��o�5�8=6ą6���&޽���5�/?��j�4�t��e@ԵC$6z������	14?ŀ4n|�5"�K��5�6�m��,6.��3ί�4$�6�i���B ��Mɳ��\��!6x} 4�?��봦�)�p��5�(��$����1�
6��b6����4�J�3Z$�ZMN5��b�f�]6G����<��e<��A5��K�����s�VQ)�9"�56�G�^��5�V��A?R5���6]����5�aA�5퓶�z3��赟e��dS6Ç���ڇ6��V� ��4���6��5�.�4PNд-]-�f�c6��5
:�6H�^3�����ۛ�1�~6�P�4Q?�5��6S*w� ��1=q��s��6'�J�>��5�z�5}��%��	>I6�<�L9K6�ǽ5Kе��8�i5Z��5<�6t�6B�4�~K\4�ھ6��46�a�5���^ֵ�n7�La�E7�E,���ѵ�vN�$s �*�5���6�a޵*�5�$x�l����L�l��Vm6�����R64w�5�n�4f7��0�����6gi�6a�/7�SڶH%��y�㶰{ôL ��q��5�d6N��6��96��:��60l�6�?��cY�6l�c���	� VW�2$�(��VBO6 ��4�2�6��ֳD�62�r��W67��"p���>ܴX15��E@5٪7Ұ����6Q����6��ŋ�,]�6g�$��$�2m���������t�P��e)5 2�3�Z�5 ҳ���6 )����ŵG��������̶$�65\u&7��!��\�6��6ϗ��c��5�E�6῕6V�q��>	��6XV/�h�7�'յ��6�b�6Z^g���O6��x3~�5 q�w#:6���Lhi6~70�5^@���=�60B��D�	�F��^��>����^�C�H6']�6Ƈ�6�?4��z�H�4N'��ë5�����p�&5���"6S��6X��f�6������ �0A�P��4��a6PN4�0�Zj2�P*�o�j�BD����6`�5�1��Sdp6�"7M&M�7"�6^�/�Q��V��n��6�������$.��`3����O���6���6�eѵj�:5~L^��"�6��6V"�J5���5�<n6 U&����a�ڶئ���6�u�6�ͺ�@{b5��F��6g�/�G�6p�=�1�5��6��䵭G6�-����64�6J�:6�h\6���7�T7��51�6 T@�<~�.V�6���"�ϵ8�	����h)H607u6F��5���6��7ی6�F�6B��d�����JM6��*�ӵ�6�J�\d����5��X���55��6�V�6*]׵Xk56tu�6&�e5�7��p5RN6�Q���6����4�f6^u�6��^6T�m5��1���7� 4l�G��5�`^��y���.��S�݌�d|��2�6��6�H�6�]6��3���6
��I�@����>"6��5X��e�����6�����B�5,Q|6���7���6AL�)���7VQZ�����X������۬7tt��=����5��68z��<��63&�����l�t&6M���H���Ah_6)'=6\Q��j�
6��	7E��|�)�±��.1�6T7C@��^dR��s��mΤ6��۶�Q~6�M���DN3��_���b6B��6�"��K6�M����6p��4�<�T��5�;�5������5;���d���5pp5�6�3�4�?�3�;6,%6-�[6%t:����h��6��86�C6Tb)6:y�6�w�\�G�7T�5(�,6���6�@�4��X���6�1�5}�6�ĸ6C�S55�6 ��6-\)74�T6���6�T�K�6�ƶ��ĵ�3�6ׇ�6����^>�)���8��a�6����t-6������ ���~5TBE5_�36�����Cj5h���973�6��_5���6�DA5�6�i6�I����[�F�4��{�4VYᶪ���ƘZ�[�+7�в���6�����}����6y���䲶�6�p*7`	�5Nϸ�=���Wf6077|�g���b��1�5�1�5�en���5���6� ��p��6���6vdm��bŵjܠ�H76��1�P]��
���F!�� �]4�L���K�$57���U�!6Ow����5�r;6�i%�О��tU�jB�6U/>7�6�7�t#���]������	�8X46���6�ꊶ��P4ȶ��Z5%�X�K�6����ھ��]�6�ų�a=���5�47��n�Bp6k�����j6E��6p����)4�O� .)5�{g6���䨶��6ܿ�2�T6��=��k���Ez� _E5[��6�D�5b�5+�6D��i�/6Ȍ�6s�v��O6������c�y�.6$@����5��6tV��%�5�64��F�6�U��g5�"$�՛5 N6�L�L\6m�t5�l����4�F6H@�TMy6�6�ɪ��{�g����:a5�7�5�gb��k;4�AP5�����5J$	6� x�tP.5�a6K��,��66�7��%�[��j35�+�����m{5�Ks����5��ŴV���Q�e�c���޳5�מ5��5��6���5�R5�C`5���5Q�6T�a6v�461|�5���.�As�5�n6��1����4��0�R
���`��ʹC6hĬ5\��>v�6?��6(�5��Ƶ�1���Y�5#=�5�;|� �(��Q�5������5��59�5h6Y~�6^L��'������6FL;6�晶�p#6߃�
�6Gv�^x�6r&�8���qsS�_��5鈭6��$�2g ���o�p4�5������4?E<6�tN�o���mf��lX5�!6鵼5��5@��6�3� �B��E'6�Y|5 ��3��5��%4N�洒tu5M� 7>[�5�+�nH���x�M�5}(5����~�;6�c�V��5t�G�&�F#�4����U76��(�qk��i�X����@O�d^B6?"�5Ig-��]4e��&=����ŵЁ�6��5�m�������6፵�$i�6|<.�Ț�,�3	붍e�4�U�6p�k5 ]���~3�೫U�5=ު5�y4��5v{���H�f6]aK5P�)�8�~6�oS5�{�����6$���f`��ԃ5,� 6��6��/6`4��ޕ5@�d��YP6P���C�e��eX��,���6E#ᵤ�B��+õU
���K6"�
�Z:L��L�5c%�6�&��ͤ5�k62{�6	ĵ*e���5�}nv�1F6�����r<����5ii5	��5�$6���,̏5$$H����6n�5��5�$�5��2����U,6�,��BQ.5z�3�Qq��ͻ����$�40���g��6"��RnK�VaP6sa�5����x��y�6UY�.w#5�ү��4���6�O6ۙ/6�.�6Z6��I�����b��p���hM6r|,6z�5�=���F��D�{7��6f,�5�V��T���$����~����|r��TI6��P���w6[�!�=0O��:���|�2A5�
%73ѶXE���d���9�6V
j�y�6���4��!5u6�6DD��Z��6D�嶜���5~�쵠u6�ʩ6*9��ϵ2�	��VT��#�6ܙ���iQ6��5��6>1�5�2�3j�	6�5�
�6��յݍ�$x����5�������ⱵJI�4�tC���x�6�4p����5pW<6��q6�xB6�Hf5p��3`ʨ3��ڂ6�? 6S��6k�۵��۵��:6�U�6�dҴ_D4��6�k}��g(6�v�6�4,6r6�7&�0�a�6�j6��.�k87Hb�4�,p�����_A�Tg��V3�6�-���E��8g6�ˡ�7����Z���'� ��rAh6�"�zi6�>ɶ�l��iW6R�"�T��6��N6z�[6:[�6������5w����_!5�7�6���16%�&��	F��;b�(��6���d��6ذ�5�9���e��tl�:d#���5K6<M�5�_v�-յo�6m�6�?�4l.��V
7 Z�3�x��b��4��x�FW�tG�6Xyz6=[���& ��a�5�1K6ٍQ���o6��ֶ,�E6��ò��P�E�<��m�6.Wj6���6v�!6aU���6n$�5$C,�ƥ'���5Ж�6..�7gZ�4���cj5� 6s��C6���q�96��5$�Y�>tJ�`�49�n68�ߵ p�6��5�Iմ�Q�6�5�6���o�����	�D���b,ݶ��5��u48�D��4�"�����X� 7 [;5$)4>o�4z���ô�p�Q='7#|�5@x����6�n����5��6��}�I�ܵ�i�	F5��060ŧ6��Q��ܧ�(s�4r���$6�	 6�G���+���ce��CĶ�1���Nеχ�6��k5^aԵ��N��K����iX��?"�0��6;�H����ψ7�2�6���6^ȶj-ܵ�,�6��i�8��4[kd6� ��ؼ�W1�6��7��J�����4+1%��f��!M���=�p��5z��������5�ƥ5\9�����5��4�ҥ�.�6wݮ���+����R�\6��7�j��hh]�^�>6�>�5a���.�`>��-4�!�����f�5�]�2�S�<̒6�Zܵ���5�J�6j�E�dT��vUԵ��R�Y2�5$�6Q���2��z6H�6d�f�za�5���5�%�5"�47���(�
��t�t��4�/۵���6+��߼��~��X_�5@S�^Y��pִ�rٶ�Fζ�����7̋�6+X��XR�HB5�=�_6�)D��\-��I浧)�6D�T�S�B6��6��ٶ�K�50�U���5��6�v�5��E6� ����A5�t�5��Z6����#\	�&<6,�z5�;�4D}��v&55��6�5r��gI�ۚ�4��Ѵ�����D���7Vֶ&�5���5�J��j�6��_6l�Ķ���j�LA6�D�5*"ȵV-a6�" �f���0X��%�|�H{��d�6�ö�9ʶ�.���5�(��x�+~�5�6
�H6�ʯ��`�6d����6�[Ǵ"���`3��T4/6�׉��sV�v�˵�5���6���5�5��V6$��5nv�׶��O:6(0^��q�z����]�6Z�t�ݛ6�+6�ˈ��L6Yn5D(5�����6�?6,�6���`�0�����`��4@��� T䲚ඔ8�5�j�5��(���^�E�L���u�6 �g�̥�6�J��ou��R6�扵afS66�7�O�� w#����NHQ6�ky��T�r�5Q���:��^��0j����s�E_5Huȴ؃�6�+���~�ȫ�54e/�W����J൞��5�!�5���5���nT�z175:`�5|6E��5�6�5�%�6�@��]|�:pt6Ü?�c� 6������Q����6�=`����6�{5A���$��4���4�&6�nR����v��Z�6V|v6�1���7��씀��Μ��_�4H�>���O����5�� a²��o6��5��X���6M�趐�[4i@�5����v**�ض����4v����1�5:���4�0�ϴ �*�˵�̴��5���5p6�����W6x�U5�!��2x���5�5e��p�5�Ð�H��68(�3a�}6�}�4*�״ƣm���ٴ-mG6m~67������@�/6��7d+� ���`ܵ�#5<(����&C-6( (�����^��5�d��	J�r�/��m��R�6��&�aQ��ޣ�50-O6�
��,�>��6R4�Y�5Н�6�'��j��5NA5�K���������5�5D��k64_p6��T�Lz'5�P�4sv�6�5��B���5x$M6����5�;�6Q��5 �J2�Tϵ���Ґ5�76  J�]��6�Q� ��4�8�O�!�@[�5P����4 I4�0�F5̶�ހ�<A�5D�4:�(6��ص�
c�M��������
e6���-����5��5f��5��*�(~��;5R��4�G���o�5쌠�7�Q5� �6�h�40L�4��5 q�4@N�P�N�����c�06U4�5�3�5��s6t��6�|\�N�����15@��4^֔54�ö �»�����4��������5�u4c:�5ЁM50�A4��'� N����ȵ	[4�m�!���<6X�p�R�͵δL6���7�
�5�X^6*'u6��5�; ���6($� ��ɼ�8�4��5'�O���6�m6�hQ6:��5D]�6��J6�4��6�ߎ6�l*6�ؾ�0fZ4vke���5�0?5�䵒�����76`J3߇�6�̆��N�g6��?���5F����}5O,�.�����6�
ϳ��G5]=6�Ҵ���ﺵ��w4�+5�� 5���6������#�5ff���"���5���4�_*��].6Xq<�4��6�j5c�6b  �$8�5<\5��h���5�����4�f�6�2�4����6��d6L�s�<05�pH�0�ɴ��e6&XV5��4��N6�k6�X$�(�6t�4�*�v���4	<µ�,�5����um4x(�4��=�S��6�E��l���(fµ�=�5&��5jze5s�6.J�5��l6�é5�q��؟�\M6P�5���6��<��`��k�5!�Q����5,J6O�˶S���%�p5���6��5B똴���6��(����q�6�2��ؓ6�B���
�ڍ�61����5���
6����:�մB͑4�R��d�5���)�6��56%�BH
�p�64�/�{sm5�Α5��D�R6�6I���[�>�6lL(�z��4�������5Byd���5�!���15�#66Dq�Y��5j��6��.��%�ڼֶ�n6��k�{݌5 "6fdG6U�ݵ��6�6B��֗��ӵ���5�C*6s�!�\��7]=���^6�0C6`?�3@m^�8Z�5��34�66�6p���)~�6c�5��A1�tݵ��,�T�j�}�5���6
���h�7a�6�� 6���5.�6���~E�5���q��`����3E��60�y�l6��i����R�6�%:5<��4&Y8�Zx��_�5�EJ4�)6t;�q[����s6)�_�����u}��0v>�d��4��F��W�60����64���6�~���+�6E�6`�/��.׵�A6�����N�f�x6��ʶSeW6Z�7���;�365��׵N䣴�7ʵ?,u��긵"�5�"6�M�5`��G��5p�$��01�\��6�2��
�D�͂���6�/����54��6���Xz�4{6#���Q��̵���37T5�.���a^���c�`�Բu�4�������hW�:8
6R��5��i6.K6��%�7���$&�5@��ͱ����F5�n5=�6V-K����4LѦ3!�t5�Gk�R_51���`l6�k���5w�<��e6��6L��4Q���B4��a�62/�׷��`�5�:����+6�-���F�_��4H��C(޶��\1R�a3|�5��µU��=j�D����ŵ�$�5:�������F4��6�F�3foĶ�ʥ�KD5D��2�xyµ�I$6�U���6n���Y4[�6$K6�_6@��(	��x�H��y��\7��5-6��5�c��[�
�P�C�xn6��L5pｶ8S6򽃶�J�����X��6�����S�EO6�(Ƶ����/�6n>96��5O�4쑍5�ր4~Lv��ԥ5E� 5�*x��S뵊7����&6���A��6��R6G�ϵ�<6d4Ĵ>9����4چ<�A�q=�6Z�B5��a6fb��Y��6�@6�.ҵm�6Y��5qh��@Dq5ʫ���5T��69����^6x�06/	���i��r;�����IF�����2
I6BG6<�<6 � �����%�5���5@߾4�׫���6��?3�e26�^��f���?r%6��6��6����RZ���F(���6$��ݤ4Y��5���6}���Ε5O���K����Pӵ
I���N�89�6y��n�6�{R6�Aڵ1t-5v��5�F��A6���:zt6����g��]5�4�6�`����5���6�6���4*e��0���*z6�n�1�5���5��ߵӅ4��E�.�M6®6�vW6��"�+��xd6�;�b▵+&�(;.�<z�4�Κ���/6p�ö�o#6m���(����6S�޶Ke�5ƨ�� �����������l6 剴����h�5�q�6am5J+
6�Q51D15�S5&�o�*z�7��ܴ���_�5Fal�F����{5�A6@�3p���8��$1�&��5�S6�É�y�W5���Jv��6p��>*6n�0� ������/��5@���P��3�q5`�D30 ��4[6Ɵm6@7C6��6-j6n5,��4(����� ����8�3�7��m�5� �����2�h���B6�m2�H�5��J���5̅��Y�6�SP� ��Pҗ5$�n5c�#6�‶�)J6\��5�5�6��5:L�5؎5�cS6�r$�V�6`�����6�6�պ5��6\�#���62�6p:�V9J������j6@=4�jS6�.�؎5X\/�a�5D`봬�ߴ�h5�#)6�F	6N�5��=�h.[�P.f4�b6>F� P�2<n�4F�5T.�5 �M4���5c�V��C6䇎5�?�52[ն��E6�}]��c 67�Z�qӶ��DL6���5��4�H���
�5 }5(ß54I���N4bLz6���t�G�:+6l
�4�0i���εJ�36�m6PSM6�A���K6DЋ5�ȶ�ͨ����5@�-���6�L�d�E5@����386��5��+�9\���X(�P36��6�B6��6�?6Dp���x$����5x�\5��7�G.����� �.6SXǵ���g5�2�d�5�=V�%a�6��!4XA�53��5��5 ��6<$6�4~?I6�15�N�50���T~4��݈�p94��)�	�;6 �6��?�5��5�qp�Ԉ���ԗ5�N6f�W��=����l��8֍6����1_6ԩ�5o���BƵ>ڈ6Ɋ.�/5��J��%�5`h��83%����`�i5��5��t��CR6U�H�^"P�`)����6��4d+H6����������̕�5 T���5@��N����+�tAY�beM5�<ȶ8�:5��5;�@�Xu����+5�v5�#��+�"�гB��VB�2�ϵ۸h6���y'�5�Q05z�T6��^6���5&� 6��X5TU��C�
�5����e��*�Z��5�ꙵ�6��6棯���m�C_6x%5sq�j#��s���Z�4�:���[5��k6x����/��)56��6((����6��6=ܶ����f���ց6Ăm5�0̶dS�4(�)5���6��D�	k�5����"�6����@��0[6-$�6pj�5h#B6X1`��Y6R�F����5;�6��N6��F���O�6I60��5YΫ6D��5��5,Q�����6nܝ6���5��7f�C��=��7��6i����6�؈6r�h6�λ��to6&�6�<d6���5P�m5�y���n��xݜ4��5���6b7�4k爵�+-5xT����6��
��J�6bS�qg�5���4�7%���M�5�r6;�68X�5?S��8�,��R!6�K|�|����5�O���צ�����⊥6�#2��G�Zv7�.ᶕ���=v��CW�8=:5�&�������7��϶Z��?��6���6]�6=�~5C7?���x䇵&E�5�\x4ߤ�64#�@�3��h5:��6(���f��@��˵��1��z�����	�����4.,���7�5F�ζ,����O 6��60�7ʲ��U�ϵ_~����F���t4!��4��� )���G{�bP7���?!7u}6@�84p�#6�86(�Ѷf�ڵ��5ζ�� Ե��Զ0W?7�/�6�O7����rر6�|`5W?�M�07v�6\q63J>6^�����5F��6[Hܶ8Qg��U6�UW�<0�Z|6V�)����6����6e�6�>��Z�6���6t����95��{ݵfC�5�� ���}6$���P	Ե	;����6����G�6�q5�L�6(#6Gݡ6�Q�6đ5v����>v�.��6p���WǶ}>ֵN�1�?\�62�6e��5���1M�6Oɶroc6�_��6��#���׵��h��t۶x/7!bv6͡`����6;�ܶK(6vD6f���+�6ї�6�k�6Xߑ5�1��ί��㘶V���9Z��e����5�p��R��a������6�˛5-�o��	62D`���s���kY��d?жgX�5�	�6�¹�Y�����5�T���=5T ~�ϩV6�7�H�����-6�#�����6 ���Rx��=ö�+��{�68���/W����6`�ѳ�J��_�5��X���0� ��f�?6���8?�`���V�q�068p��oP6V��� 6H��6�S�64W_� ߛ��;Ҷ�?�xpҴe��6)���rF�5�b���AR�*��54��m��6�6X2�0Z�B��_��(�N4 Hn22�^�������6��6 ��6@E��颉6�+c�n�,6�����I6�n��'�6���6a>6�ȶ�ꤶAI6T��65c	7�Ap���95@��5u9�5V��6��5�;:6���4��)6���5���06�k�6���6��<6��5!�6�ǣ�8ʻ��D�5���6�����礶�4��n��jq�4Uֵ�VJ61aA67�a�my��*D�5�	�4 �C65O��-!�$��J뒶\�"6�rM6���5}��6���34�5"6X5.�,�ކ6�)���H�<4�޽Ͷ�c��P�$52��B�7����ƥ6���6�,s��[�6��7�6Z�M4��5�ǵ �V3d��5�ض��<�H�l ��n����S�Ȼ6�������6te�6�~<�CR��i���A~�6D��@'�4���4��k� �3��t�ll���ǳ4A����Ѵ�)�6�}|5 �״\(577$�5�)6�R�57"��6ͭ���6ڼ`6`}!7�Z�6�W�ʞ���޾��q�6��%6Bl�5pw5�Ԧ�����pu�v��6�8 �Z�"7#�6��?6Y��6�1���2��zf�b����<=65��Z�7ʖ�襃6�Jm6�k��@~4�Ʈ��G�60����6�x�5�S�6�I6�t�V�5�s�6�#7��6eZ7�����St5_��5�2[5P��м��=�58�(4/�\� �2�K�5�X�5�]X� �r� ���w�7�>/�kv7���5��|5VV4v���������e�`I65�lt�:h.5j�O6��Z6�B�5>���>!6�zt�@E�5gw��55���5�4K6�/�؈�5n3��ѵ�9?60H�5~k��q��1�5�X���^�����5|T�5�56��j�E�N6V6�� �"t5Z��٣86��36*6@�\+@�&�	6�v4~y!���=3��6n�5��N3d8��] ��7I�#���ѵ�6�4 6�o�����VT6�5�SƵ�t�_n�6�W�<�Q6���4��5ddִ�5V.]������5,��5`6��A�96`������ۺ��͡��҄6�	6�!v�p4r�?56ܨ�5J�ֵ���5s��5��5�8X6�t�����y7C�Z6� �5ŕ� ���F3�4��[�5�i%���_�O�86v� 6�`� ��29p�4���f䨶�XH��r������F�{v6�����A4�%�6�t�s5rJ.���Զ2`7��9�505ɴ�Vw6���5,g���,q�͡5>�5 �4D�7�	ܵ��
� *|��FN�!H5Co���`鴞��6Ļ�6��G����DX96(�5����̹�j^5 �6ཝ�S�l6�]%54(�6^87�^450��5�
�6T(�hN��Сv���5�(��@յ�r´"��5�1%5��6T[6�Ȧ�P��5�۝��4��4 s��{6�~X�T3�K��5܉5h^5t�5��l6N��5���}��5��µ\e�6h-��U���TY�(x��^��6Л?5Zm6� ���g5*,g�o��
��6����u�=L�6��ѵV��5�r>6$\T��w4����6��� �a�]ދ��v�4菏�'�6z=5�O�48b��0�s��m5�ٵ���5�<"6�3I��+�6�ޖ� :H5T���Bꐶ*���u�����x���)6x���D F6xK�4�@�6�7��H�-6hM�5��5��������\v�Y6b�	���5}� 7��6�w}5��6�6�986~$�5�~�6��R6x%������ק���ɭ5��6��9��6ɧ�6Sݬ6����R7۶>�7��6�(�5PS24 46��G?�6Т�6Ԧ5�p��ۡ5`6�8�r�5�[���{�40Uq��E6���6Ѷ����6�aj�*���>�[6Q(�6�����D5���o��5�"�b2���S���k	7��6��ҵ-���7�b��5��6lc6������6�]���5�.��VDc�ٙ%6
7D�E���I/�R�*6����y:��g�����?�5H��6��ɶ_��4b�}�*t�6Xy�D����0��w���� 6��쵊�`7t�hM���1K�9�A��oж8g൯�w��H��6$��Oz��˟�6�T�5��讞6��	����6�J)6H3�5����٢6F���vMH����6��6HǶ�叵v�54 7t贇ň�l��������U�(� ���
���7L�.���	6Nd�����'H�6��e6�O�7@I83��G5����Ά��◾��W,6P'4E�22�ܵ[V�6/��،�u�X76��P6Q��5ڸ���~�3�-�6@'��������4��5S�.�6����e6�Y6�G�6�fC6�
[��$7�6�4���6�4��G6�2���5F��6<766��6�M�5��v��?���gT6�8�6��M7�>C�H6!65����ɣ6?S
7sP�6BVo5#�f6�e76�������v�6a�n�L�74Q6���5��6�Y�jH'���6D�;4H�2�������6_�S66!��:6D9�"��61Na6�ҕ5��ն��4�&6��Y5 N?6�b�6�x6�r�35
+��b'{5��O�6n�6H��6����|~6��6	�n���67��'6 m�2��}��+�[4�Eݵ��δ��e5��c6���ۃ�5@�5F*\��鵈�y6P8�d@%�r��5����E6v�6�q� �ֵᮁ6%"��B(۶jˬ6��4&���k��J8��x/y5�͙5�߮�K�65}v6`GA6�ﾵf��&�56�$�6��`��)��4(�6�1\�C���:h6�h�5��Y��6p-�4W5���30G6��)�HG_50���@X�@�3`hU�MH��0ڜ�H86�0ŵ8���y������4i��6�6ڶBUN�<R�5�Y�6.5��4Z6�>6�(����5��y��Ϛ6�ڇ���6��(��-�6/*�6��6�� 4@8�2꒓��͜6�-�6f>��m5���<�ڵkYt6��x�׵٪6&�6�x6�Ŵ +I�b�6v0'���'�}�����p5L�}6�)6U/�5�R����A�126��6�#���i60��5�É���$6�6��5�,(��x�@V�4fH
62!��ؿ���'M6�}���46�J���,��6����.�����6|_i���g6�/�=�Ŷ�#�5�i���6�$�6״���6���Ҹ�5��6H��`(2�hwc�Uu5�'2� ˂���H���5�u�6�A4+�6�Q���|5Dr6��{6(�����5� 66"6�|�6��µ��6��3�r��B�}&a6:R��o�6��F�p�����J0ĵ���5�-�5��z6�B�%�Զ<��5l�6`��6W������6������_���V�"�n6�dB�<�L5v\�6�7F5ئ&�7y����v�Y�46�w�68�4�>㴄��h�$ߵ���5�궳`��3E�ӵ�55d޸��YB6���5G%)68�49^>6��]�$�|5�P6 #�4�J�6�ؕ����43�G5�*Q�pХ5�0����S6P��3	�_���@6\*5�8�5XK�U�P���մ��h���L6`�)���C�IjB6��,��5.�6X<��X��4JE��Ԓ���W��ؚ6���5�mѳ�iQ6�����75|�̴>\_�n�/���m6p�q4C�5�a5��4�6^0����u�E*����N6�C�4`�j��΋������K���63�6������5�z14�����5�&%��d�����"e�66p�rqc��Z5���B�ߵ���5C�r���4����mw�M���[ٴbYz6�t�65%�6�	5�[��l�3��ֶ3��6h�6�t輳�H��B�6zR`��K�4%Ω�z��4x��6�vѵ�5Ѷp:��96U=��}��}�5� ��žൖ�7�mζ�߳�o4�k���/cI6U�T�B۵f.���$1� �4��2��K2������H�j�j�q6Y�6"�5kq�5B�}6�t%���'5l�N���=6W�<�����D�6H�����6� ��N�4�=U6a��Ay�6��6I3�6I�i6,Jd�>i���6	ݥ6�z6�����,�4�l�Ś��Db6�5�ն׻T6�2K��s���6� 6^$�6������]�z6��S5��ݴ���6�uA62x���s5v+�6�$��1��H���L�����6���p�5Ǎ��[��w�6F��6���(03'Ի5|g��n̷6�؎5?��6�����6A��Y��4o�ĵUɏ���J��6(�E����Ҿ4f�46(	62Z�6-&��~A�4~��6���6�B{���صoζ;�_�a�B��5vs6`�˶����'z6�iݵo��5�5�Y3�ݪ�5 �/6��c��3&� 4_�U~6A��$�Y6x����J\5��5���6O��5�,6�U�5C���L��5�(�5v��5�Ln�V�7z������83������4�n�5U���Y7�V�6+v��Q��6�^[5ď�ԏ�6�f(��R�B�?6���5jfw�175�2�..�4u5��5��I6���5�"c6���_3tH9��W��W�~6�66�����6r`���~5ȷ�4�H�5q��D�5�>䵿f�6�h6�㶼�*��@��3��c6�����6��C�4:�5���k�;u6+0���!5D��5e�p��خ5���6�lW6�v�*��5$�h��l5��r5�ῶ��45�4D�E�����Q��į�"1�&̼6T ٴ~E(6�+6d�|��J!3U�47�kq��A�5 d$�O��5��C���Ru���e�5ۗ7�50G�2�a�6"�{�5V=Y6�3��j�a6 M�2�h����6 ���{^�6����kr�:��M�5�PK6�6f��5N���<r�5�̒5�U�4�Դ�;.5��x�μX5�A�4鰖6�$u5R�5 �i�G�5��M�
�p����9�4���5ĥ>�SC�5��˶%Z76�x��,�4v�B6��5�I��ta��Jr��5��=v6�b�'�'���`�� 
�Y���8�~�95V�5x�56���Ϋ����6-S�5H�04�)�4*%���<�5$����@q76��K6@�4�l�4@qS6d*�4&264�=�O���i��6�6|�Z��`��@�4��[5���5JeR5�ص�"�59�6�×���3�ke�N����A%����3��ڵ�,������7��$I�d����4ۧ�F׆6�l6�>�6�V�5P=g6 {,4���3�$�5@��5�[6l��2�_5�익K/5c���M|6��6��6	Ϋ5��6�-�5֥b���6�=�l
K�����))����O�5jz���P�5n���,>�5Z|��N�5���6c$6�7��j�*������p5i)��~B%5nBK6��5Xk�5ri:�N �	0�B��5 �.4�ʆ5� 5����=�5�+��eǂ5��e5�6i955�辶@hw���0�/�p�| ���83��QY6��5�)����Ƶ\9�4�-�5��_�� n�N��4��5����&��j�S64�w�HR����c_5���0u5g����4 ?�6�d�5R7�����5�	�p��j�26��D�d��6z�L6�|6 xv0�U�6[#�6�}F6 {�3�!��a�5}��5�k��d�=6���5�6T�l���˶�N-6�eJ6
)�]�^�¾!��^��-�1�I6�f���݊5^��6�$64�F6�6B��&�`��4�U�6�I�d���5ِR6����@���R6�u�Hz=6���`-4L�|�OO�`�5��$4��5k�6\�P6*p��-��,66�]µ�����G�4���5 �H�q�6jpT��吵`U-4�[��v�����#6��P6S��y$�6�\�*Q^6�ל���V5�M���c6�� 6b� 6��	6@�4�Kn���M��?�4&S�6��.6�0<5�׵���F�g6���@Ě3�6��6�����l���(�4�(��ĭ�6B�6삹����4o���ԡ6E�5�ٝ�4JH5I⏶1L75�H�5n<5 ӥ�zz'�J=5�<3�g��C���@�5�Ķ[��6��޶A�Ѷ�����鯶t�6ݹK6!MT�,r��B6h0������4^���#�5�A�6�X=�i����M&6޸õ�{ӵ���W�e�� ���� ��6�|��ߑ�4ו��C ���+��y"6�!6,��62[�t����M6v0����P6h�5[��v6^4��ܳP�۵�0O54�k6�����e6hG��>}K���3H%�Bn�5>L��׵N��L>4X�4��6`f��6�aS�d�[5h� 5��o�7:[6�(n5�@������U�6�q�5�*6���0�x60|a�l�˵xF��D��5F\d6o`5�6@�"�)�6ȳ����7A"}�`�&���q��e� )�j:6�����6�Ͷ�
�6 %�2�o�4Q�4|��]��5I�=��.6��X���p5�9v4>Z4�ȥ�n� �N�S�>�Q�$��5H�k�Q���k�~6�W��D�H5�Ӌ5�^��L�4x�&��gw�H:�4���5����6 �2������u��f�m��PD6ز�c��b���#��R8��M꫶��6�����6���5*�2��c��5:V5�=6&���\54�15;zh�A/���ʴ�G�5�9ǳ�����"��^Y5m�4���6�Y5���4��n�X)z��8"60� 5�ڵz�W6�7��h5q��5~������"a96D�;6G��Z��#G�����6�3�mx5�6���J�{����6iw7�Е5�4v����`qU��U5@\�07���62*�6�â5�F<�(�V�@��6����9�6��!�>���S"6�RN�B��4��`������6���3��6�%���]6|&��LH��@��4N�6m쩶 N�5F��6�߿3�О5���Դ �z�8�J6<�����4hY������5ٗ�����5��=5����l!5�6����1����}4��ִ�憵b�@6P��4�x�5�=j6�µ8ܚ�C㌵(U5L\�eO�@�4�՛65�|6���5����� �6�4�572�8x 4N����3WL�S;6]�E6��L��5��5,�صM�Z6�E{��M�5�r*����ȢB6H$U��7�4ڵ]��6��6:�5:��5��_5�M5��PT6��6�y6���3�5qX6��7� �8��;�5���6�9��Z�6k�5I6ɨZ����%3/�0Lp4 P 3�̂�;��6���6��˵�̆68��5Ҧ7�ǉ+6�H��s�5�N�8�D6j�ʵ���7��5��ʶ �6�{�64ą5���&F�4q���o'6�Z�jpn��360��4�4K4��6����j�R�+��6B:��<!"���5i�]��#i�e�6dޑ��=w6Э96���6(s25g�6O(5$�A�RL	�*҈���5��f���U6x,�4r�6��5���30��4��&7���6D������]�6������6���4�e����̞6�-�O[~6��6�96�ǐ�8��<4��i��k_56GA�����<.�6�����5�6^>�<27��;5En\6~��5��<�<J5��w6@i�3����{�����,�7���/�6�0�5��6zC�6���q,������7�� ���u��G*6��"5����U
7��<6f9�"��6ށ��ߌI�8-6�ĝ�>�6��16�w6,gônM3�xW5��5f����އ6��n5�˶P�5 J*5�?!5��n���ش��ŵ�#N6�h��,q�5ROf�.#�6�p�6T��68p����5 ��1��5<:Q�3�7���6��'6��6|��5.X��0�5JᇵP�S6��5S�6΅��h�5��(7d=��87?6�E����]�kD�3�o6��6 ƱL�X5}�8��ط5>�(6^���ص�Q�5����´����5���5�>�6���5������6
/�6z�p�!h�6Ih]����������*5�F�6�	ܵ5^��$
�ᾶB{6)V �)�+��eZ6x!3� ���f�6�9õ�1�4��궄����5��P�A��6g|6Z�6��o6����b�D4j�G6�VZ�p,��**����5�? �y�ĵ����`}<6聆6�k浦{�5����e`���4 `� ��3X!;6 �2b�G�
6aϰ5�5V�6�%6�^]���?�ZJ:���\6� �4��-�PIX��ki5�8��v(6����n��xr5�S���N���2�6`g�5$륵��"5�5K��� H6Қ~6N� 6aH�5�3Ե@�����u�j��5d.5m��6�6���}�ڵ���Ť5؍*5v�6�ࣴN��5`~����6���5vWz4�6�C��Z.Z6�	I6Vy��wĶr��6!L�6¾5X�5\�B6����v�s��я6�7 ���4J�6��T6�6@��7*�5��q�r	/����3U�6��5|�b��ñ6�"ǵ�\�5(ʇ5�y!5�����16��\��	5p��4
\�5���`u�2�X��q�5k�:�˞�	��,66\$�5�s5��6ۅ��n �54�������aQ�5��4�%���+6�4�4Q����� ��6ݝ6D'5>�յ��T�T�E60��������5�E��������l[N642� 9�(;��h즶c����5�T5�􉶜�յ�	���֟�^8��(Ҷ�^6��;�[	�6"ó��;g��
6Z��5\B���򒵹��@0�6�v��,i4�.6��P�<B|5h�\���r���ڶ�`E6��~�����牱5&�*6] ��#��5�(���T�̢�6�!�� �6xQ{��~���}6�D�5"^�|�36�����1�5j�I65�K6��4��p�����Ƶ���5x]��s� 6$��ZT+6�������5�s�4u���&遶��)6�,�4[�57� a�5Z�5�,���5�KM�q��5�٪�L� �46q"�5�H���(4���6����Jĵ�g�6.3�5��o��$��}����P�����5�~��`o���!���6�:�$^��x�����t�v�5t�&4{��{�5zـ4�6�5ɵ�5�d�(%�+���>��5�x$5�6W5f��5J�$�S����06�b���56����4�\е8�t�\��5p7�!PԵ�5��ֵX�i���L5��\�0��5��´Y�x6�6:�6��z��N�6�^
��zW��V�����а���
7�r.5t�J�ĺ�6Y�5�;6@�X5�'����$����5�0�6�kĵ�Q5��6�H5W1�T�6F��5�����4<Kܴ%�o�O�l��W6Y��5`&/6|�ٴ]�ͪ�6tm��%��5|~_63X�5�36䅫�o�H6��,�6���5`j�5_�赠֝6�{���]��n3@�F3+�V6��6�/�ڌo5(p�i����5������52���� �3h_��R�������r��5{�c�� D� �8�v4��83C6�(�p�5elT�l��5�!�5��H6񗅶댝6��L� #}2\n~�w����Ug6 rX4CZB���52�i5@6�#���5���5]�����~��j6K�i���p6��5��W5*��6�*d��PP6ha7� �?��
o6
sr6 'ҳ�굈���G5�>�� a4@�̳4Ň��L	�늉�ZO��z	68Ƴ� G(�7�0�U26��
��3䶸�յ椶�oa5 �?�K�5�ɚ5f0��(�����;����
���2���5"��g5P(#5t2z���7�5ӳ 2��gO���Ꮅ�:�й�5 �Y6�~5|�<�����|�6-h46��&��D�`	5{��5�i2���5|��T�5$�E5�/����$6"a5W2��&œ68bE�.�R6�!���}� ��4RY~62T.6�G�5���54Ͷ �w��B�5b��6`'�4_6�H�5h�6l���� �6�v5Ķ����絢>)6�x���@6�:ֵJ^ ����4pQ�4�q`5����	$�6��)�6�C��sT�>6�5 ��1`��{�5��ƶ�ʺ��My���6m���� c��8�6 �$�CJ��h�6�3���}��@�6d#���}P���ƴEgP�4�{6��%��*�5���5��W��f�6�6��F6�%6d^6��W�X��5\�5,�J��c+6D$(��)�� h��zI��4���C�5I� 5�l�5@�(6ʆ�v��>m���l�{�,6�1 6]p#�_��b��X��x젵/����6Hu�5��Ŵ�����#� ڇ���5��X6�Ǵ�`�6`R�O�7�>6�Vz6DY)7X����D������m#h�Qa����7���ݤ5��6��L�c��"�k6D�е���6h0�5�a���ތ6;�P35�*P5 xO4��6>9� }6<k5��B6��76�N5��~67�� 5Z��@5D��;�ɵ���6�"�!@B6FA�6��)6K�)��LB7���5J$�5��,60�15�E6 �5o�����v����<`6�댶 ��3��v=y������Iﶦ)�6�W����H���p�ͮ��J����3|�PJ�5�C��-u�5������6L$�6�t��}�LO�5�f�{P6�B5�hZ�9���f5P%��'A�x2����6�A^�~26 Ҕ�z�O����5��6b�~6�u���z�  H1L�[�n�"6����ZBt6��ö`��5Ĉ�6`v�6�i�֍6�<Ŷ,w���`w6��6����ס5hq�6��� ���ZŶ���6��C6���5T޲��w� �}�S��%��5� ��{�X��4�5Ћ?5N�	6 _f��!|6H�4��ж��4��5��4�K�6@��3�N6@w��rH��г6��N6�7z9M6P��5�+�5.@��+6F���u�6�"�5�*�){�62���6���6C�6�,4~�	6YɵE� 6d8H���5Ji6,bO6؂���C�ƀ�F^�5��G� �j���J6�����x�� ,�6m+��X4�����X�Ǎ��M��G�6 lJ2F
صĩ�6�m�2
�<��٥6��S�>��6�x�5X;a����L�(�|���O����p�]R7���]�6���6B�t����5:!-7���N6<����?6�H��ƛ6�v�����4.�v��ۺ6Gau6"jV�b��5U�@���[5X&26�~�����6�460Pa�$��5 �55��X�*V�6й��ES�6����v���
�x��5ИM6e�D��5��>7��|3��Z6t�X4��6\�P6�>���6d�	6.��6.�5��1�7�A�<QO6)�6R�6��Y�(r�5H�'�8侵T��5������2���6w��6x�*6#��6��?�&���6_���(���i�n8n6���1�x�"6� 4���&5ʪc6r�6Ȉ~5 `��t6R�6�]~6D@��Ѧ5�B86'K6��Ǵ")(6�A���(��:d� a:��D>6@�g5�%����K�

�6Hʁ���q6�	6��4����)61_���l�Z4�6��t�-5��T������6�P6*Op� �O6�H6�+5�9ʵX�m6����4�5�9N����5YN��8dV6�7�6��p0޴�J�5�t95�f������n�s�����W��XP6:�|������96&��L�3�Z�5��5�����6�-��W�D�,6[@66��6�B6���6@��3w~��r�6�y���C5"	~�3�x��1��z6�l����5�g��s �6*����Ĵ�<6�(�5�(6~�66�f�����5|�6�6j!���۴Lh'�(X��>ش6V6�p�ǡ6$���4�,ϴxra�&Ao6��.&S�JKL5�7�˶�63���Ƃ�����F����5`�ֵ8�<�Xj�4�^4h�͵?���Ճ����5~����̵Ĭ��<8������.6�ɵ ����"�\2x6���i��5�#6���D9���bL64s6#M6^��Բ?�`���1ѵ|Z6�A���s6p�I5p1T4��5#n
5H����{�5Z"�5p<�N|6�,6�㶍C�6���6p��5M�]�d`�:<6���� W3*�%6r0U6���3v괭��CH���M5`6�LRH6}��6�8�
��6
���l��5���4��@6��6�R��8t�062��;��h6,a6��=J�5 ��5�5�6n3�6���5}�A5��5@�X6cd26@ғ3{�Զ��O�I�6�25����7����5�� ���zs�5r9#�9#���ö��z6��6���H5�p�H���ʧg�sX�60�h4:j�6T�15��µ|<(6j 63A���
!������� d3�M޵.x5L	�6���BK�5 �4�b�55��5�,4F!�5H�ﴚ86ۺ鵔8>6b�5Ɲ�g�4�,�Z�5�.\5+kR��!P�Յ�5>���n�j6D����q��N�6�[b6��3ġ+6R>��%r6��6t�63-	6P�6�島�1�bඈ�$7 b3&�m��ܢ5�.B6��6 ��3̖0��c�6���@P����7<��5�s6V�%��@5���6�v�6�6���u��Zc�6ݹ6� 7U��608��)6�%6�궦�?�Y�6\�h6�¶�{L�6	������#ᵠx�����6^}�����6�S.��n���zk6�H�6a6�v5�����c6B�)6/��5�I�6�e"6�#65�RL�� �5�Ӯ6@v�3嶶<��e�3,�C�x4�5/:^���������$�5��C����:��6�Fǵ*R�5�B���K���ѳ�7�5�����ѡ6�U�5t���5lꪵ�`ڶ�L�5�*x5��p6-�x+,���t���ߵ����.�6�P�5���6�����9�4��6�ܖ4��n��@c���T��ye6|ߟ�P�6�6�"͵��e���ƴ�.W�,�S50+
7��y���?6��ڴ���F�ĵl'#6������,���u��6����I�j�L6P�S�Ƚ������#�@x�6��鶚�5� 7�$��/6�m5����S�6���6VV��-j̵�-���|�6vo�5��5��#7�X^�D�L�{s�|t���J����68���j���oBd5"���%��6�ĥ6��6���i�.6�$����6�8���=�6{l�ݶ̷J6�6�6Y!N����6*�	�8�%6�6�b6���6�А6�.>��J��q5@��3���5S\�n�6�ݴ5�Í�\Z���G��b�6�b�6�6��6�Z6�AN6���5�+�6H�δH��6�r5��-76o�<5l�S5^�N�@w3��44��"6&�37�X6ga7�I6f� �!�7��j�F J6����Wي5�9n�6���5p6��Q��g����5Bnt�F!"6*.��~�#5ŏ�5`l@��,62J�6<h�5Z�?6��26��6t�6�Z�������4P�&5��5��4���@��w66'r����39%6�K�5��x����6�K;�4؅5���5����W�5:|�9,��M����϶�$�x� �t毶��µ�5h(7xN}6f���i�o�T�ϴ0+��ؠ�cep��������y��6�~�$����|�5!�;6^��6/!%�9�w
��w�5��5�a����5"wW��0O6$=5���6���*����)��K�8��6R�˵��k�h*�5\)�6��Ӵ�`6H�s5ū�6
��6�}5=�O���	�l!6�.(��VB6ӵ$��5�k5�V�6�����K�5��M4�6e\��5��F��ن�}K�4԰�4�6����$����6�ڿ5�P��:\�5 S6��6@������6�ZP68qe6��5�0 6\Rx�=��5³06�Q6%�6I�v6X��4)7�6��6P�4Vi�6�������5@��Tc��@�61��6��<5Z��V܉��m6.��5�VV�t��5|��45H��C�6ZA�4h�:�q��� ��5�� ����67W#6 �4<6����6\�`67nö��6���T2$��]�:�_�Ҵ��@C{6����iy5t-6��6�"q6u� ��K<�q��6�6��c6�$����ʵ<�$6�B�6���5ֶ̝�@�5:��6��ֵ �ղ�F9���5�s#70h�3b'��|"�@��
��).6�z7�5�994h�*�Gن�'�w�l�	�J��6�����䡵��T5�+�5�,�5�#׵o}6X74-�^6D���]ˊ7�6E�,��<�3�C��Tb3�"q��y�5�܊6�H��W 64��5|e�5��c5��6��K5���6�
:����p�6��h5��+6�ب5`���4��ݵnW5n��@�U3��6N	�5����j6����2�>6��a��)a����5Xb~�|��5}�Ŷ��6���H�6�������|6
�5���5N�g�8�G5*.�5������F6�U�5%��6� h6tʗ����4A&C60�'�xI��>6�}A�bB6��z�^6h�x6�:�5��5���дf��5ڦe�fk�60�$��>�6]�f4.G#�^=6Ń����6V��zFu�&�36Pcn�U� �'K�6��9�����7ǵ=^��P�6l�;6Eʎ��_5 �쵧��5p��52���I�̒S��#6M�5��5n�6x��4�����r�6�"��fD�����ކl6?'�����>��6� ۴L&��ky4�3�����@�����o6@�6Ěh���D6���44�4�2m��6k�6��4������5n�l5c���0b6t�����3J�06��/�<�6�0%5�ȏ�͗�6	�>6�_�5bqJ���c��w�5��\�4�v�$�����65�6B�6TlT��,h�H��f�R�xU��15 Rµl�l5G��5�߀���H5^:��ª6(R�4�(��X��r�26�������4T3�5�]�8&�|-5Uw�6zd5Ǧ�4�\a������R6����|�5t<�5��d������Y�ҿA5p�1���5Rg6�M�4p�K� ��4�W��<�6X3S6@��4�sf�0Ȉ��R���R�5�V����6&���
��� �ⲬL�w�ڵc���eF�$Q�5,x)6����φ6��4��w68
`52����@62k���M4_M6,V��A51v5Πe��]�5|h��8�6�5c6�X����5��u6e�	�O3�6�U�7���Eֵ�:`���_6Z8�6ph��6���IE���Ͷ5g��
Y���򵠛E�\�y6n�5�B6˜�6p�N4������� 6ȯ��-�5 ힳ,ԧ��.�5���4!|���U5�R�5&{�Rk�q͵0��4�3�����6�= ��n� ���}6�����紤z-6D��5�%�5Z?�T��6I��5 �5��6�4��֡�>��6腨�� ��j����s��2�6 �6�|5(j@�|�M���4Q�(�k�xʇ6V]��z�̖�5���4��U5.))�C癶/��6\6ζ�C���k�� f84��e5z�6�aT5Ȅb�#��5�>6�G5�f:����t���sJ��5v��5�:H�0�H�-�6�$��������5��,5\ˎ��� 5�8�4�i6@��5�'ǶHt�6���4��5���
2�C�����H6�6�i_152��6�5��T1����'6�^�6_1�v[6+����<6�<6���5"-��;��r��?64^Kg�bk5���5�n �Ul6��k4 �0�䠴������ ��3�f+��}�6�wA�ı�H�4fٽ5S�5���735����Q4�8�s5�����p�3���V����6��ȵ�S5�`W5�*�5�^45qֵ�Χ��4ΐ�5��a4b�H=�5?O�6���b���I��1����I�������B5~jj6�;����-4��6*h��'�	6}�4ơ5.y<��d��56�������7��Q�:/ɴ�� �ପ��ۧ6��5LK<����6�	6�Ѿ5�;��2 �6���5@U˳#k���J]���q���P�p�p�F�X4��d4ƨ���<6�/�4�ڲ� �=5ʋ��m�6��U6�����I3��*6`f���;f�,dF6�_���	ϳ���r���"N50,�6��{5�¸4v5�~2��K��e)�67�4d�S�&�5��5��W6�ݴ���5���5d��4�F�@+5H�40�5���O`�Z���u�55�����;����6�s�d��5Z��S�
�ŵʹ϶�_����4xނ� c�3Zi���߶^��61�9�b�X����4�
�6fH`����l�4��24�e��b�R䵰si4v��(Z���FM��Ԓ4��l6ɟT6�wx5��p4&N��jC;��M,6�(�4�l5�{1���5���� :j����3 O(4`�46��6�z��A�D�\)�8��4p&�C�6���5��ζ.7����X�񶌇�6�6O�71�R6�|���}��I綀��}s16h��5V66�5��X�6���5tyj�.�ܴ4��)6Hq۶�Ѷ8�ʴ�T\6=��6iz�[�$6�6b�j6��6z��7��5<���W���5#��5 F�љ�6eCQ60�<�� 5���5�����a-6H��?F���*�|/�4K���1�5�5������ص��[7)�,�< ���6TV6��鶜��5g�#�6��'*������"6�Ќ7� ���9���썶�k����6� �6�j�63�5�x�5�D��O7���6���5��6�u,��*5�x󶲝�6V5�B �6���'���I	�`6�I�2��6���1��6�eV��ö�e6<T:5��6P�#6 7�7v�V����(6��7���6���l��ȶ���53	B6^�e6��6���5G���a-6L{6)$�6�B6`�N�Wyҵ��X6�\j���5O17v��5���P4*����6��7P����6�H��j�;6�pJ6���6,S 6�w����5+�c5|~��
7�J����J�6|�ǵ�5��"�ٶW��|�R�糖��:6�j���6b��Ɩ5�F��Q,6f)5B�G5 �2�c36y6B�6 �P� ������6D�u6�D4o��S5S-�67�z���5 '4 u���$�; %6��B6�+�6���54�����/����W3�6w�46y����6�Yീ�ڳ� =6�J�� �c6��6܏�6wB7(w��'`7���5%b6uZ�6�<��@��3��v6��Y�6h?�U� 7h��6xh67cF|6�E���P�6�%6�����%ж��p6�a6�n��� �3��6�*6�]|5�I����
'���H5�?M���5%��6���������c�5VM6����&.6�q��d�s
7�W�6@}��Z%;7ѳ�5��"���54*��C�x�jJC�^^6�QI6!�-6�۵28�5�6 �4<�N�*"N6�tK6���+�������V5�|�6�8�/�(6:2�6m���v���ȶ���6x|��𝊶�5/�p��4�!7����9�69����L�M�u6��59��D!�qS=5 '�����l�5J�ϵ0��5��6>�>���6���5r5���/5S�ŵ���&��a
�HWɵ j)6EAl3��2��9�6s�׶��o�@	�6���5�'�jiw�s5����6�hH6P��`v�*�X6�+���hʶ�j�6�ή6���5N*6'6!����5Ya��������61��6�?�5��6q�"�h6����@s5�*5�.q6��4��6_�r��Լ��|N4���6�3�6l�6��t6��\�7#6�M�6���6:#�4�',5�1�52�� �r44X�6aC-5��5�~�6,��� ��3:W6 ;���~�����5�=�5�|�6�64��5 _��ѐ0�E�V��m+�V�5��׵c����4�5�/6w�6�5�J@5b��vqζ���F�6��5B>6[{�6�W�����Rq�6Fе�7��60_����pc6F:6�����6~�W��t�5�5X���ʶ6�җ5�T5����
7���5�tF5�G5��5��16�b5������1�d��5jW ���O6�{@52�\��f��� [�'�b�W6�-u6��Q6���c����%�'��6�����5�v16b�E68�48�6�W�����5K��4z7W6,��6���#G6$�\�bpB5x}�5�26&�¶�\�5 t�2���5 �t6����B�ҵ��4�r����6T�H6�]`��P585ۋ
5"�õ� ��7D6:u�����~�t5�[�3�5�d�/����������6}��������6����4T��6P������5B��5
��5����<'6�۵2\� `6���Pn��"��>���Ao�6�4����3��S7�9v�pqo6�P�5m���P钴[���:�6]˵���50���6Af�8���1h��t7���.�4	��*iO5f��[qƶ�C6���6���6$��X��5X�/6 �5�b��G�*��9�6\��@�5_,K��Sy���4�������5�o 7�)�|�#����5�
�6����ݵ=T�G��V³5�����:�6t�����%!����6
C<78N60o6@옶SZ�5(��FP�5&6]��6���6O6�d3�n�����5����EUV7�6���)A5�5݄6�<�5B�򵠤���U�6T8��P�6�E���7�5z�����6�/"�R	 7qX��H��赱R�5��Z7����w���X��f��|G-�����R6#�6�OŲ��c��U6���4Z>�68c�68��6�����z]6X��c��~�^6�6"g�6�G���M�5��B6g�7�0��.76��f5Z����P��5��6� {6b)���s665��86������������-i����6��C6�;���J^6(f�BЃ��S�5�>����5:�ܵ4s ��2��[�u��$Q5Ź ��p���T�5|֬�.�6�r6ֽ{���*��-���P�6r�J6v����6 �18�5�o��;�,k�l��6X���mt6�nJ6����z��������ⶏ�7O06I�_�H��5��H�x�4�56%������'6�VC�D����t6μöͻb5�M73b����ٚ�l��5��*6'1�7zS�+}}�)ܵXi�5xMs��5��0��=�6l�G��0�6��@���۲��"6A��56d*74$�%�y6(;y6�C6���6<ļ5�_ �A���F#���^_6���b!���:�6&�54�f����6lђ4�ag6�� ���̵���d�G����6 �1�b��r��6;�ö���5��86j��U�[6�B5��4�p���F�F{9�s!�5~��5���HF�6�3�4 k"5�����Q�y����t6��5h�6���6 :Y�\N��σ6|��4(�ҵ������6��V�b�5v(�6�i��&|6'����Za�6_誵�|�����Pzp6� �5+�����J\�6}�6O�Ѷ${50Ҵ�����Rr0���d�b7��A6�%�6�����P�6y�6p;�4��4M�n��q6��0�/�46� ��e-��o��P645h�H6/6M�ᵱ|�6P�0�cS-�jKն��6�/5���`�`�?L¶9$��瞵�X6����2��5j�̶{G��h��Q�6)��J�2��1��,5x<�5(=��I�6`��4�΢��#6m%������)���x5�r?��y�5�Y���}R�Y��6�.�5�5 {!��<���Cs5r 6���5P��4_g.�<�5L�۵��3(9	5�C�����=�ȵ��*�	!6�F�6(�l�����xO6�d�4�آ5劝�v�6��u5�p[����u�6u���v�5f 6�)6��5dd_���6˔���~��5���J#d6x��jj+���5��j��ٮ6a�6֮�6W7c6P�"6J5�z4h�%U�fӨ���/�,����>"����ˀ�c�~��V뵠��4<�3��$� _�3���??�6ă��B���t{����E4�:\�Mr�lM�5 ��5��c5Ȇ|�%9�C$7X���kX�U����6 ������(�q6�ɟ��)6�V�5��ɵo��t��Ryv��Wq5�v5]��v����W�6�ӵz0�5-�K�=�|6� �� rb6�[6Az,�b��5��0���޵�$h��HK�����ھ5~	�qz���fص�����nʅ6f�i6Ի&�R$��m�S�hdI6]=�r���*�5�;�4x��.�.��+��p�ȶ�M�5�C6��5|[6*�P�Ha�4�-5l ���T55�i6������8��/6Ǎ�5������v��8��/D�@��&����RP6��̵�+�����2Շ��,���U� �Գ �Ӵ0��|����K����x�M\2����J�5�Ŗ6�엶��5
Ȃ6ۣh66�ײ4��е��?��oM6�5x���x�:6�x5�`���8X�l��5�Xö_)�5�y�PA�N�5빏������6p����5���4����qG6dN6^ ���穵��N�8w42$1��:��+�6<'6�y���9��.��H��5 .�5��T4��D�ȉ�5��5b#���f��V(6�<:6�?�I�*6�{�5�<�c�k6X������3�ԏ5��k�\d����+5�5Ұ]�e	6p<�p&6n!���6 ߇�LrG��|,6L)5�6T���5^b�5�+�av��
�E6�562�ȵ�i�_	2�Ɇ˵���5�6�5�'5��_�%��60x��00���6�j��O�ȴҽ��ݔ3`V6������X�4��X6��}�p��5\�|6��W�pj40��>�������_v�D�6��E4�7'�
V;��!5�"��,9�p�6�k��Nߵ(?o5�)6��6���4��W6�z�5�OK647�5~>�6���n����5�u4�k&5N;���aX�bk�5�M�O�6p}�50n6�Q5L���>Q�4W96�Y�����5�GW6��Ӵ~t�5�%1�퓓�h��6�*d6�G�R.��6~�5���΍6��L��4�,nQ�r��Gnk6�e�L6Z\q�xA9��'�5ז1�n@	���,5l��4�o��`���4���Փ6��V���9��വ�`����ȵ�@��W�5"��5^"�v���7��x>�n�064���6��
6�̳��25ӵ�f<�t�(�`ܸ5PV�D��4˙�5"��5�n��aqϵ���5�9���>l5\���ݴ��N���?�6gi�.@5����.��5L�%5ʘ�5��g6fK(���5#���n�}��"����Ŵ�a5@�p��%̵�%6dr$�F�<L�5@����\�p��6�C6 V����K-�v�5@���D!�텨5�ބ5Q7�w�5�%���sڶ��
�(^6NmJ��CN6*2���5���6����#����<���6r� 6Hj�ȵl� 
Q5R�H6�tJ6"~�HD6[6��6��6�005l�6 k�4��4X�6���d6
6���p^6���tϫ�%Ƈ6�%�3��t5_�����W�y�6?2.��;ٵ j����6�@�6��w5ˁϵ.OZ�jWF���W�kU.��^�6�76Y�c��ҵ�h�k�46��:6.58(4����48��`6x��
��5X������5>E��C���6n���ꪵ��60G�43Q6pj6eS���6��do 6�Զ5��5h�����f6�� 6h6��Ď6����";�6?6�.6>��6��4��k��6�p�5nh�5��]��52Ɏ�`��6B~���R5��5���4�k�=�6�ެ�M���q��j,��bw����n},6 �6����N5��0��5o�/�с7V��h�6V��6w.�5�d�%�����õR��5Fj>7n.��wȵ���5����V"���'���l��;5;9�Ȱ�6ε��!6���5�3�58-�&�6˦�6dfY5�� 4�o����+���S����h��6Ξ*7��Ķ�r68?V���6 ���Z��5�v�4�N����5K�`�r�ɵ�x�%�ӌ6z����q6u�y��6�45��αHU<5����]T��p�6���6i��%�6��>͉�x���]���̶�2�4(��B�����J5�/5���v�Q�:6�B�5x �dY��l6L�J�25�s󵎜b5�T%�&��6P����4��^Ě��A;����R���I��ţ6n���;,����t���
�.I�6Ԫ(6�vN5�����T�5`����4���3��G6W�6pb4�eֶ�ڜ�H�L���6��絓ß�i�6���Šo6bI���-:5t�e��ƫ�:�'��۶����836 F��ir5Ү6ľζ�,5b< 6VW5<7��m|5 �޳��ж�I������l��Z�6-m���D�46�\�5�'!6v��5dYq6R����A���Y�50//�Ɏ��]$��\E6���6�k5��C5�fF6 9t��؀6\|�j;Ӷۙ�I�4�y�5�(�6J;���["���g06���6 ̞�x^�6H�6�0����-���z5-Za6��6O�26��̵�46,�߶$��6��i5��6���6�Ʊ6(St6�T1�6.6�P�b[!6P�5���6q{b7����@��4ʡ�5� |�S��6��?(6�!4�`Յ5 �����Ӵ���6�7v����6�w���5Ԑ�\[��)ˤ5��"� K�6`z5��b���5� ;6�ʗ��
7��8^6�!a���:5�����R�3�|�6���64��4�CH6@Q=�.�w6M9ж���5"�6��^6vt#6=�e6��Q�ݘ�6�T�56�5���tO���5��{����6���6���?36p�쵗� 6@��3�2��4:6������o5�	����"�/����>�6�?��ا6�j���؊��u�5���5�6�ƻ66#��<��6p�ֵ�T�6�^I6���5^��6?$�:��5�76�Y�6,�ϴ�eض�H76���43F��m!����6Lz�6ж�h6���6���M�c��	¶�_���s�6���p�@D��i��5�y*6D��6ft����	��6l�"6晡6�q˶ �u�$�n3�5�&a�c�6|���}��k5��µjf�6Bc56���6��]�(����aj���7p:6 y�6iĘ6�Pq����\�L4������5@a=6cJ�5�*�6�xX6<�'7���8�S5n��5]c6��E6�i����׵ܗ�4+
��i�6ޞ6&�5��R5�}6.ž6�M�6o�X�pJ1���3���6�̲4��6�0�4�m�6�.B7��˵��6��6��56x�a��(�5�=��",�����U��Zs37��p6���6_��6�5�
�5�}���aR6^��6�~l��54�^����b�q��6|T�6ح7��6�#�6<6��7�I�6Rd}�<�6E�)7��r3�z�����jՑ����7ѭ���?7㋞�J�|5��	7���8h���;7����5�Ӷ�26P��6��F6K�Ķ0X�� �W5dZ����5"\����=6�`��m06�����5���&�3�5�Y6$v?�����&�#�*B�48�6&�5|U-��L�5D��4��c69���D\�����<7�%�������E4Η��p�\�A:��t�4��d��k�����<�{6��5��6��q��춱qU��zٶ|tM���5>��6d "�T���}���伉���p�T���%�Ԩ�4��j�6𬦵6%7�H>6���;�#��ε��e��O6X��44n6��5�x�	0ӵ���6�U?�/�@���@g|5�9�6�0+6���5hb\�'�	6��U6�#������赭F=��n7�c��Ŧ5t����x��G�6��S6���XN41ն�Ω6*�.�D�0� )e��y�6��j�Զ?�����6|��5�:�� ���9���|-4�����BѶ�6,�46&��ќ6t���G��1�6 ��6�������Y5��<��]�6	�7�y[��67�C�5�ᶬ�-68ԙ�~X�"Џ6D6�5[��u 6��06i�<�ض��<�16���pv_��g>�����͌���6ն�5@f�5Z���i��5�ᶋ#����P�����b5Q�����x�J ����4-�g�`���S56��H�~��6�B����@4�V�Q<s�����^�&�TyQ�R���7ڨ�6���5^��6�qu����T�5�(8�����ƌ�t����zl�pb�Fۚ52�jSx6���2�����5v/�WX�6���I6�Pa���f�4#��P'�4(7&����5��5
^7�n�6˩�5Ж�5���5_�6B����\e5}��,ׄ�y�6�5���5ы5�
t6�o�t�5��<���������1��Ԟ��;��5�w�4�y6^�b�hߊ4�D6���n�̶����i&�6r�ܵM_۵�ꕶ�n��0�6H�c������������ކ�2�K���6$sҶ��#6�0@���561yƴ�rе�ϵ�ֹ�fG��8{_��L26bT6�16�����o5�ҍ�k�ٵkU���Uȵ�2�5����ߵ15U^�K.%��6F���Tϵ��5�JP���}6�]D4�说*�75��2��/�5�X6,t��p(�4p�O����5E'��b��5P���)7!$t6���D�>6��G6��������Y5�?�3m�6a806#:����6Pw�R���\n6r�Ե8�� �W����3���6Ps�5a�<6�%s���5�R����5��Y�5�1��p@̶H�3���5aZh6[a6P5�}�5��h���<\�6z���m��6{�6�?�����4���4�6�$��Lq7���ǭ���5�d޴��5X��+�5W.6"/��,�6&5�5�!�4j]6�Z�5N���c6\[�5+� ���5�­5�o9�lLŵ���^�26~3�6�>��[�����6��6���?��5 ;^4P^5���\o6�*���A6Ha�5�k�����6I$���6ؖ�z���c��A^%6T6�W���̶��6op�6<f#5�ә6I�r6�ք6�W¶ׯ��Wj-6�E�'K�6o
ҵ1˵�_!�<�5A"�5zR5���97�6d�6B���S��5�$ 5�_k6�&�6�R@�^n�5�mO�I�0�z������`�R�w��^]�d1�������6,�S5c��u��5L��5�T���0�5R6��`����6�զ�)#µA˴$��4`!3��53^��:v�4� *����4pH5�DI� �22f�46�[��eY�ᒵ�%�5 4�0:�V5�UY�r!�&k�4�Q�Lg�4�+�5pQ�5��5�@X���n�^6�Sz6㨵�ܲ㵢!��PV�4>5v���Su��>����m���6�xy�f<N��j�5Ү�5�^A6�|�5�|6�0���6��V��4���6�K��M�5q�6��5]��5���U�P6��
����6�{t6�����g6(w�5�Hs���F6U˓��2�5��Z5I��5|��G�e6�Ah6�\5�D7��
~4��5�6�8�4��:����5tD5�B�õ~⡶�6x5�5�U5��9��-��d�4�p,����%�4��h�d/#��Л5 �5(gQ� ͇4L��pk�5�xZ4r�b���$9����״ �i4Z�5895H��Rx6�m��@8�X�5�@��g ��AB6z��k46�f�5
����[�5�s<5hK74(fu4<K?63�.6� 6}66d�J6��[6^�`�/5�M�
��5>ĵ��J��5��5��t6�6U}յ���6_�����5���5 lǱ��õ�r5�v��P=�Q]5<�P�`h�3���{�5pd��n'��s6�b?5�5P4�Q6�x�8��c� P���e5������xh5H�$��ǵ�]6�]�50R[6�a+��a.�,P�6�Ϝ5��?�@+Ӳv�5h�=��66yIg6{����a5���5
�&�>��޻�m<n6��6�V��1y�h�5Y/��\���p�@�t85$P�4�4�ä���ӵ�ۼ5�G��q]굠��8��4��Z������6�5�哶I6�w.5��4J>y6���u�fO&6=��5�b�By����d��4| &�����e�3���6}!5\���3�4��崚�p�^5~�4�ę����5�G��������4��o�:���5J��5@|3��4�V ����邵��5�O�3`kW�L��3r�6����A�6�;86�玵/�5�K�5_�m5�>����>i�5#���|��э5!k�6��7P�Xm53�M6Vi6���5��6���4���5?��x�ֵ�.�T�´;5a�5T$P6�%�"M6K�����6����$6X 5��5���5 ��5����4L"�W6G6RG�[�5�G�5T��4C�ִ��5?ܲ�=-�R,�5�ݛ5pv�3��׳��5�ϵ{`��<>��}��wx+6nn45"<�W�5�ݵ�75����4J���%�6�砵�\N5�4�!��d�6c��ˋ��#�36u�6��<Gu3p�'���5z��Ոg6��j��@���{65S튴��4���5S��6�%4 3L��2
��Y�4B��4�Ln�N��5L�����5�S�t8�5���5з]�6i�5��֚��8�S�`��4@2����2,r��Br����5���5	�>�I�O6���6����j`�*ݺ53��5~�9�ʱ�T��5�_�2��/48|4��Ze��% 6� ���R65��4�{+���-6����4��X���UD2�w�6�]q�xځ���5�68U�4�j�5��6�j�z��5 ?��GH�5��õAtŵj0�5b!�5��%mٵ)���O5u�]5`��@5�C�5P��4�c�5�4D�h5ج5��6��ƨ5�6+�6�o�<|����ʵ�&�45�ͭ5!��5������5�V6{m-69�a�5LE�4_5gc'��:���=�������@���6A	�6
���y�5����,{5�Vk6��?�X�63��&�@�5Z[�����"�5R{(���6�6��*��{6	����x58e��Y�������S&6��E5��6(5���;4nm6�b��9*6h+���J6���5��pD�5���40�س|q�����4��4�1��q��O�k6�0���X�V'4m5�c@5"3<�y�C5����6�R � E+���S6Ƞz��^t�ĵ@6�Y��ȴ̴��V���4�4�$fj�|�6��� e�3脪5�a�H�� +�5����P��4DO��˕4ضo�jF]����3*�+6C�+6@$��25��w��״��[4�������5P,^��=6�>�k���]#6"�4ﭵਜ਼5��Ķ�W�5�岵���6��/�:	�5� ��,��50π4[=w��[�5r��80��Z&5|n��f��6.tI6 �\5 �:4��#�y�5� ��̧ϵ{�`6"+�6�]p�B����k��[6����gr����\'���G�6���lG6�Pw4�mj�I��[���Y���:T@6ѡg5��5��4�f`�`A4��P6S��|���S�6*��6y�:��L�{c�5������b���d5�D6�����$6^�4���~5��5Ϛq6������6/�C6�֎���?6��-6 "��i�5�g��̣\��u#6���5���PzI4[�K��a�5}�H���r��6<�'�����TV6��.�o6l3��@�4���6Ӣ�W�r60U�2�=4�u�6F�1���_�h�5T0C���e5���XZ���T��u !�+o�6�!���Q=�nȦ6��)���G3*�\6�B68�&��#J��|��|�-6��B��`�6��Ƕ#+�6s�=�4�4@N���6��v�G�T�Ӗ1���6��v��^��[�65\���[61Ұ�X�I5@z`6DpI�.�qZp60�n5�5�q������6�[q6�y͵�6]I�5 ��q���<A6p3�4�^�6o��ܷ\6�M�6F��6�ȯ4@U�3P�5 �Ǵ�Bw6�\7ĐU6�*�	��5�d�5l��Kn�6_*�8��s��636��$6%F�6�Ǐ5���� �6�
P�h��4xdb���58�X��ٶ�h)6Kā6���5h�/�e���ٵ��N�
��6Õ5����H��6�����% 7
.x�k<�m"268�z�d� ��2X3���=���6b���<ߢ6b>�5sk+�t�6L��4����z�6f�5�6-�
\ƶ�`6�7���3�c ����6f8�6�=n���6�K��9�61�l������϶!�ʶ��5#�6Xg6;�(7z%%��-��7�7tI��[�ZW�6�8�5�Tд��6Tvr��p79m��
A6_v��?4rT7"����ɴ��[5n��5k���ҳ|�HA�6�/6����e4�һ5�Y���T6�6@#�������6X3�6��1��Un4�1�6�É6,�E6͔q��<�on+65�	6>F{��o 7R��6L�56����Ǔ��aH6�c�6�X7Q���T�P5_�ᵟ~ֶ�𒵐�\�8�O�T��6RfE6�Ak�B��6�=���P�6��� ���܃�+ٖ�3c�5 �����U6ih���O�P�R4&{˶�kA�L��5�5Q����T	X6�Jĵ�r���O��{X6j䵵�A��מ��a@��6�|-6���5�e�6Bk�5�W~5�Ju���q�	sA6�O���"����u�6̒R� �ҳ#�6��9��E��6!�6�R��񸔶�������5`K�����3�+�6v���?�6�X�5�+µ:ʢ6��=�3�7x�_�j�x�h��6�!`�8cL��Xe��u��p'K��3�5��1+��#6������`�-5���5P�@6C����sr4��6����,��6�0�{Q6(㪶�m���ҵ��7�7l�Ͷ]�65�^�Tw�5�յK�d��9Ѷ�5$�77��:�	aƵ�6�Ն��m[��)�[��5F쇶�h�6�:�����;[��'�5��:6xGt51/�6��<;�6m$F6��6�@%5öt+�Џk��pݶTB��x6�R35X�6$�R����6A;��ٍ�5�}u�9�6��5 �1�(�x�S?54G&�C���=�5���� ��G�\��O�����a[Ƶ��Z���6��/��%�/�6��Z�Ƙ�5��<6d����8��N�?���\5�#ᵤ����ꪵܱ�5����B	6���*���`7F��<sӴ
yq6�j�v��6��"�ZH�^�ֵ`m|�5��F��5)^I��}6W���`�
7~�4����=�֐�4�A6j@��~c���nIL6�M�5����,eS5'�R���5GQ6K6	��@�޶��=�2庶<=����趜d�5��ô0�5r�l6F��6��϶�(�4�g�/��5��5�����:���6!7�YZ��#�5��_6xV�Pv(���4?����ڵ��y6�O���� 6B�*5���5�O�6��4ڋ�5�6�5
�&6T䴶��J6�y���5�7��gq��5*b_6L���j>�]��5����􈶳}6G>~6D�?4�nе���6�7L5�Hk�� 4�2"6���5��(���86������=6����pȋ4(�5^��5�Dl�X�ٶ4}6���50[���9�6��6� ��w��p�S7b\}���l6�C5?�6����4�^��o�6w�6��̶o������5fw��H/6��T6���5@���ۍ�5v���A#��c�4�g6������s�:��
Z�6��Q��ǉ��o6b����z�����8��4��8������!6{ڒ5�Y�F��3��5�B���X�5J�5(�6������5���چ��I�Ģ+���7 Ð�*n6<��6%\�6��մ��5��6W�P�(�V6���a䶐��`�K5(e6��6N�6������,4���5�=���h5���5�`εj����g�(6b5��6ո$�!]���
�&΋6��Գ�^H��ൾ���ƶ6��6^!R6��j5،�������r�5�� ��Uݶ��P�n��@��� 
�t�L6l�4M5 ~����5�`L6��5�C�g�5D��5�X�5s��5�K4�.�6#���������5G%��6�6�����}6�(83�6~��R7��61�7��+�M���˶ f�4��6�[5�5{��+������Z�ʶ��`$
6�N�5��ݶR�ﶜK�6r��6Z=
�8�ʶ���6B��࠻5`�86�	ӵ�j�ʠ����NM��Ƶ6�A7e���q��&ƶv��6���.E�6�^ڵʲ57�v6 �4�:�Xs����6�y]�XP����յ8*6�϶m�	��U7�׸����6���-�5	�6)�7vq�6 ���}	6��#��tմ ��3�o6�jl6��6"�5��$�6Q�}�����i5?�3�O��5��7{V06Z`�64����� ��{�6���]ԁ�� ��@l�6l��5�Q��w"3��76���68Eֶ��"5i���(�5��ʶ�'�6���6{Oݶ��6H�W�d-7��]�P�5�?7EQ�+�6P����(7&�X��a�6�:F6Ȇ��ȉ5S��6�ޣ��l6HN��<�4�׏3K��6T?6���4#�6���p<6C�6��5��4a_�� ����P�G��6�R6���0�ȶ�C�E-�6"=z6j�6p��DP66͆5@내�x�4�1U�X�a�:d7rܻ5
r���d��L��#!���e�M�6��o6"�l6�U�608��a�0�k���27���6�3̶�ƺ��6������^�>9�6h���o��6��M�<'_6�915 :#7	�7�ua6 3h�������6�Kc��5�6�ƶ����7pI>��-{���B6��5B�7(_��WO6WX���)ǵHO�5���6t�5pSO��46��d�G�5�iY65���@)6�� 5���4��6`8�6���5=͵@������R�H7-6����n7��0����q���5lm#�e�ٶ��,�ɺ�6�
����6@UG4D�,�=S����t�1�G&7#��.��o��j37<|�6�R6Ú7��5���ƶ<�5�?1��ǟ6\:'�����L�$7,�@��Q3��$��5a�4�E&6�C���I�6���*��)v4�36E�96�4���4�n�5�58*#5�%�54Ũ5����w��r��{�5���5�FC5�*6�玶2�Z5�I
6���5�`P6��X�e����J��K�26>5�
Z6�����63;.�W�,60�z��Fh505$��5�*�5@uM�`"7 ��P�5P�Z6D45��6x����S6�s�5�T{�?�6H`��q��6�y]6�����������5��۵����{6`��d���>5�W�5ʡv��}�6�B�PX�4k���hCW��� �*���8�6�(������Գ4��5��
��)54���M�6�7��C^%��f6;��5V�|�Ă��r5�6H��^	�6N�� �i��i 6�t�6�(�5Ty��מ6���F'�x+4��6�ŉ����4�\+����5�_\5�敶9p�5 ��5�tN�@1i5��ص�)6T|r���G��<���ɂ�r�6{�K����5d��5��O�E���;��T�d��I��0+�3z@��k�5Li��@��8*6rN �^��5 �94�$�6��6j�;���B6��6r�����r��6��=5Ћ��f��
W�QE�As��t5I��5���i��&V6���6h�5s�õ 2;4pA�5���t�4Cµu1��,W5�GP6��L����5q�󵞡��=vŶ��J���6�y5�����0�2��4r~#6rFb6:?���B�wP�6D��5Iy-6ǻ5�撶$�5c7#�6�1u5��I6G��j��Ƕ����4W�]�xŶ�F���#6u��6��ߵ�v7A�����4�?��M6Ep��z�5&jO�8��Vb�6��F6�t�6x�/��/h5cs6��n�������bV�VU�6�A�b	f�hF����6���GX涜�}6���2a�]6PR+5ha5���62li6&�6 �W3nͫ6�h�=M�6��6(����4%�m���5`n`���e�V��@�5Ԭ~6JU�5��{6�7��TF25����,)�6��;6����27�����+6/s6�l6�])6���6s��5Q�6C����췵`//��6���5j���z���EͶ��6�Z�5v0M�,�v6 �汕�۶�D6r�+6o����6�d6�^��A�5"��6?���m�7�{4��5r)���k5��t6'�6��	�[86ˑ5j�A�0�`4+�6Ȇ,�t���69��L�46ㇵ��6��6 n��,������ؠ���<�4v��t��$�5��L�l���d涠5M�5Ȓ����5�d�5za�5*
66����^�d�Զ^��6�m�����5謶� C	3�q���m�5C71�:ߵ�nk��K���6�����`�50.�2(R�T@��[r��{�Ԫb��$�6L���*�L����t���*�����B�E,�����@�y4�~*��A˵�f�ZÈ6 q4��9��8f���ҫ6�u���5��06U�26�9�5�dQ�Z�5qx�5�n��n������t 6*��6���8��5�7�UN�]�$5H�c���6��c�5ph�5b��5O����|5����������6|o�5է��o������a튵��6�ב5l�5ާ�lC/5��{еPh��X��ዶ�����*صpǾ���@F���%6��6yp�ȓ5R:�6�I�7g�6�X�4���������6�쫵$֖5���6�^��YZ
7��5xP�p a43)ҶDG'��a6H��6����V6_��6��e5{���T$��c�65sC�(׻�ʛ�;ᰶ	�� (�5'1_6��6LzF�F]�5$���Jz��W�������������R����5=y6b�-�&9�tr[6s�5� 61����Ҷe�6��t6 m�2�)�5N���Z�p��Ft���b6h�ϴ���Ŗ�6�:�����MնR����>|�x��5��Ķ���t~x��f��^c�5@��3
�H6C�l�	⾶J���Z�6� ��Pt8�9��4_���̴��6`0��~"5�S�F6Mw$�ˋ6L\p��1�,����c�6h�-5X���W�6 r=3�"�3ٿ�5��50�"�5����,^�4�"�5���4-�5�J�R��"P5􈽴���4�>u���`��䋵؀�4R��5�h��?�6��5�F���A5r#06Js�5`�z5��5GĶX��5��_6 ���R\��5v���R�6e�4,T��X��5�Ì� �#����5��4NX���u76 hs�ĕ���.6�+��H7��4�fI�z�P��!�N(�5���5P�6�R�5�p2� ��5��ִ��5`WX3�}6�i���.6B���gp�L�}5�D�K�6  �r�V5��B�Z�ĵ���C�*�r��\5�OO��O������P!�@D���5@P�5��w��b�����Eb��պ5�
f��I�QF	6�7F64��0�5���5пP6"�5��i�5�|K��n�R�6X�4�'6��J5�촹��5R$�5DA�5z�5h#�4h]�4L]
6�%����
6��:���M4�y5b�!���D�\�5�(63���@�5h�,5 ��jTg6 ���A��rp:���<�X\<���>5`+���4 @��f��4��6�߻5�Ƽ�K6�-g��GI5�J�&�]�Ϋ�5��5 mW� B�3<�Q��@��N��ֽ�5#�� �9���75���5��U6��5��5�2� ��4����N��H��5hV�\{��!5�`S�RSu�j��5J�6�zZ6�W���j�|��5�����%�`κ4�TZ�؅�4��'6r�6�f��:"�6ب	6���4�+ 6>u�~����4�}b���6�[�6������_64m5��4<�x����5�Z�5�7��Q�J5�ؔ4���4�^5}36�m6�W���ٛ�w��@2F6|�ٵ*���q�
6zյF6�m������ 4�6��6/�H������6�f�5��;��?�5^v�5v\5a =��<=5/�O6�H5��ࢶ������7�2By5	���� 6�Ĵ>r6x��}�	6�د����5��>��$5��Y5�6�p�5T��� 5x�}����5�n��8���S���@�5B�w�6k)6@���λ4,��3㽰5W�96�J6��?5�7�4nT���P ��M�5������)6�Ԙ���5�<]6�s70��3��5�5���E%����X�j���ϵG��6�;t6:���5^�4�lʹ��6^�@�I��6����Bߢ�H_ݶ�ۿ3��մp�6I4�O9��t�߻ �0�4���5�(:�)6>�L
���B��#(��SK5h��5��5�������D�+G�5 ��5���5@��4�ٳVpu6�5Z���6�R�5�z��w�����e_6=�6�u���85��4��� ��6�+�0�"4����4o�.��5��c5G!�g�ϵZZ�5R�R6�2�5H��4ň^5f���> ĵpf#6����,+ӵQ����g�����5�R�%��4{�5��$6J�#� F�1��5櫿5P���,%��*��-15�����5��)5w�w����X�6��5ø5 +�7(s6��)��x?�{��]'�����F6�7��x�r�/��t�4p�6�X�ְ��P6�(]6��4��ݵ}!�4�b��1�5���+��Z�2M�Q6�;��(yƴ�\T5"r6b6J�˵�G���5|��58�L�E�V5�\�4ǘ5�Y`�Պ65X����6<4
4}�O6�f5+���nB�5��3�d�5җ�4-�O���&���H5R*(�sf����l��J�4��&6	 6�r�5t�55���6�N�4�c%�g@�6���5�4�õ������#�ț�,�&�T1�4���PG�6�5���)�6 @?�fي���6=L���44ڵa6>1��X�436����34w���@�76Y��6�8��Q6@6�֦���L�����k`�6T��6�q��i�7R+���C6/�5���-(�6�E^6Mq�����52�Y�J6�µ#��6��5,_ݴ�)z�ʸ���?�5Α���M�4=��5����L�5�����x�6�>7Lj��Nl��_�J�6�ζ�U�6�P�6��S6'����`��LR���J�6RY"���:��6t�̵Z���)�6��E�q�����:�U�6�n���s�6W�ĵ�a�6�X�3:x�6j�����ȴu\�S��6<�������ѵ��D6�,N5���5jn޵p��5x��������
/����5��X�>�!6�ڵ�(����6N'�6��(�  ���=5��_5��*)���B4l�D�,8v� Ɯ6X}-���/�ȫĵg15��n5�0ŵ����n�Zpc�_|��g�H�,P60�5B��5 �ٲ�&66���5R�6Hѵ�X�4jQp����6����k����6:i̵�\S6���`Z�3�66'ԶÚ5�>J5ꏈ6�D6��z�B�6]Y�Ϋi6#5�F���H�%�6D��5hk��(.���}ݶ�aZ6
�ʶ�����ӊ�6�'6� z����4�R˵< ��������L�A6Ϫ;6hJ4���6o���m
6H6�6u���S������ж������o6jo��HŶ�
7|"k6���QP7&�w,]5S�7�C���赵�"7ȯ�L'6��4o쫵r��6:����><6J��6@\6�u���¶ |�2��i5��5�ڗ6���5�#��v���� ��F�4nv�(g/�	,=5\&���sݶb%�����4�|�c����5�#ӵv;�5��V6�$�4~/��ށ��7>���e6^�+�� @6t�Q6�K�5�`�6|9�5j��5��6N����˚6/�[6��?6^��5�0$��q6��˶���܁��G͵KQ$6���6�����6��)�nA6=�6@4���)5��6�����ո�L�A5�\���b�����3��.n5�
5�r�����6P��>l�5 h��ർ��5��N�u2�`+�3�z�5�6�������6G��6��6�����&�?j��,����\�I�'�T�ܶũ�^z�����C6BC6;A�ڼ�5�Ե��{���4b�	�vk�56���� �������W�6RU-���k���H6�Q��`W����62W��[�˶J"���6��5�6��� ^7���5����䥶����a��>�a����6�Ř4�C�5�.����6BGD6�7�f��5��۶j �6t,L��6�a�Ɛ ���@��ه6��$�{�W6̺6M�!���;4�F����ᵖ`��#;�2�q�`6͙��|7
��6tq�6,�5e*�����Gr� ��5zb�������e5��5�%p��6��v5�Զ�w۵Jǒ�fs6[�µԠ�4[ʈ6 ��2��q5;�5���6|�ǳ�,z�
�B�kLC�$�5 '�h{6�ᡶ��/�W����26h�����c4���y��7vɵho*5�L�?��۩6��P��4a�P5�/7�|�I ��"�6���5�1��h�s��)6ź��x����L7qB6�6�AA4쮸4Ҭ ���69�/��5����@�=��[_�؄崊0�6�o�5Ѣ�6�+f�(v�6 0�4h=�6ұ�ED��@�E�@�5�Ŋ6��f �����=6@I<5t��5���5 ��3k</�D��@��̔����4��(5����{;�5h��7J&��A���v�X�D��ζ� 2�4�y���(s�p@鴿(��nC��n�5�׍���6F	��w��L ���0��蹶M�^��;�5�O6�P�� ��5H�5� ���z 50;]�Ք�5��>����.4o5u�N�17�����6m?66.�3�ö`�47�Y5����1�5�?ֶ'���a�6RAD6YgG��G�x,Z�0<�������S<���w64R��=���Aҵ�6]V�J��5@�25�/��LA;5l�u�.�Ƶ4j��G6���5D�5�g���P����� �t	<5f]M7�E�6�c �/#����$�¶{Ib�G��6�G̶��I��F-6D����6
6	�P65��6�6Vc�\T6 ����o6�PA���A����5o�A���5���5��6z���E:�� ���+6�@6���6�ԛ�覬5����>�60q�5ñ�5��@6��j6�tL�@G׵[7�6FѰ6�q`���4�+�� ��9�6X'���4vr��PN���]6*��6�A�&C�6��E5dn��'�6\��6�M�����$��6���4��5�̏��;�6�95�7%����6�i'6۫!�P��
vv�"�6�,{�6���6�Go6;�r�LwڵnJ64�6���6���6���5^���]P6�̶����7-�7�[6��)��t5hC�d�x6��46Bմ�F6��p+I��?6�ȇ6	�5�&"��"ֶK�5���6j�&�:v����6/3�6%\5�6�o�Y��6�:���v)6��7�7Ͷ�C���6Fo��F+{6ćж�k�5���6�S��Z"�~o����6�	4��=��O5WD�6��6�Kʴ�5�6���5�@�6C�Ӷ2� �酂�����|%�i��6 23B�Z�H�6�D(6ɇx�yq6y�E�_w��0��6-�����5P_᳔�,��L5�2:�M���ƥ�6����@�4��6+0����'6�������D.5K���5�4�7��F~5;���[N��~�J�3\�6�0���6��յc�5�Tg5���6Z�ص 3'16� ^5�ۢ6 �T4�Զ��6����d�\�/6���:�6Ќ��0ɶ͞�6��6b.6�"0��Ƕ~������SF�63Y�6J���N7�$d���$6��=63����c6�86����0\�#�ݵ
6u��6Zuʵ�G�6��<��u�5���.1�F�6���5���5���6�����ĺ�4,$5�r4�µz\W���۴Rk7�A��` �4��z6�D���"|5|����h�����U6�Pd6+S��#�k�P��遶+��!�~�X6�	�bǆ��$>6��>5&��ヵ�µ6�6��>�p%5�$����6@]�6��L6a^L������5����T��5p�Q6ތK�i��d�7�Y�����6<��64R��������p6�&?�v�ƶ��������5H�8�P���4@�ĳPkԴ������69�~�������6�2	6�f�P"��=e$�$��5�$$��h84EY35@t��0J����.�,�fP�6树6��L6Z���2����d޵R;�6\��6T�>�t_V6P�96ժ���e��Z�j���b���E7>���ʐ6�Q쵾���e���'��ĵ���l5Ж6�6jF6�	����̶��6�W��)6�~o���d)�S#5�A�6j?5ƾ̶��5
 �63Z<6V�76X��I�0���T��u|�H�6*�84.005�de�H�5��!5�;�6��5EJR67�V6�6���6�i&�F#�4=����*�l��5ާ8�ym ���5~f6���4�U�5�J�6�L�5�?��E#�#7p�J5Nζ��A54�նCq7�l���㯵_<a6����s�5є �BG����6p�8����6��-����$^�5���6w_�� �@��4�+k��D�NB 6����խ�6�gB�b��5�dR��8���6����Et6� 2���6���< ^5^�6Џ� ర�%����Hjô,���򛌵W��6p�4v k60���1�3�4�@6�>�h� 5��6bft�l��6}9��y{�6@��4m$��&6�F6fy�6ꣶ47^6޾ζ��5�&j5��-���6V�4�u6�����e!�����t͠6b"�5�N�5�~ѶPmQ6�خ6�Q����6�>6H�E�ԙ0�=e�<�M6�����B��8�6 @յ�r���Y5��X��t�62����
�T�.7`�4��6�06x�d6�I�5@������4�������	o��?X60�������r��������>�h\7N������5 �@6aN�6�H2�ĵ��5�\e6���3��K�`���g�����5%�5� ��`)�6�޵�k����W6 .2�.dն/R�PcO�9��ދ6�C�6x�7�F3�LC�6��<��QN6RR���PR���R6㗵�1���U����5�D6���`5H&36����%1�xW� е�a��_�,���"�v�Ǵ�1#��J�Kur����8F�3���6�36��/�t����6���4d��4)6y��5�9�5f����5g.�5ܯ)�����۔�6oU�����f�4/��60��4D��6Wl��./��B�T6}-�����7+P&���6����\��<A�5�^a5�s�5�_x5K�]�dB5O-�5�?3�xk4�g6�4:6
��4a�6���f�����dA�D�*6t�.�]P0�Ą�5����<��,w��v�6<(35�� \�2u
дϿ�5P� 6Zs[6�����_��uW5��̵���3���5�h45�-5:�\5*W�5��ֶ�j�����5�L� U�|C5�7;6���6��>4�(�6�y�����6y=�����54!�5a���9�
��3�E�4v�$���L6�L6�a`��*�5�~S�
�ϴk4�6�77��65-�6Ն�5��y5��\�+6�bM4��m6 ���z�6��-6��50���Ȱ���05D5���6�|����4�E�4���7�6Ѐ �@Ew�]%��:`4�'4P4�6��е�÷5P��4 :5�P6����G�5N�K6�:�4<�ɵ`̮� �豯a�4�)��8Z5��Z��Q�5��N�DƇ���v6�6��5X�6���K��6��5qB���6t�r�`�ҵ�R65P޵�$6��)6H��H�4IYW6��j6q�6�*7hx�5���6��+5�� �N\���h��ˁ�6X�ĵ���6j���y�ݼ�6ٰ5v��5�ګ��p�����٩6N�6j4�x)�����X��4�p6 =5�!i���3Ғ�\8ɵ$����5�o�5�w�6<���0�S�8�P��76�A����6T�^��YA�Hk'6"󆵒-/�-��5��4,�6MV�5�^�K���ѹ������/���,��S��]�6��aG�6Lݥ��nk6PN6�}�5֏�A�!��R~�+�6A�6;x����$ځ�L��5��7���I���7����:U$�.BжQ	����5��6v2�6�/>��ֱ�@LӴ!�6P��5�L�6saٵ$6��d���`5f:�5~NǶ�M6���6��L��� ����(�7�����P��&���w4`�]6��5䠥�Tj�6�(7%{����7��G�~Z��%�@�|3�r��R7��ٴ��6l�5\��p���n6U_7�M?v��Q�6��6)'O�pԶ�����J5�� ����(1���$6B~O�O��sU5#�k�:6H-���ĳƣ0�8���!���5
�6IH8����6O-�6&꺶@�F5E�*�O�F�(�
�%x6�����Ѷ�=�6"��6�wF6Z�4�252� ��:ֶ։v���F�H�	7�팶Ɩ��ε5+�M�f#��X�B5+|��8�3��a��7�6n�i6l����Ra���r��57�	�q�7��5���c��ζ 
4z	��76vA6���7Ϛ6���;��6���q��6qKw6x�X�n	46��W5�Mµz�%�*<�������6T$�5cH�6�Q�4�Y��5��d6��?�5q�h��f16F{�5�?�6�=�5z��5�	<6��_��i���V/6���R:5NQ�6�Eh�I6�6z�6���6*U?� h	3��61�6�6�5�3�6��48푶�o�6�V���F;6��#��5W�6��쵟�7(����D��Ґ4B4���[ƵDk�5 �#3��O6��7�����b�6jW�6`V�5@���4;��O���;�P,z683�6}��6T�6'��6�/��]-36�?:7�,��8�6�\��{2�6xL��n26�h7
�6�Q�6-B5������7�G��_�6�n��|�ᵤ��5�@6y5="7��r�4��^�76�6���b�6l����жfz6Q�6n�5x&|7vK�6�#��BA굪�ĵ�7���pD�6T�9�LlM�<�#64�g�f����6�1�,��6�寶 J�5�/7|�O�8?
�)R5e�a���M���7g�B��"���C��A�5-���7�������&����/���JW�6i�����5���̿յԥ�6b架�u#��:õ����y6J+����U���5�����<䶐C�5��s����?0�5n�}��t��c16���5�$=�@�ᵀy����6���6�Ͷ�r6�4����6�k6L��4��f6�f���6�Ü5-�O�9�|��f7�W!5�?�B�۵R��6*Ap��&�H{еyŅ5����6���6b��6=�P1:6����`4$H8���6@����6�`�6PG�5�ǅ�XW'���$6��ʴ� ���A�Fv� �,6�0����3����pҽ6�D�6�%����l61�7��6��h5)শ�A�pM���T7���5Z+��d�5.D��,���)}���6�Q�������-��FO���������V&�6������+��d{���3 )��g��6��bi6�+96�a6��6,Ř5T!���v����6V���*&v6# �6�`72�6�>��$[�4bTP6���58�6�]��/IZ6,�� 3��5��X�N5eg&6 \Z3� {���<5s��4b�5�m96�6C�H��6<{�����5�N�.��5z`ٵ�D�5N[�6���U�5�ß��i�66h\��m�5�z�5�#���I�T�48���䆍��R�3�k��և�6B�M��*�щ]6��6��:5Ғ:�@��4� �5�KF5^z�5��Θ^�]�6��P��B$6\��5�⫴ ��5bz��UP���4 @S��姵r�1�R�M6����>��-I6ۤ�4=8�nOH��hJ5�^5��̶vt6H?�j��.!��(�6�#F4PH6��a����jE�-�5P{-���6@S�4D$X�_M96�pU6�'6@֯3��5`�ٴd�3��m&�
��5`1�5Xd��
�5Z5��u5� ��/5��6�"ε�4汵��9�$�5P�'�Z�+�dJٵ�e���ĉ5��(5T۾�̦��r�3�����������5���5 浼5h=����1�>��M���s6P-��;M&6$�x��-&5N�$�p��4�4��1��\�86F7�5.��5G�6(tU4@�Ե��m��&�6Y+�@]�3��6�n?��6�sN�@��4d��4h'�H�65��fA�LL��I�5�3c�x��5�>��d6t�n6� 4�6L��61ڵh��r�5�?:�	�66��C��n�5(<E6NR6�š4��5/J�k`�5��Y5�8i�׺�5�X�� �#�z;6�J6t��4�E���N6<�I6��g�6 ��3ǐ06z>�5�� ��h������岚��5�(	�:�96���6��5�96JV1�d[�6�1��z0?6�Ì��#V�6��ٸ�5�XF����4N?u63~j��x�5�� �>yɵ���g� �X (��S��H���x%#��>Ƕ�dv4H�u�HӴ5�wе�fN6��K�^�5P �4ز85Ӽ�6���5~�,�׳�����������4�a26p|�O���Hy�6��6��66Q5�N�5&r �(صH�e5p�]�t	��YO�,uu������~�6P�Q5�[Y4�%5���3�NE6h�l�r �jŶ5@��>AO�id�Uv�l�#�6$�ҵ�{�6���`=M���56C�\!6�E�5���2�ћ5�*E52x6;��M�%6��>5�-�.,2�>M66#���&���:���� 6a�յ�+���0f5>cC�~1H���6��n6����6LKJ�\�;5�H�6�/C���Q6'�4xH~��OO6������ζv�36+�6F��6p�h�!by6�{u��t16@����Q�5�P3�d7��I��6ݚt6;�ⶲ,����#16C�6��r�`��L6Ue�6|v-4`��3Ϛ6�Q�<�H6��l�")���(�5�S��/*63�6 )�2Nq�5�l�� ����1ȶ`��H_ȴ.2�D�ö �74�$�UK7�G�5D)�6.�G���ɶ`J�4K�J�f�6�S$�yZ76Dq��V^�6眭5t�ٴ�[�5�M���ò7�6�����V�7R�v�:��6m�����z6����g�D۵�2��!��WLy5]�5��5v�ܶz[�6���4��x��B6��
Ϋ�U-36�]N5tI6N܉5��������5-헶�֜��<����6Z0Z5B�Ŵ��5ڑ�4d~06�zs��7~�Lx�H�������Q�5Q��a�:6=�6��^��V%6k�4|�Y6�5��A�v�6^�5��5�p�5Z�C6X����d�6�ڗ�B���ϵ��/6�vV�0�6K�q�Ņ���(6��5�_t6���5�s��A�H�.5_D5�͎��	�4���5W�36�nM��b��E����6Z�5<0D6Pve�� 6##5b�]�^�60N�Ĺq5��=6�u�6�Vh5����8����p�F�7�m��(�)�U6��(��r�j�5&��:�޵�O�50�5��&6���5nn�5�XԶB�96Z�16�bݵN$��Sĵr�=��v(�a*5��5s~�0$�3��.��(�5�z״���,5�r]5B�3�~�C�5�n.6"�6�ȶ5��=�����6*N#6 �R�j�r�8���e6t������<O�q�6�d�4�׳5�5�鶃e76�'*���5��"���ִ�o���<6PҮ�� �5� �56Ђ��(H6�N���̼�Z�<6���5���6(�6MLj��+�}C7�@+6�+���#{6f�t6�(�5��#�O�������6��޶��O6Yε:o��د������76�A���a�5]Ѷ�u60s�6�.:5�-Ӷ��5���6����h�5&��<9C5�����@6߳�50I�j0���'5"�#6�w�58^9�G�6�UQ6�W58��4z�s�L8�4�3��l�6�6�r���U�D�46p$X����5����ݳ��G���r�b�~�f	�5�k�5$����4��l�@Bt3���6��Q��n�Ȕ����3eD�Yu6G	ͶE���|ѐ6~��50���{�>�y��^f6L�жBy˶Q�O6�Γ6�d�5��s4(b���Ф��ж5ձ5�j6��6H?g�$g6O%6U�5�T�5l4�6�[��ff��|��`Va����������j��6j�<�������Ǵ����~5�&m��R2R��p������?��t����6����*����85�8O��;���37Z�5摛���5�_�6�Lε�l�5趵����D%ȵ�'��|����4��7ۚ�6��6Jڵ�J�4����D��6tb}�`�4B���[ߌ��B�62	�6	���pu5�6�Pp��Zr5�����6~���>&�������5���2�$�|[>���6TXL6Au���5l��>Q ����,86F_�5'yh���X��8Sy6��M����σ6���۫�6/,6O轶��Z���N�_���@���i�ȓ�6�Z����4��}5�w���(59�86�m���0�+�V����6�z�60�X6!��5���şF��S�5|���6Yr��m����6n9���܋�3�4�/60؀68�6@銶S��6�՚���/�+a7@��7f�5�}��$/�Bxu��w�g��6���5�7��*��51�ʵ�c6@��6	�~��6x Z�]*f���6�_���6⟵r�~6Ý;6'�96@A��@`^����5o[�5��Y7�ɶ@�)���v�'�N�a�5�҆��Pj6�9�6^YC�44O�s�6��6��5��-7 IX��(h��u�6�wd�0����I���޳t�6 V5��68?���F�6 l86�T�)��6V��U6��d@�6n�7ګt���46�-)�,cߵ�W6��}6��Ŷ�%���l���2����6��5fk��� ��P�6n�46�y��oö��S��,�6�.���s�6c5XA�62�ɶۼb6��b7�O��H�+(����Z� ��)V�*����@��������+�jH7���6��7�<RP6�(J�]G6Z���>��x�O��6�5��66��^�|}ն6|뵎Z@�Ċ
6lڧ��������� R�2=�t6/|�5a� 6��)�Ͷ��6i�������m��6��#��s�6`��4�s��7��6(��̥��l�=��6�T���;5:`6��36(��6:�	6z��k>���WӶ�5�6�59�{6��#7Й)�N剶@*)�P����x�3��6!叶�����768��&���GS7���6-{͵u�6~��bw�6�C�������/5�e�����6�%��0/Ŵ�!�����Y��5�!��\}��n-�5 �V��޾6i�<�N̕��Ce6��z�Q�9�*� 3fV���U�5�05`=G4�6�H}5Hp�l��5�A6
���g6 ��6~��6�e�U"4� �5�x�4�v�6rr�4@�I45kZ;67w�5T��5x�:28-�� .�6<`��������86�V�����>��5N����C68���4��'6{g�5�6�Ņ5���b�j�X��lk6�>���]�X�j���c=5f�[�@�6�\�Y��%6Twy���i6 4e��D5��r5������)���6�S6qYb66�:����g95r�62�x�r #���-5xё56��S��6^z5]��Q9y6fQ6���5v��4
�޶ ��4��5��$5��6�۞6Xϧ5�0���(�x��5�2�3\J�oԾ����5��~5z%��!Ե�k�6��~6F��5X.���c�5=k��T��
��U�242L5 ���k��`��5.�5 *^�T{�"�4�J!����6�� �h�-3 ��2�. 6��6h��jf���յ 54��ڴ����wo	7`h*5 <�� ��ݷ6�Ql5GX62(�6��.�6𡶺�*6+�16��6�{�6�6�4\CE��av6ؙ�5�6��2�5�!ҵ<��4�����_���0}���E��0���fֵ��6&�b�3�_d$�E�O6�/����4�E5 �b2�e{5��w6�+򵄼��^��z��	��6�m�p���by��ů�B��5D�׶A����A��<&G��Ս�~:�6j�5#m6p��#3��Y��װ�+�5u�y5��6��h5:�J�Pr�6YΠ6yC���5~�Ĵ�	�5�ൾ8�5�C��+5�V��5�\�T:�!x�����5ܣ�6����x|�4l�6��~V�5�+�v\"���68�r5���6�cȶB��6v��5��6�;J�U`
��՚��B6`���0��6]S6t
��W?�`�6����)7�nC5��"5N[޵J�涼ʄ�xI�4\�z6����h�Y�PK4���3p�C3��D5�`�6$��6��׵��ݴ��(�k�NA����S442ֶv~6`�2�I�����5̽o5V�ε�Ȩ�	57�I�6|V50�w6�lP�I��5���5}����6#6���%s5���z�4�i��	��~��{�6b=���B�X�ĶZ���aP�5�H����6w��6�z7��e�6UBѵo*y�B�-�|CI�Y�������������5��ٵgo�5��<6769�6+��I�!65˴;�9�!p�	Z�4�
��V˴���5b������6^�'6(L�6'��6bN�4|n�5`�ٵP���웓6������M�������e�r.�6Z��6�<��a#86%W�5��6ȫ�6��6b놵tq�68�z62����9ֵ_���_��C(6p�5���5=�ﵖ�ȵa�A6��5��5�;���ƚ�t�����4���5!�5G̶����C�6��v�R�5�u5��;�x�õ�S�5�0��u��<�u�v�ݵ�V��@p3�T��$�6aM5nĉ5j�6���X4߇�5��z��K�58�0����3���5�����{558ܦ5׏�M��q�D�O��k35<�˳pTi�$5��R�K���0�5܂�VZ
�h�5�h���Z5�
6`�M���[5P�����t�4��F54䌵������?4����t�v4�+���&d6Х�5f��Re���o4O=5z�~�?4�\�3��d5e����紊Nc6 v�+U����y5�!D6�AJ6�>��* 6�:�Q2׵�87�����7��hL��͵�!�6k�F�5I|�5���u��6��4hy���A6x�H�P\����1"��x̳�����z���{��{억�1,6TĆ6����-A�c��o�s6@�ܲr����?1��l�� ��$n`������q�6�m�5:%�55鳴�(��$��5�6v��24�6��'5��*�F�6К5.�W��cx5��δ`���C��~�6)�ﳎ�O�_�Ѷ�a>6��%6�sr5@������4Lf��%P/6T��4�h6򩤶�)�5�7P������r���̊��7����+�`b��5��t5�86冚5TE462���ӵ��6�	v�X#�4܅/6(��4�Z���4���S�|,����5���5\�(��f�5'�} D�Hdp5<J���������6�	�ě6��	6���Zh64��hE6��p�^�6��:6 o(6�g���2��#6B�@5�&K6d�ݵ���g�6�����g�R��>�5[A��ٟ��͛��$�`��5%�=�ر�5��\6@-�6�!6P�A���	�����V���48���P��Ʉ�ы��`����A���ސ����4:�r��IĲk������4�46�u�3[a �^�#�T5*�j6%_(����5f%5��la��?�5��6�!6vL>6�b06�c��W�5@��2̎���6B�#6qL��d 6�r"��܂���K6�=�5Tb���=��a�µ�5*��#�6��
6���4����'�XЍ�x�?3�`5�:+���r16g`5M|P6R��v�[���`��M6z�޵��4J�ɵ�
�5���5醴�X5��5�`�3$�U>?5���b���*7��,5������+�!�6�=�I�(6�Q6/��� ���	��R���>��_6�DI��=ĵK~6�W�@y]��'6�YH���3�|�6�Y
6G4�x^���/�z�P6VJ��L������6K:�5����Ͷ�&?��S5�<a����4ȟK4 �>�|��D�M5P��6�[�4�(�ge�5fyK�M.�5|����H]6���5̓�6�wg�mT�$��4�ӶQp.�u�2����4��W�է��xּ���6(���*�v�Z��5�?6�i~��a6k�P����5bW�����5�5�41�\� �a�鶑~U6P������6�����G5 ����E����5�ȏ��C46�0@�%26@2�5pSE6h��	�6��'�5���8Ri6@��!5�pn�5���6?5�P��5�D<6���8�6ؓ����4`H�4�N6���m6�@Q6 ܘ/��N4"6�4ߺ6NV5r�0�H�i�O6���oe�58���c	6�*�5P1s4��(6&X��=�<5���5g������R� �|�32�5N)5$"�5�/�5~hQ6h�ֶ
2�4�*�6 �2��6��}�	�5`{_�YH6�/�5��7LՖ6
_ 7Hn�.�1����6(5�%��|�������/#�����[�64�`6O�`�2��6�P�5�6�5�P���$�V��6�Jk�l!.6��N��Ro�c���"�4,%n5b����:7�"�pӶ@mS��j6i݄��⏶��6(?4�ё�����!�~6��xj+���uT4�c���\���|�ص�y���1�Ծ�6�IG���b�26 8�4X��4�Mb6�n�6�B=�^�6 ?�3V)�5���3TSn6�R�6r0ζ�,6v����hU7��B��¬3u�@��ON7�&6�޳��u(7���5FUS6S��:�&6�>7�w6,�S���6�C'�h"��z��6RS׶B�5�E.���е[_6�����,J6��C6^86�`�z����U6/��5o�6&( 6���6�d�P�3��^(6��368R�4�W!��ޛ�H��6��Y�	�=��~�5!@�6�\�� �3(�#4׮;�$�E�#��6�>�5�е�C��DOz��D�LݴA�e(�6n��6 �4�c���t7(?6��ŶfmP6��Ӷ �1�|�nܗ��w����p6��B5Ѝ���[����H�-+q6�͵��5i:6c�6�O5@*� ҵ~��Wb7�f6�	6�����-�6���6te6nwt��8�R4��I�l�6�<E7�E$6$��"�
�S�5*߭6�k7���Վ66�5��a�7������5��#7�YԵS6�����I2��Ǥ6�!7Bܔ7�Aڶ�6~����6�Z�4��ȶ�~T6;�[4�6rc��	���%� =γ . � ��4wf�6��y��mU5��6fL0�D77�`�}��(qD�?2r���e6X�w��A�ܝE�E�5N2�d��6D�$�_�U ������06�ͶPN��$��6��ˠ�6�2�3ʠ����4���5�ҶϳB���>5��S2E����V���L4p�+���5b��64Ù�]{6p�T�j�P��s?��6�h^�Cx�6�m���f�n:�6���5��ȵΏo���v�?=6@����
6��g�<8��{�6,����5x�S�(�7��-6�FI����5�f;��f5��E6�Y�60H45�6~U����6D�
6����"�6��E�P60��5�t��6t��p�7<T�h{=�j����5؏	�T�.6��q�D��>�a� �]3�4^6�����$�6%5�?|��� ��5e�B�n6*/�5��5H�5�6F�%6��^���r5L�#4D6z��5`C)5��R�.'�5�� �|�5E+2��
��;��P����6���2�|5��e���6ۭt5�2�A�%s�6x�5 Uܲ�e���^6P�4�596Aם�D�g�95"	�o޵w�5z|�5(�5�s�*�մ�0A��P���`6�;8����������6Жµ�!~�� 6n�ѵ W�4�ζ"&�6X�6�cU5��\P��/ߴ��i����4�J�5���6��G6@�3	̛��g̶C9�5��[5\�(�C�F����p��F6�����#6޶ �\���<Ć�R�5p�̴�QA��~�5��58�66]B��]6d;��Vw�\��6��ӵ08V�P ���� ����5��E��.�5��-6jg ��S�6`o��He�6p|� 703��5�)��hJ]����+ ���N�5� &��M�6����Z2(6�V���	���ų���5С"7d��5�{����5$�|5@[��=J5������)�C�3�;��6۸�5��'5`����Ǩ� �6�2�5`2B��ff�$i���q�Ll�6��y�e���r5����JUy6�H6�A��,z6^�ڶpA�6��Ͷ�j5{�N6��ЅP�P�����`6�q�5�8�4�t�6���A ��46q��^��)�4Lg6�Lb��WE���n6�6|>��f�{�����|�26K(�%�6�S�����6|X���Ԓ��öd�6h�5��:��$6��۶�[�4��5��C�Q���m6@³(z��ڵ�p�6֐4�d�86O><��+�6���6��#�6P6�m��bv�x!�6qv�6��궘�(��.�4D�6d8��4D�5W�5�|"�$����|Ю6d,�n��6plP��<� t���>�4�ok�$T�5J�_6�@��߶���5t��*A6���k� �3<�B��5]X�v[�6�#�4g�5���5�%�6�0�r�ܶ?Q�6 ��1@y���a�����.Ⱦ6�^�4�Ե���4۔�5�%�6��㵺��4���5
�D63F5�Ҷ`�6��6���"�6:6;�5(������5dn�6r�F6b�*�x�5K<�6��6���6B�6�)�0h�q6�65pD�>�6ļ�6L|O6��F7j�b6`C�y96Z
+�/�炵��6`e5 �?/��5"�]��	6t�F6��.6 �6Љ�y`��z�6�I76�#ŵ�q���7�5�6 Ay�@�6��4Y�[��#�6謫5��5 s4<)Զ��6��_5��� >�к������6_�6�Le7�Z�*t?6��%7�5�s�5H�6H߹6p&�5/�ݶ4��5�z�6,�37L�q��Gc6��5"ޯ6-I���y���G���?6X��g�52�K�B�e���7�lB��������6޿6��D�>6M6�\�z��6ڮ��2���5��$6�J
7�1z����5 .-7�16 �5̍o����6n媵��6n�5]��6Nʓ6�Ԣ5����^֣���I6�6�h�6�|ضj=6��5���.m�6L#嵠�M��:7eY�6I��6A�"7�+���ޡ5�n��1���昕5�
7�M 6����E+�'`66:��^k��z��l��2�+�/���6�z�6�L�4�w�6��r�4
6{��6`�1���6C8�Th�5�q��7��Ѳ��a���5�?��j77x�5�@+�2�K�6�M%���_���ö�:f�vN7y��6|<�je�d��6Ƭ�6\��&0�|�R7
?^6,,S����6�@5���6�c5���6��51zO6�]�6r��6�΁��7�157�'�6���O{�>�7<�6w������27��6��2�6xg7�QB6B7�B��~K7��16$枵��p�x�6�4�6h>�6 �;79+�?�8��k
7��۵$��Q7����j�6�6�3q�Β1�F�7z�� ��7�5�!�6V�u6t�6(�������̇6B��5�ȶ`�ɶkZ'7�O%7 '��xY��9c6��	7���h��5�F����5F~��Z��5>V�6X�е=�h��6��]�6`;p����{Ư��c����Y���7��6�<��xw�)����B١�0u��1`�����6�j���5�+7<uw6;�ά?5����.6�6H&��k 6Ú_��&6R�}6�u�5h��l��xs�6�����1U6����?��K 6/�4Lmʵ�t6T󯶚_%����5��6�б��q5�/�6�o�=K�6���6���ץ�V7U�l,�5I�Q��UP��63�i�X'��^!6݅���85��5u䶅t(�cd�6��g���C�#�W�J{�6���45�O6��n�x/�5g��6�T%���T���6�+�6�M�����bm6�{�ʟӶ%sw4���.o!7�8�6��5�7���/���6�D�6 gų��@��3������6��R�w8����U7}C��ȫ5��`5��%��:M��*�6�
���g�7E��6��/5J7�'���5���6�K���Ƕ2��f�k6���6�96Up�5. ���5��"��Z��:����fW6����?45`P5�$ᵸ��5���5��6�[ö�Qy4r�4���j�5V)��}k����6�5�"�v�����<�6�|.6r?�5� 5���5��/7�k����8��J36@�b6�L��趄���9�O5d?6����h7�7P��6��/�`,(���7@��4�+\�2&6U���@N~����s��4�6?7T�G�[öh�t5�*�6��6rE6󹶶�F17V'��Lz�����`z4益�D�6��m7�"*6[@���x�5`v�4���6 ��޴H��c�h!����5��b6+��l�7���h4[��D6`7��5m��6`��40zص�\��6�{��tR�l��L7��P��3�u����h6Y@�6��5�w�b�&5.؇��D6ΝO����|N���y��;۵@�4��9�������q�����5���5F��D��������D�D쐶�*7PG���2��6�66�!N�?B66�u6"�����2f�Kh�����3��5���U�����B�4�����'6�����6No�6'p�6n��=�O6@�n4+!�6Ţ���J���6�Z�Ȋ6@~63iֶh�m6�4oJ�6N�a����w�6��ֶ@Ͷ��5�+]����6>ͽ�|b�����6����*5�=v�eu�69i�6Z\=7��n��V�i��ZmH��7��!�?�5��%�0;n������뗵�D��ؙ������6�\�� ��P�m5�zD6���z�g6��6�Wb6N�Q�rx�6�:	��i��m�'6���6���.��N�̶��6[���(=�5�*��#�6 �I4�Ѷ�RL�T᫶.M����5~'s6H�5���;*���*6�_J7e���"�5t��5 �j�S[v6^��mZ����n���b7 ������`�|4��o� 3����@ڧ���74}o6�e���E07��/5J5&�*6��q5h���"��6������6� 7��@�xo�4:0� ��5yzz6��ӵP�5����}�5�4��6�r6���5�ϵ�y���8�6�}��h�I�Ւ6A�V?050�59��6f�5���)-7W�tE�5���R;��3�5�S7�y�5w����6���xč�t@#6�w���I�������7�=��	��p(��<=6�a 7)a���&7`��?����!7�״6�᣶��s5<�<�2���q6��p5�ڨ�D,85�0 4����a��6^�y��x7�o���$3��#6�.6
���*Ό�c�N60{T��i��rE,6k'
7�����5��95h��!��������˵����|j�6��6��6��"7�55k�����"6r�?6��4ȵ]�<#
���w6�w�5q ����z6H�[�F9� ��2��U�-�c6�`G��t�6�ה5Q�5�Q6���:s�5sKP6��5��ɵ�`�@8>6����p�N��'���6NI�6�\+5,��4��Ƶ0�3
P�6^<A6
䇶�6�N��/�6E��6��&6�Ȳ6���<�j��b'5���W/64���6��q���2���n5�e�3�Pι60�6��x�L"��	��b�6|(7\��S�5�䤶��n5��5lB�5�eP�:468��676����S�nr�5��v6�7��u��)��ڛ"�����>�5Xz�h�
6�l@6����Sh�60$�����6���5�?�4C�6��f6�q�`C0�/H�6����ޡ64���8@�6��3��ȶd5�kf���׵L�6��/6�0t����6'�52ze���X	��c-[6ت���%6��4���6;,�6$�Եab�5Ce6ߖm��ڴ�:�6��i6r�(7@�_���'7��62 ?6�2�6��-6GQŶ0�5r)��r�R�q7o�x.�6��"7��ɶ'��g2�6i�A6z�ĵ~�ŵ�I�6�A,�̽�4R6�$��p-�6X�[6�Q����Ե���2�,6��B���6y[7`T��L� +�4�n����x���7�ش��16Pi6�s5$�M��GK7�kD6�gM5����4 #W��D6�.�6���6�P�5�n�iG�6�5���5�f�.[���Y�6�	��'a5꺅6�yմ|mi�D�k��
�6�O�5BL�� ,�6Ǒ���6���ⶔ����,����5T�/6��4���6�%�5��4�������6,d�6��i6��y�;A̶,� 6�9�R��4E'2�uc6����Ӎ����ʳ��õ4ޘ�e��J/ٵFv6�~ȶ�6��� �y�Xӭ�,'6�05�|�lZ��/����P�P���������&��
"��0�5�y_���e5�$6'����9�Т6��6�R���i6��_����6dX�P�c��tz6��6u"����5 �k�v4H:4�25�5%��rL�5����k �h�O5|�-6��5PK9��Շ5,� �␵�)ӵ���6�X{6��6z?�P5�4�z�"κ6�_6Ȍ�5��52
<6,���#���\5?6i�mk��$n)5	X56��o�poG���5`~��e>\��'���V06��.��۶����6��ϵ�8C�\g����ٵ���H-5V��5i&�Z.^6��?6Ɋ���̴Nٶ ��� �g4�0^����I�6_k�-��T\�(�5��Y6�/���9t���54�,����3bD�������Z�/�ֵ>r6$i������>76t y�P൶|��6����Q4T5 Ǡ3��5�"��X�S5m����k��Ӏ6;ߴ��4���93��
6��6,�϶��<6㘦��`�6|뢵	h�5�!e5wv}���H�ب	��z�4��4��6$�,��:�6�$6��7�i�5 8�4���4&3��F��L�6 ��6x< ��K�6��6�?6��5�Ձ6lM���� 54���j�2����6-6��ߵ��4�S�1`o6�9=��_%4��v�x(�pi���5�I6^�q6)F� DE�
��5�A6D(?��b�6�U��'�4���5 ƽ�4;��Z�d6I+@��y�������6t�'�"5""�� 3]6�8ܵ�1����96=�g6 ��3��Y��y����%5~I������5Zv�5�	)��T���58H15���4696�K35��ݶԼ@6�ҝ5Z�U60s�5̔ϵ�6�[��Uf6R�5Z�5 !1��R7��$���5�e�G;�(%�4$��5��ȴ�"h����5�us��⛴��ȵsn6)�6 a4�������ڗ��v�J�t�(50~|5��=6 ��3Ўܶ��6r2&���y5�(��b2��j#5��`�6�혶�Y���?�6��5R��������䵷�6z轶�
6Դn� ���n':�b�1��>�� @�5^7��n��5�C5Nn�5h�15�B4��/5�9� �w3O�����(����?6p�\50>E��p6Pv�5p9�5n�	�DuD��[?6��"�H�85tw�5��:��¢3}��6�����"����� �� I�2��x5.<���j�3�qg�!L���Ύ5֍ֵȋ�&x64	�5�5hIT5����Q��l���m�	�6s�%�P����96�=6@�14�/6d\��xB3��V6�	���Q4R{��0E�5�4��x4pS��P3��H�U��0"�Fȷ5��6t3�5�+)6 �´�-P5p;]��� ���6�Zv� s�0��pb
�� 5@.� q��E��<�6ќ:���ôV�x�P�/4���A�6/_��A6�N��@��5N?6�&���O���25B�<��5�X5��3�c5o�06Չ�OO���5��5�}S6��q�V[r�B7����B� �_4�*"��J��Զ\6�5)��L�6�����T60�4�/�'������5� #5c��,j�5��ӶѴ�f��5$��Ŧ�5��4/�'�6�C�3^a�6h�5pʵ �|�vQ6��6��4oP�5(B��hJ��X�6��#6��e��.�5x<��pA�g� 6o	Z����5`�z6 V�5lg6`44I�Y�&��fLF6M�6�@ݴ�?��;7����J޴=���h�5��O6@F���&%5:��5�Q�pf��%�����5�D 5��4�0��|��6<16���6?��5ȁ�5�DC5/��6pl�(���[ov�F�5�����p��_#6���6V~e5�ʶ2�6��T�$d7#E:��N��.�5&@��Ɂ:�$��5���6��{�6�e�� ���3�6t�H�.ٴ�	Z��r�����6���b�N�|v26�<u��_)�	f�5L�޶Fς���6�v�3r��秳��J���5ܽ����6�k��=n�v��������ҍ/6R����6�6᭹�	N�b�Ҷq���`��ă�6�$W��ڵ��5��Ŷ��5w�6���6�5�)�����I��Aδn3��>g�5Z=2�$�+�(�4|(۵�@�PВ���25��0�,B�XcĶ�>*6��1��Ӛ�T61����p6>0����ߵ��6X�g���u�B��6 �50I�T��ة����q�ll754��5*��6��������/�6N��6���Ĳ6�6^���N#�L#�P���B�X6���[���<o@6ʻ76��6�����F5"5��6��=�$����d�6Rt��]�6؉)6�bv����6�Х� �Q5�8�5@�����$6G,�ړ6@'p�A{�6bA�6�0��^������5Ӭ�5-��6,����� o6�L�5�6��B5�7��6�J#�sC6��:J7@z{3�9�6.z � @=5�J6��7�摵v�趪=>6���5 �-2�2�8l6`�k�`󽴚�5BW�IY�6x�P��ul6O�C��k,���n6ti6�i`6�J�������h���X;�5H[������6��+���5�� 6Y����ޢ6�j��K0��2�5� �@γ �p��e-��"�5P��5�k6���4��4|(��ca5'm�����26T{���"6���qʵ���4�j�5����$6�׀��u5b�6��i���50y��8� ���G6��4��w4%���}5zq�6��#6_$6h6Z6�ߵp��6 Z��
���\�ôD6�>B5��\���յ4	6�d69=06>��5PQr�~��5���F���d�5\c>���2��Jv4F� 6�յ����50���V�8��4Ύ6Tϵ�C"5$��6�a3�l�3�=�%��o6�<w���F6@ƿ����5��x���$��p��K6@�̵F��5`	��O6 /���q6\��5�����X�!6xH�5Ě�5zh/�����.����3���Dc�6�P4�ȵ�~ʵ�2�F��4��5 	o�Α�ܥ7��͵�>��v,6��B�\ 5��D6�%������D�(��b��z��5��L5 ��1��j54�6���4|��5������6H�N�K���;5�[y6�/6�'x5>�5������5�L=6��x5�A6F������6�]r�t��7�����6��||�\��*FC�u�����`�5�e�4�IB6�V'������&�3*��`�g?6�7�#5�S���A:6?��=��Ե\*�f�ֵ�r���Z����·4"�$�f
k��O��֞5�y�4 �A�|�I��6��5B�5O)��b~�������6�ӓ�����G���ٔ��w'5
��5B/�5춚5&���"?����_�.62"��������V6������d��U6�.��:6���H۵���v��47��6g�#5\��6$<���\D5"N^��՚6��P6�Z7���(A�5�s0��H���nv�ڎ����˴�������5���5|lG5���5LjѴ�)��@Q!�Oa 7�򱴈D4V+�6`S���։6pe�4 ����68���1�2�ع׵�+Ǵ���4:�q6+( ���`2z���[ٶ���u����&6�'|�6ۢ���;6h���v�5]5(6`�Q���X͵�[�4��-6��&6ܢ�6���6�Y�@�7��37��2��D6Ԭ5���2���{̵�W&� ���L�W�6�#7T]���ô6hU5z��6�D��|o�5-���8Gz6��6>_�4Cf޶!����9�6G�a����5,�X60H�4���6� �6O�6ӏ��G��6�p��>ҵ����6ã��/�6����#t6\\��F.�5Z��6>z	�F����W���%��Y0��6d8�6�3v6��d�f�N��L�-]6�L�6�����pM��O%�DO�4��;�$���7�Nc���ضB�������6lPⴻ6u6��v�Rl�E�6Bo6)�ݢ�6[s��M�56��LYY6����v���d<��q����d+f���6"`f�(۝5s�5/�865E�6`�4�%�TT���������6eͶ�����= 6�)�5�����0���T@��z���U��+�A���{��#�68d"����4������"_�6�4vy�56S�5u�����i60|(�}-N�{�6
Ď��˳�g��@,5̎�5VW5��{N����;'7�Ƚ6
��<Q5��@�l`�5��v���|6�/Ƕ��"����6/�#7$^I��6.5d_�5j�<6r�!�"�����6^�6��X�@�i��jԶHF`� �V�QŴ��K�Y�=5��F6�W���u����6�q�5�t��
7�䶴����7��V�L35�Uֶ�:}�(�6+�6�ـ4mE6��97�M4��ȶm�6�a�5���5<?����6��6�̕�6"�B6m�#�p����?�C6�������6Z���]�L��V��z�5�E�5��6��6z=�6���>�5���6
�����q�m6<ѯ�oc�4J���`��4��6R��볾5�!6,�ض�<���?��L��4i�O6g�6T~-����1��ɰ5�\��4��ʶ+�:�a�6��4���5@޵��7�A(6���PTT��6�5���5d��tِ��K���W6-@�5w��6�����6���4Y��5����Z_�5H�4�=7#�5=��|��6���6���6qtT�	VL6�+6�V���6YQ���4�6I'+�D䉵c�@6v�6���6 �b5�X�5y|6����i��6���
/7o$�44a6�﵋׃6�]�5 ����G5 �'����6|���h���@�>���f6�Z�Ĺ&�����ad� 66�~�����ӵHͶhb6���6�^L�H�,�, 7��F���5s��6 ��w)��Au6���"S�O67b�E$��."�63��%��6����15�4i��57�\6^E ��E�6˦
7 ��6�<�6'9@��9���4���$�ea�6ݑ�6��ζ��5	�77ߴg6��X��bo6c��6���6LN?6$�|6�-�6*������6�y6����d�?�j78�h6��F����6`�����h����6��S=�6t�6����眵��%�|i6K�	7ǝ��i!7r�*7v��6��$���a5�	^667��#�H�~7,�ƶ��6D�6�Ѷ4�:�E��6'�51���f�J��*<5�6�b��kj���jW��Ȏ��b5686l�
6���6�_!4awm6��6�������,5�6M�B6�)��W#6J���ϵ*>�5dX#�D�6�ڶ��/�Nڒ�.����S56Y�h��6	W7*���w6ā�5�O~�@��2�\86qU�����58���P�6�66�@ж��b��'�͈7"�?�@Ɯ�_�70i��mKb�`C������kR��Jȶp>���o 7��>����5�5�4Zv6��6(v-7b�&���ڶ0%?6�z
���o�����������5��6G�7�Bt5Ⱦ@5 *����`6 C��X8���p��v�5"��6CV6a�5}�7x�65����h��6I�F6���!�5K7tv��} 7�>�6���M�6�7�0ն߆�6XG���6~p'6L�T6��B��+U����5P�4 �J4�(s��6���5��Ŷ
�6@��5�ӵ?Æ5��t��D�4��6l�ɵ����0(5�M�4�䮵̵�5�x�5�<�6����-V�x ��3n55d3��	�5��4]�Z6�����\6084��6���>�4|�5�h[5 p����4�~�5j.Y��f�8�Q5���6��5h���T�<��6 Gf���N6�.D����5쭄�V��5(N���-��*�6+,�6�µX���"ʦ4�g�X�46�'�5dr���i�x�5�B6]�6���6`�c��6�hI���\�6(6J���JK�5�`5���5 ��5�9j5�����6��&54���6�y25XF�5�Z16`#�3P��5 ���.{��:��5�� 6��{6�W�5(�n�<�)5�Я4���@襴�6�3n3A��`I_4��D6�%�58�`(�?����-��XB�4f�4�15D<��u6��6�@6�P�6�t@6�9�5�4V�H[��`�5��s5$�����6x�5�"6��6��7�6J��� M�'��`�54��5T��61�
tl5x�7�#ぶ�Pd���5<��8�6����J5��������&���l�B��4;?6�t��n��6 34\�5T�4�3|�$�1� c1⑤4�/�4$#�U0T�J¶،N5�75�68���鱶W'6�
b��
68l�4��5�.��'�5���6�3ĵp�Ķ\��񗵶P�6ءE5@�O4h(6:2;��ŭ�d�r��l75}��A�Ƶ��6��
V��vXߵ ȯ4��54�Z�4�c̵�䵀��5�46��f�P6X ���j�5��1�8b�4�=Ե���,FW��0���A6�����5�(6�?0��J�� �������,�p��5�϶�36-�3�fͶ5`A�5����A6�p����6����������.�0�6��5����|���lH5�,B6m��6�������5���#lõ 
��L�ර����c�%�6r��5�9��e��5��t6��ŵ�+���O��dp~6�R�b7���8���+�5�F	6���5[�6X�6��j��C(^6��P6yp䵪9�5^O5�l�5&|�����L���HT����5�).��*6kl�5µ���!6 ��6N����P#4�����Y6 �4�
Զ�w�5t�#5���5��|6��6���X���k�ȂQ6���6EŶ��5$�3��}�5&�6���5���5x�4�rc6���5S����L�U��6�iV6
��6�_ϵ�� 4-<�Sn�5tBj5�6�\�����5bS&6�Ξ6�����t�4�ߒ5p�4� `4��6���4�I6��5v�5��5�H��V�4�y��o���ώ6����T�����94���p�ԵC
�6�(o���S6g9����	���,6���4;Sֵ�%6��5.���z�5�>5؜e��yy6&�6�4��\���\f��e�ߵ*�+�E��466����5bś��ٰ5L$�V�o5�ʷ��k#�H��4!�}6"�R6����)��g��O��A��5l���fĵx%��[�6�t�H�)����&����՗��؉b��O5�D�6�A5�1��|f��7�4[��'H�@x�5����P�v6�ʜ64+��Z�L�I&7��z�(��5�S6R�5Y��6��@5rk����6�,�58��6�ꩵ��?�����:q�56��5^9��L�����5گ��a��5T� ��T��6�Դ5� 6��鴄�h�h�66.�6��k���h9^���5��������cE�P�B��4��5l2D��F6	6���F6u��6V�Q�:]6۰�Pu��gb6ޏܵ�r 6��8ƶP��6�����5q�6@�T�0ux� \�5���~��n�Z��;H��N���8�5;�6��Ӵ�Ю���6�Ď��p�n2m61ܼ��	~6��
�o}�4�۵���@��l�K6j��$�5�e�5D2��h5�暵X�}5�I+6��ߞ.6(��t ��V-*6vR��pK5` �д�_J86�J��(��5�� S6QFضȌ:5I�ĵk,'5*6��a31!�5�G�5����l7���"�5f� �494|���hUյ�;}�o (6�g5�E�6!|�5Ev��YGf6h����5�x9�pO���ۣ���6�q55&6��;5��4����Ƞ���7�6���6��5�i�X66� v2S��6��%��m��k�C灶����d�5�c�3�6oK ���268���ָ`6DcS6���4�\�TC 6�&���H�5�U6��np5H$�5T�N5�/�6 'B4R�K6/yѵd/@��ܵ�!����P6�,	�$�6��H�����w�6Ο�4�-�5��A�A�6�e�5�;86�	(6=�4w�16rr{6�ځ�l��4m�4����6�5054M݀6~�6$�$6R=O6�̈́6�Q�C����3�5������4t�Y� �L2/}��<��6 l�5������ �u5�CS����5��5�P�4��33X�����ֵL����L���A9�5({26n�a� r^4h]a5쥰5P�Ѵ(����K]5��5�ൿ� 6��16�V�5Rpx6��6@'��H� 4�V�5��!�Ƕ�=����9��W��,U60��6dF���5�M6.;5K��x�����6�c��n�50�%���3�ʨ9���%M���β��ˆ5ȉL���{� ���|��5�5���l����5�X���#6(�S6A�I6M0��Z-U��v�����3�hh�0v5"�����[e�����A��p���/�5o*�6Bү���#��p�6�:�6�cr�[fv�����_F�<��� iҵ�[6�ַ��3F6��4Vqf�M6�~h�80Q�\[6-\�5N�m�LDm�8�6#B��dJ6�����r��=��Į6�諶�y�4��5��̵�-6&�q�bz5��?6��4�O�4{g���>96�e�3���5Y�5\����� �X���ε �53�qĴ� '� x6r_6���4�9���GY6R���ش5�@J6&�εT�����6PL���"���� ��oQ��n���Ύ�Cݍ�B���@L5���C6�
U�`�3@�ֲ���5��5n��6�p�x� 5�:g�0*_6,�3���
�5�
�6n⸵��d6�DU6yx)� ̧�������6�6Ƒ��*|:��Qu����6��ѡ��(x�44=�����6*y96D$��f�
6�ں�j�W5-��6BS��Ĵ��j�1ݽ5p�W6��>�����X!5��е<�̵i���o�3���5��u3P�y6sv60�J5$�d��(?5�	�5���0覶h����25!�Ķ�fh5D��50��6��4���5�N4��3l6��y5'�6������5#j�5�6@㴞��5 p�����5,�6A���^�t�C{6�k-6�rٴ�|e5_�46�5ݵU\6��5/=
�E�<5(W�4��-�d�35.�&��nF6��6@iF��6������l͵�!!� �Z6�v�.:���O6ZX5�c�5�8�5 ��5�Qڵ�j64��5@�14��G�?x��x�5ZZ+66�0@�4`�ϳ<��d"&��Č��I5��+6�>�5)h�5��5$�c6������56���Q�6�Jj�+��� ����X 6�sX6��z5�6��)4�B�Rŗ�`=6�ū6�U$5��>6H3r5ʵ�d�6��B6��炵���5E,�H3�4�P?5gb��X������56h�u5Z�l6X�����v4�#6#5֬�6��	5��65�F6�M�5Pd�6�q6�T}6�D׵^���zc�Q�T��5{�65 9p3˥��h��eR+6 ze���Ĵp,4<sD5��4����$��5{�G5���\�ʵt�5@Ȍ�p�b� ��4�q���5T��5���`o��v�@=�p����85���@������������6�*���+�@�P6�L3Z��5�㈵����N�5腛�"(�5��f4p�:Y�6X:16��6�356ɂ�2��LC6�M����6tF5�4�� 6�3F4)�����}�6� ���䴉/�6�H6�I�4�@�54oJ6�H-��6��� ��<h-��VY�"��6J��58�6؇5��6� I6_T�5#�ٶaP�5��µ`៴*Zõ^�6��5B���&�ݵĆI��
�5�H��\�V4�%�Ε�s�5vK	6�M��.�6�bг@��3����XY6 64`��3�l�6�G����� �1@6  1�i�4䋈���6�M�8��5�|
6���i4��s�l��5>}6�R6�۾�qn�6�����5v�����鳓L���ƵXa��,��5�w6����l�59Z�0 d�h��5L5���5@�h5����8v�5s�5�=�����������6.���`y�����$�d�A%�5zG�5�E���ר5�sĴJ� � 5�3�i�5���3q􀶓�	6���r^��R6O8�H��4v�!6Z�5����6%��d�4�N�5؎4@���͛4��9�:bP5�^Z5�ҵ�K�p�K���5p@6��v���N5p64M35�M��1G5 Ј�lC�����3R~76���ا6x�5�T��*'^��� ���%���4|ȷ5d3��@$<���� V;���5��崂z����5�F�4Jj�H�5���XQ76�?6Qy��R}�5 K�3J��5��ô���5�(���)��6@3P����4�7,6p�ֳ|;�6����E�5�}I6�xH6gw�6��K6f^�5�6�h6���4�e�5vl@����5�@c�.�16<#�5�P��0.�4.6�O����� ��1�U�5���<�����k6 �j�\6�r	�H��)6Ĉ^5)6n��6t� ����6L�X6�6Na��I�5�	��`W5́�5���5��{6���5�q���&�2�🶃d�S 6��Ѷ�	�(ˆ5����� �(�VǊ6���5��Ƶ��W5��69�76�]���Bg��J�6<��5Q�¶A
�6�XT6(�6��6p�P�(6'5�y�D�嵦��5B�T�k������ �6�.� �J5U9Q���>�0(,��5^o>�����.5�u���􏴬�����̶؜�403f4
�57���hgH����J3�򟇶*U�6H"յȮ{6 -�5���6`|4����p&��_H�6i6��6��3���4^V6X��4�B�5|	��c�6(�x�f���6�;�629�5c�4�:p��f=6�b[��u�sZ6��!5lM�63
h6��ô0R��I>�.�06i�5A��6����ܵ�wƵ�5�ɘ6z�׶ П���3�jS���R�8��6��l�����|�5~�b��o�4�F'�V7��M�5�M~6���[��6a`7����	����6��d6qQ����7v��5\�6<�6�6�����6	jݶw!�{��5��58�ƴ�N�3,�F�d5n.�6�����%��}�$�/�פ+����6�&6NN��4��Hgj5|7عI4�u�4ˣ��y5Jy���4p2�4����<̶[�6H]���ö���	+6�V6<K�~�� �d��峳ޫ���������5�F�_��t!�E#�6@g]5Ji>7_� 5@ȟ3͞Q6*B�6sn۶�bA5˶8<��8�5�>6��#��?_7�i�3�ƶ��˵ J�6�6��;Lڶ����t��5��$�)�߶;�|6B43���6��˶�x6o�� �03��+5�L붊��5Ƕ�!54��ʵ���5�c�6֛ ��S��N<�6щ� 4�����ab�6�܁��7�֘5:f'6�~�� dB4X��.6�X!� �=675^�7镬6&6 s�6����ר���6p���ͺ6�@�h�?�67�%w5;	7�|"56��+�B��6"|�������5"������u6xT5�!U�Ѳ��k�t�R*�px��&�6��8����̀)6��?�0���p#���]��V�%6]F<6R��6��4�Z赤��5��4�J�6�4'5��6#!3�� H��~6�Ϳ6 Ԙ1 8+4�m6�3�6�%�Ăw6�'ᵈ��
Y�44=���(.7�66A�6���@�bS6r��Ӭ5�0��Xf�*ݪ5������o5 '��"\6��5�(y6��~�l��H�6������� ����x�6M9D�@�ʴ�;��,��6��|5�k�6��5����1�5\���_x�����E��!e5����o� 6��4@kK��?�Cgc6B롶*ND�a�ö���5��q�5���6d�����JG����5�	�5�2x5�9񴂜{5,@���ul�j�6��06�ぶ�Z[��܀6	6�=��=�5�6ѵ�u5*^T6�!6.Nw6(86l����+µ %'4�PJ�B�ѵ��n�F�ȵQh�6���6L�5>/�5=�47�6�ɶ5� 6X����x��4Y5��(60Tv��.�0�5�76�����5�e(5�	���v�6+'�5�P*7M�õP_�3� ��\֚4Q�4�"h��P�p��5,	16�=�~�)�T_"��6�#_��w6\暴ۿ��F@�4 <V2N.õJ̖6 ζ�ҵU\���q���1-�����b��d}� e$�45$i�5�6������M�2�5㜿�n�6������
��5�n��+�q��Vʶ����1����ԫ���-6ظ6

2��nK���6�f"6@�W44d�6#��6d׍5G��� ���mq�6�A������)g��,6hJ>�_�͵��(�2��[n�HD'6���=�6�[�6�I�5�/^6ZxG6|��5���5�%6��*5����S6P�\6A��6E5�6 \c1�%4�%V���N6�;��8��6�4�j�86�76&h�����6CZ�6U��5ā�4F����F����^��5@�3���U���/5@V�3���2᧷5�p�5���4ݪ�5�v+�n{_5�u'6�H�����v�5a�I67��5��f6�e6"�A6R���M6��5u賴X��܎r�F�5j������`�66y�6$Ǒ6�w6r�#6���d��6�y6H~��F���ߧ5V���~\�6���6����W95B���0;d�`a5���5�-�5eR��3#5+A��>�6��#6 N?6l���CȤ6t��4���*���µ��}��5 +5��$��&'6��*6`�p6�@����(��ٶ��`�6��5�.6l��l�5l�@5F_�5��d�α�6N~����6N�4Gn�~`�64�6�)w5=��4(|�jb����5nx��!�8���!�5��a6{*�&�\����=�9�-��f�6�>��vG65V����iȵ�u赉����n&���۵8�����*���-���E����6n9��@4�  y2���5�V��^5�c�5��-6���е <p4\���T��4�e�5�6J� ����\6��4|,U����6��+�*����{6t��W60,�5�-D����5P��5��5������4�䢶\�T6��1'�Q�f�36�k��Baȵ��@�6��6�\����E67e/��qʹ��6`��wK66ŵ5��93�kص�q����E�V"=5�0�MNڶ�=��|�!�t6��Q4�C�5�V5X)r�B����5 �6%��C*�6Rc�����^��6�i�$6Δ-6l��6p!�4=��54��_�T6���4��@�ʶN�'5fOX����(u6ޔ{�pV�ѓf���@�������%6��ϵ�:��Q�6��h����6*B361Z�8��խ�zP��H��6���4��6
�H�X���	�.�#5,�洤ː5���4Po���sv��B6�|�3T�54��5�1�H�絮�������[E6�9���µN@�6�Ft���r5���4����ۘ쵖鋵��K��}��F{��[�6�D��g�5���^m��~�!5���5��5�T��T8$�t�6�K���4�Wp�<�ŴD�n6��
3p��ɋ6.��� W6���Te��1Ҕ�\)��'�5�Jm�d!����4skm5�-ն�2��
6��v6�#G6���*��4�����޵v�5�����2�6���6.�/���?�=��4��6�i��X0�6¨5Bi�&�5Μ5�����6|�Y56g�5O��'���+6C't5�Z6P�����64��-�3��\v�v݊4�>�4��l5��ѵ��7�h����}�A�q�F����	6��$6��}5����3���`5{͵�G�<��5"�6��U5�V"6{6��5LOô\偶X"c5D(-4�[�6x�n5�c�5[�-5����[��4�zu5p0�����_5�u5|����@���6n>�5f?�5mޣ�ܭ���-̵X�Ky6\�\6�oh���� a�F�=��_y4��`���q�lG³'>��w����Qe6���^Cô���5�ӻ���j*)��r���
6696�J���5	��6c�`���Q���յ�,����g�6�fF���M�by�5�[ܵ)6 4��n�5�z۴'��뽴62G�5E�6����x�:6�փ���-� 6X6�y��� v6p ��,ƶʺ�5/y6�{@5��k�H3~�0�6i~��{7H�ᵫ}�����6x*Q3��q�Llw5����~�>6���Q!���6�jZ���6l"�ȎZ�݆�|��6%?6 �6��6j�o����6o����U�I�(�,�5�$�S�"6A{��/�*C��)�|5�.��f��c2���&��|6��g6P�5$�85�I������{e��5ȹ�5��Q��3�4
� �j�6�M���L$4H�V6��T�Rj5�C�(G5���(��5��F6������!64Ƿ�00�4�3N��ؔ�����y�5��G�@,r3�~R�"h�6�ŀ5_ 6 |�U6�0��ҵ��y�6K��b�6���"���G�/�*6��L5�i6���5�ܵ$�W��#-6h�5�����.6  ���M�X[F5Т������e4R�ε4w�5�d��~4v��D2�n7)6(���F��67���6I�ϵ ���4���6O�6O�����P��HAe�t��~�2�XS�6�dg6���Ѳ6������152�����!���c6����Xֶ��%�	��5��N6j�ζ(�5�Z/�Jc���4�5N0F6���6"�76#xT�(���q�� �"6$/���X)�A�5�Yp43�F�����ضT+ӵ�O��R6\Hr�ڄR5ny�4�Sn� ��kY�5Ɇ�p+е�A�4�S�5�~�6�Ԍ�H�6�UʶZ�6�Is5t(3�2ws6��C5��5�v������}�5�T���=�$e4���M)6��?���6 �4�\����5�U��Q%� K6$I�C��f�6�A4E�6���5P�5�ȍ��Ŕ�>�۶g.��1s�<����H�5:�6��g5'�]60G4L*6�@�F2���=�5���b~6@8մ�Y�4������[���q��#6�j�������g6m�632��J�5�[�5˲϶��26�V߶^�ŵ4�F��P��E*��ᬶ�qC60e��NM36�6Cc�5>3����e�������6�2N�Od�6
t2��Y�W���J�6�j�5�蘶r,6�N��6��6 <B6=j8��]�5Y6ȗ0��t7z5�r����ö����_��|`8�"�[6RXn��ʾ5�'d�[n?6���5 �&3Z�6�vU6i�E��F>��66�+�N_ ���=4�@�b���<G��@ճb�����m5�H����T���o�4��p6�a5(�50����!�6��,��x׵#��E�5L^�5 ���(��5Ty��6������B����5�Y�4�)5�0B6�O���#ݵM_6rAJ��R�5��.4��r���ѵR�K6�� �=f�5I;��"�������6t��ft6��ʴ�n5F4�e|�������6"i��K�"�j��5�	6+
f����5�!�3�6mkb�&��5�&�5�8r�d#<��FѶ�jO6��6B��<�6`+6}G`�����^�5�6���"&4��ӵ��5m�6*#6!�"6��4�3ݵ��I5�$D6W#>� �e�(��4O7�5�bs5&t�P���g��$t9���6�\6��˵0u��6�4�({�5�y���6 #6XN�5���5����j��δ�6=���H ��.³���5��ʵ!S69ε\��J��4�{5д�4=%4[x6]��۳6!��5,�ീ�I666-;�x\K5�t5�A�����x-�5�ɚ5[�[6<��4E0�5�S<6"��"/6CM����@��2��=�w�q�ᔵ�jx�66[޵ l�2�3L6G����D��l6��m�3񖴾f6�6,�=������!<���y��4l�f?>5G���u
5��ŵ)�4�����M6ډʵ��൚�/���5%~�6"�K5�h� ����H�)(���H6�ol�|S���,M�`�Z��W5bA����<6&k�5`���D�&���4g6�HC6{\�6_t5�J�5O�a��#�6x�6�U�Ç��,�5Hu����5$r
5�q��x���O�  q�ڇ�����#��0��5@�-��t�6�4�5Ns6�T{6��6�o75�ْ�"m/5�-6���6�	C6��V�z��5�nL�+@��i��[�ڴ|�д�u���ʈ��Y����p?��r� �Բv��4��lp�R�	�u�D�ٶ�uq�CM�6X�[��-6ĩ�6jc�5Zh��!c���'��~�5�5��8T�Ԥ�OGd�^�	6L�"�0˒��D�4ܧB�����-g
6�10�	�F6��ٶ�+�6�@k�̥6R�5rU���4r>I6�ɶaص�k�6�5|�Q�L�@6���5���]" 6������V�I6�o���	�68�6�]ܴ�zT6�؂����6��ݴ(��4I]+6#
6Ȧ 6J��4
uf��k�5�96�'���b�6�F�����3���5�4���]��4d86\��f���)��r��53(>6N�76��R��f~6���5`�4 {G�&f�Z7 �����&�Ι���`6䑐� ��3Q\��)M���058�u�)��5�ε�3g5I�ε�^C5�Ƕ�<�5o�J6Ko��Hr���/�5ƃ�6r)3�:�@6�x�5o��6	p#�H+�5��6I�6�N������6�@G6���#�5})��r��5B��5�g�5,�6��<5�G.��ψ��}w6MS4%/���5��ζ��˵G��6�Wc�́��[����� ������+z6���6�
E6���|�5PV��2��L|%��:6�,6N��� ���_�t�x6��6Q/��\�5Z�^6�I�3��6SõHԱ6pF6�U5��	7�6P݉5��6F\ֵ%[��0�6V韶�pD5U}17b���[J6P7v΋�����f;�4�~�-��횛��5�6�1$kֵ�=p3/w��f6��6zbf5��6 �%��62�6M�X5aQ�<�<�*�(6�%��Q�30��|���?�5�����7�
��s76�{��Q�5�.�d���_N����5� ����6na��|�36��5~<ʶ�~�40Re6bD�U���,���^E4�g 6Ù�6y�/���&��~�5�p��T�~��ʶ%��D˙�_�6����Z6P��p�y��J��v��*��6�	�6_ef��'Z5L�w4��!����5�>:6[�B6�����۶u�5]�������>�6x�&4��6M�$5��յ����DV�6�-<�س#6�F6��6}���Lf��ձ�
?M6:�6�6۶.�~5<�0�֯�����5�bN�"WI���2�;6Xɿ�
]�5��y�0�����4��O6��5��y5�@-6?q����
���82�;ݼ4�"�;N��v�[�,5�<\6��'5�{�4npϵ�ô��5\4��F[��*�6�{ �
{����6��B6GO�5�>5T}�4$��5���2���mN6G:,�$�մ��w6��V65�6"��藩4���6�i5\���֎��[��/��8����y5R;$���5�K�$6�
�5�̣�n��5� ��.�D�6��^�5$���8��N�5�$Ե��Q��a���5��lZ��	���5�o��5�h6C�u��S��F���3((���P_4�r4��ᴈy�5�`�����i�
�L�ɶp��5�n+���6��{5��W5�p1��I&���p���$�5\[R5e��jݚ�G���@<��6�o�5�M6PAx�vP����7����6�,6/�=�酶H�86�76����n6��h�g�A���ĵj��5���"K_��U��@i�5�H54-l�־�6����$�X6rY56��`�?�5��5B�B�^q��Pf[�����6 '�������F�B��V7��R�����Z//��n��-6��G��g6 !��q�6�
��$�d�5���T����A��6�5)6o6����26в 5��4U��5\�2��Ed����5��=���Ƶ�"
5�!��LIڵb����B65�6��k�8�4;�6��5C�K��fѵ�D�4p�*�D��)���-�i���T��6�Q5���
�W4;P�4a�&6���~� ����5�/�*�5U��~(�5���4 ��~+�6�A5 �i�IE�Qݚ���5�J�6�"�� 7��׏� <�4��J�`�:6F57��&_�z�}��y6R�9�����3
e6�z�5���6L���8��&����y�3�J�V����V36lh��Ɓ��PC6�5r�I6��`6{]6�e��k5�����6n$5-l�+$/�x0��b��Dܵ�Y5ݝ�&j굪M7�6=7���6���y�;7���5�dh����2�D6޸@6��l51�A�3��6���6���6f��5?oy6�η6��#��[7����63�y�p%�3������5��?��S)6D��6[)U���76���6y��6��f�u7x�f4 F�����65��$U5�q�5o �T͵���6�fu�I�4��76�7��6�16cc&��6I����5�=�5����L��5���b�۶jm-�9�� ��u/7����>VV�>ь�t޶�Ĵn�C5�X�5b�}���׶��(���@�R~	���{58�
4|�n��5Ե��*6�}5f:�6�����i�����66�54zU��\V�sƞ5��O��w�5�{R6��:6\t�xya����6�w6�=�5;綀��5�*7ӵ�6p�4D�7P�x6�� �%3��7���"����6�_6�끶�"6�o#6߈�TN�61�d��ԗ�/Up6Nǒ5����&���.6B��6M���?�6�ǲ6K�����6�h5`�5I�7��b"6(�L6>���h�a6t|��|;1���5������7�?����@�H��Z�6�T6����k*"6<�5���㒥6*�R�0�5�Զ�L�6��p6�����Ǵ��Ƶ<<�6���5�O��H7�V�O6z�6 �2C����6 �o�99��(:ﶅ@y6�u�6V���ϱ5$t��`�3�f�4g�6Ð6MK$����4@����D6�S�� xd0&@D6 +1��Z5�i��0Ɯ5��%�d%�6���6���6��S5�~�4�E��H8���� 7��"5��6]����5n�?��R�5<�64ٵ�í6+g���36�	6��ζy�f6xҶIMX� �=4]!�6]K�6�؆6��$6�K�6��� ۷�k�.���I5XB�޼�50�K��%6nF���x���9�g����`���Z_6dM5:�6��4z)G5�v��p�ɵ�6�*�Jr�5�Ԧ5���5�
5s2 6&��4��൞ӗ��^b��/�6ފ��!욵Uٽ�.�x5��5�k�0��4i����5�P&��F�ޚ�5�	�S�.�W"�ܬ5��:5Ђ7`��D6�;�r�ϵj(���.�3�6B06��ٵ@!3���q�ⶓ����6�?!6���6D�26$	�5s�Ѷ�Q4X����Z�4�:�6^G�6���5)|���Wٵ}v�6J����6Թu�0d�58��5�6�+{���4���8��41]^��-��S7	7�]4��6>�ε2b 6Ǚ���e����5dp�� �[�lZ�6T�Q�>��6\Wp�Ԅx�漢�X�6�'d5.�464�5�84��6D�5*޳���Q��Y�5��4��5ܘ�W�6�~�(Y�'�$�jm 6��a����5�E�5`%�5^�5��c]a6���4�����UZ�<�i5�6�I� ���i�6x7�6��?�<@53q5*�ɵXW��[B}6�TP6U��T���*v�zi���6𢫶ћ���p5�q���5�6&���f���/6EF���m5@2J�&I��(2�6��06'��K�6�t�6� �3{p,�Py�4�O �*���{6�8ߵ�iǵ�I�5���4���"@�,�����4�o����6jQ
6�_w4*����6��ȵph24։�6�c����5���������8^4>΅6��463�6�����&|6Uh2��`67�ȵ��H���6�
C������`�6�����4n �5r�Q��"����ҿ6{��E零�4!���36��z5�,6R'}��;A�MÀ6G{´hl�5�hu�XVٵ���P�U4����Ƭ�52��0ؼ3
%6�*4��4�F�5�	�5-�G6�Q4�e��m��'��@�G��+6�l5�x6�k�5�ߵ��6�ŶWQ��`��<>"�P���4���Դl%ڴt~�6�`V6��o� ��N�������)6q�:���f��a�6����µ�/6�Ǯ6ط����ą�4�L�p�{5�|t��6�6̀=���,��Yz��6�Y[55�6ȉ�6D*�5Z����\�@<[4rxx5b�ʶ��4}H6�u���܍�Xӷ5;�6 1����5��4|t�5�K�6f�5�d�5�4|5g�6���5�8�f�l6�5�� �3Un��፶���5�$6��5�x�6b�������K6\G}5hgִ�0��H�;���N�ﾈ6�bx�*�����95�^h�$J5@9��i�5�h����	6@� ��#4��V��|�>��6��_��;�^��5n�x6���2}����4/������|�+�\��4��4M�R�f�ʶ��6��l�;��5MK�5�ƶ��ǵ�VH4N�55���� v"6���5ӛ5-9���.�3��䯁���u���5��5�q�5$��5�?4�׵x�/��B�6;�6N=6�0
����>�c9S6s�j6���F$6p��5�B��ҷ�:9 ��a�5 ��C����O�pc��@\36��W�:6橻�;k�� U�6;�z駶Hx66 v���@�4���6���6TA���l���聵D�}���5�W���3�5X�*�ݦ��\7^6.R16�"�. 	�fg��E�ǵ`���.���46�
��􎸴X4����׉�5�ī�㲦�g�,�53U�e�$�8�E�����<�5d������62iݵs5�~P��|25�r�4��G� �2Pl5�@�(�)��x�Z`��y6^ϵ 5�3 yf���16��L5�t4��=�@�3�x�����2g�5�U�ʂ%6x�U�ߖ�5�h� C3pj����230;��~<�cL�4��՟5�� 6���k�NZc5���5{H��4=׮6��5��5tT�4`@k4�m6o)�60����c�v�G5p
a���Y�mc6:i*�m�x5� 7��m6��ò4>H6���� w�7ʌ6!j���m���U�5y;�5&{�6>jt��F�������۴����S��5P�P6p��5��y6�fc��6D8�6�6>F1�r|���\6��S���%����5�����rZ6�iy�D �6�q6��d5�ڨ�eq�Jp#6�	Ķd�6��`�@u�5@#G��1ɵ�����\�4$���̺6,�6B�46��T�ʹ��е S�2��u����5j%6$�p����5@:}�x�D�#X�6ɵ�6p4(�5�t�6Ku��)�5$س6�)6�E��1:6x�5��H j���0�|?��3�5l���D��8����>6h��53���56 ��3�U�F4��{�>�Є��=��6�سh�(�@�Ƶ��6Z��6`���>V��i���]�6�Ye6YvL���6� I6��6�V64����R�5A��1J6Vf96o�6-c���I���Y5ǡ*6�j��J�6	��5���Pa`��]6Ǯ%��ټ6�BԵ���8��6�O4����G0i6'���Ph�����}S6L�5����+5�q,�V�5׫���0�F����Z����L��6d�w6�Lv���z 6$��6=�e�\X��ؠ�5r�6+5ʹ�5d��6�W�3�9���Д6�ܵFN����u�B�ҵ�6�0p6���ٱ6�׽�P#4��`6���0�\6p�;5�_6$95��� ���l'���.7��75NI�5ͭ6��66pa�4�*2���'���x6����&�Bː�+'O�_�6H��5�q���M�6�A�5L� �q.6����=��p"6�����٩5���6�_(�Hգ�7��6�3U6���5.���45v��5	��1<6��m���7j5
�Kv6 ܬ��꒴D�F5��5���6ۛ&��e'6��S���}��;6�Fq�\]ܵ�[62
6�մ5D�6ș���U��TI ��_/6+��(����4�M�5^w����6b���r�4�L��y�v�h+61_���Y�6v*6lJյRѴ6���Pvv�&SI62�����k� ǝ4$J�4h�0���w��͞5�6D^b�+>6J�[54]5!�X�Phv���b5C���l�j��5��F�Ǌ�5��{�@06�.�5��6h����������?��0Op���v5 �)6��5��5&��5�|6 ���#=\�T=�6���D�d��=�~]���A5��`�%յ��5�5p�4��55f�@�t���׵�.l�׸�5ĎN��K�5�_��ԩa5��4@S�x���`���I�t���Żµ�h���ҵ`�6u��5T�������5��5Tm6�Fڵ�S�^�"�(*�h�y���8���5ʇ�5�ޛ6��5�wt5�r5�b���"���h60���Q�������6+4@q.�0�O4�3e��dm��A|�4��5"�&4HU3���´D0˴ �%�Ͷb5V��5�14A�D5���*��5U�bq���i��1#6��5�a���6��(5�/ 4(#j�X_���6v����"���$���A5�*�5��.� $l��f6�
�5`;f���6�6��4-}�5v�ӵ1�M������5���5V���_5��6��5�'��������5�IU5wq����ZG���T�Ƕ�+�5��j5�%���5�:�j�5l��50��3ى,���\�`23�62��\6B��5��5#�168_�N5�na���䵒�Z��s�\#5=v6�?*6���9&Y6����A"�Qb�rw��H<
5��95ty:5��5��1�5��4O�Ҵb��5g���s��d�6D?�5~�*�׊�6j�16�?5^�ȴA-&6	�6��5&8B�����x5����(6�N6@��4[#9�\��53�������4���Q4ȅ�4(�5x������5\_�5w�6e�4��e4��6�K<5!x�7޼5L��5���v��4��:��a�uY^����� ��׀6r&s����4X�ҵPL�x���0�[4?����M���f5P����zj��6LF�6�a6��Y6'5��E�{6���6�5�?��6�I5;���}�5��;6\-����p6]g�����5�U.6�ĶK-.6�6� �5�4~6��e2����b�6��6 �ֳ�c��5S��6�j�_\���϶�`6�ڡ6&ͣ6�a=6�qɵ���5�j6���6"#x5Iƶ�6��I�k#�5�t6��i(�/�5��J5R�ɵ^&l�.V.�Ug����6A�6��6*���� �d˸�RY�5м}4̝o6]��� �X6�����T�Uζw�˵��5�D}6;���ع��@�+��8�5h���Y��̓��;K��8�4D(�P�^� �H5	�$�^��6��4��f6�����E6
�ӵ`k�6O 6<�;�*a��~���Q5[�
6<�66�Ok6�-��dB��d��`���.�3s�86كE�c��6�ҥ�@��C,�L�6n6��.�n)�DfJ��p�j)K���6l1A�`��gd��(LB�X�R�&86@���h���4|���.,��-�ҶRI̵J�U4���5�b�6�5X�
AM5(k�4�M����2�(��!����b6J��64�����52�4��6x�s4���6�	6�����O���gi5B�F6���5�Y0������6-��61"���3���9�d���r���	�
�Ѷ���o�P6��ĵ�uG5rc)6��O�;�%���o�!Pڵ�5�f6�.��"��5DYC�0����1��m6PD���G��6!5,6���0
6j�_5�d'��6�:L6�r6|��,�嵆$6{�46��� ��1�i&6r�6lAȴ�-�5��a6􂨶�oϴ<@��M?5�F�����L�����!�ep��k-5X���i���5S5���崴R6c5��浌�구q̵�G6q{y�s�5�����׵3��5{���p�4��6<��5ʀ�4Էֵ�n����A6�5p6'ٵ`{3�WK��M6��m5X.�����5��Q���I� �v2\Zw6�tI6�k�hd�5�Y�n�6U26H�(6�a׶���6"�5��D�6��s6q��h�'��?�66��\�,ڟ��=�6N+6]�k�7�s񶢄�5X�B��p�{�^6
2
6�0v���,6 I���E�5I��6���:i�5x���F�5PR��3D嶕��6�K�6�g5ƹ�5&%�6�6�jG��D�6,�� Y�5⾉6 c/�n�c6����5��'�y6`1����϶�a�6��L6J35>��5�VH�g�i�_s���u�5��6Cә6Ө0�����x����ց��9�5;27�����
?6�g���(�;H�6�
�z�6�Vr��5�6���V4��7x�ŵu�6��B6.ɤ�<�*��Yd6VC�6���N_��z�5͋����Jж*��d�6�Þ�^��6؝�5S���ۛ6h<x6e�����5����$�r36���6O[��?��*R�68��3�}��e�+�=����+�5H����6
ɩ��B���Ꮆ �"5��52����6@]�5df��PD6�'����51�6�f�6@���l��5���6$�6H8)3��ٶ��2��6p�7��ߟ6�h�4��5�
�F�E����H'��S5��6���UV�����5�&��F�#����6�䶦j865O�64綨'���ˍ6n[M� ��5p�6��V�̶n��4����I�6k˶�͵ค5�@d�\�����57Ѹ	�1<�6h������6v5�C�6�=�����96 7�mK5<M��Z+��>��9��6r��6r�Ӷ$��6��϶��'��Ѷ޸6I�ζ`�ȴ� 1�3ضD���v�53��c�����6r7"�6���"j��J�D��Շ6��:�r6B�N6b��F�`6��� \.4�ً���3��m�V�5Xo�4�ݖ� �3��>����6*[6ӻ6l|/4��>�hm5VFQ��նH��ڥ$���t�ص6�50˳Hz��i�۵� �6x��4��i6�����6N>ȶ�ɉ�>Z��Æ�?�W�w�6|�r�^]W���6��m6�U�6�q<4([�6nҵp��5x�;� aŴ��ڴ|���,�H6���6ŕ�5y꠵���6����T��5��*6X`��(ˀ6,]�5��?5�ĶpI6<wA�\Z�5�>��_)�K�6^}��&(5�M鶠2��~g�6��B��қ6gs��P�6�`ٶ.���G�P�@#S�+)��_(7_g�Ng�6X��5��ӵxw�ઇ���&�69�<6x�\5腞4��&�4⁶۩�6� 0�D��5T�i6� 5C�4�Z2�6Ӻ5��"��S.��Q��6�M����6ޟ�6�36��3�Uڶ�G�Բ��L�p�GЋ5�V*����'��/�6F��6#�6V�56r��0P1��!6��4J~�5D,O�W٠6|�����5004��85�u���c�v�6*��]|��T3��`62) 76����7!fN��ZR5�w6d�w�E�6�׆�'�h�5�6�_6K݋6:��6������!5%J����Զ|TO�Vݓ���26��=6(R���յt�6�3ğ�6��@7R1��S��i�6���5Fж�7��R=05�q�Z�	��U��:�'��|�6&DL6X��5P��4���6@N�4�b4�$�5c�5@�y�LԐ�d�3�b�*�����G��5���Z *7x	�56�@���е�QV6 9�|�*���'�b���fՑ�D(�5� �5�}�4��4(��5 n�46����ݶ�V$6�JM6��6�)���� ��x&7p���ID5>�5�*�B�޵f�6�]�50綵P�V5��0�ގ ����6 �%�#R6.�.���4�d5��z�5j�K�Lqn�=d6016P�6R`�5|�5�ˣ��KI���(�T����sL>6л�5r묶�z����,6�n�3�s5?�5[f<�P~�2n�5������!�5��9�б5�c5����� 6�z5x��5���4P�ǵ��67�υ�095�����6J���� ���ZQ����5z+�6�]O� s"5:yv6�S�6G<j6��?6?ݵ���
�����.76%�4�^6���1 �'7�9��섬����5�у6p��5�N6����"��F�D6@\e��^�4 -����s�5�Y�6rg1����V(��>O/6�_7�����8ݵ�5;����5�7_(�6���Ķ0�L��5� �5�A5��)����6��6��05��^��9w�p�Ѵb� �o�Wmt� t0:�z��5��!6�C-5��ε�^����58e4��4d6~lյH�6ZD/����N�8�_�ٵLx����5�j6�ʶj@��O11��5�ݜ��㫵��+6�4g�¬S��숵�D'�"�5���5(O�4t~�66N�u���ª6)���s�յ!jж�e@�y�u5���4�?=�,�E6$z_6R���:Z��s�}E66�Y����~5�86B{�`����õ6?�6tk52w-�a�n����
�07z�T6�X��y�@��5�e�5�6���u�g������z�6�3�5 ��3X�W� ���l7@�&6(������4�E��+�6tO_5�,5�6�pA��>6(�6�
Y�@`�Nj�5v,����5̼X5X:��(D�w��6����D��V/6����{�5�Q�����<��n�,��c4^�&6�H6��5����#�6�QU�#nG5�5�'S��QA6�(�63|����5�(
7�P6тŵvz~���5D$�<��Z�6T�f>6 ��4��5BHr6�L�6�T�� gų5���B����������@�˶ �6!�5�II���5��O�@6��6�A#4i��6G0��*�D6t!ĵ�;4�j��T�!��>>��Ǟ�����ã�60��6.�k��6:2�����>6�;��c������55�vN��$�ݵ&�5ܦR���J 76h��4t�>�ܷ�5��V5 ��4	я5�8��A���8�b^�6�A)4��6h�5�i���&�e�P�=6�hڶMu�5\��5�{��(��5��δ�z�6��H��q����)��m��7 �%95�66��?68"��|��:I�48i5ؕ6��n&5�g&6�{@4��K�ܴ�
6��6X�4$�T5d21�����T5)�����X5�g@6�C.6��l�J�}5ؗ	�j5/�6.�5D�6�(�5��
5p
�4*��6��g���+6T�6 )˴�����6�4!jl5�46f�5v�e6a�A��5��
��O6��52,�5��5(�4�y�5��5��2���B���� 6B�۵v����9�4n�5*��5�656y�6$�ĵ�7�� d]3�͑�Z����8��i�45�nI�rEB6�
4� o�6=��t�5�P굧f5�%5�𶚮R6̪�5�z��[��6�41�D�5,�յZKp�4��5�e�5�;G� 6ͲN���O��Z�Pwa6�	5��6p������5�:�������_������5z�M�`7�����5�9�5+����2m6��ص�@�� ?��B��5�r鴢^�5jО5� �x��4�=��^�4�$3��-8��"S6��V��ڢ���5��47�5\�6\��sSJ���5�Vc�D&:���L6���3L�e6|�[�̭�x�6��5�*�RM��~+6�fe� f��X�66D�M5"<,6�JM�ā�ɵ�,�6����:60��4R�d��_��/5�Z ����4ĵ��5��z��%��q��R:���r5�p���6��"��jj�HWӴ$��5�ŵQח61�A� ���"r6}�5Ά�5D��5��`6���p��5�L���%���]��;(��6k�$�=�|6��B��95�)F5`v4�V5��6�ɍ�H��5.!5 �-���o6�<�����r�5���4�1�5 �M5�ǵ�ۯ��#�6�~��J6l��@/�N�6g�Y�N� 7�G���g�qd5�#����Ü�6�X6԰6�f�0t��n=�6`w�4�̲5�l޴�
6 '�6��ȶ�h/6�x6n4��RD�#k.�w�D6��J��#���Q�L�7=�6����=+6O�J��״60��,G�51�46�06,�I��$�5��$6A���:7�3�y���F6�)�p��5��T��u�6J(�54f<�P[���p%�������e7��4���ʟ �6�6^��\Rh���7���5d�յ�A&����#�?6�0�6`=�c-7xF�4�l�6!ީ��d�62[6D�)5E/�H�25��	����6W3�5�Ye��6�"D5�H��Μ6��̶8 2���7e{~6���6� /634���� '4k�5@hk4�l6*�6C�6�qC��o�5ɔ����6xe%6�鶀aE3N�6��6�yS6'����6!6��{�0�B6.�R6��26��]6������ ��_6V�4[�:6�M�6��p��6��6~Q�5�����_�����qo�5�	?6�O�5~i7�����5��N�X��@�H3(d�m���j��@?60��h�P�7�ʶ) �6�5�6�ص,r6h)1�����DP��0��6F/6OV4�_�5�@�6 ��4�%�5�m5��յǞӶ(J��=,�hg5vK�6�ʏ6�ȏ�D�D5AAi6`Q붂��6B�t��6��$�㮦�|��5*�7�R��dW� *=2��d��6��b�w4����6�%G6�_#��е|k5��k�Кm��T�6xu�6/(�%���#ζ��H^굈�j6HO6U^�,6�k�+n�6L��M�}��6�7���t�õAN�߿X6)g��A���Έ5茓3�%Դ4'#�TP��^FY��Hǵ�K	���h��5vq�������7���62�L5�+5���6���u+�6��b���o��R��,E5�u���X��苔�tOi5l�	5S86v?G6N�ⴚ0�6G-�5��w�h�4/��5ӹ�5�9��U��5�$5���y��6C�m��:7��[|6�.��̂����!5wzD����4`�6��6f�1�^
6z����6^,6(4A��_�5T�ߵ���5��u6�5Lߘ�hЎ6�V6�n5v*�6�r6�K�5q�����"��p~�6�4��%��6 y458��u�5�16Y����U�5�,47L8�ݤ���54�d6�3?6���y��LZ:��M(�*�A5R�F���"���f6���6���^a�}86�2N6�@�5��4�O6۔���F"6ȁ!��*�5��\�Řg6��6&�3��-���?�6��6ph'6�:�3�ٺ5���3���5*;�x�{6�j96�����u�3=ε�@6z�R�jh�5�V�@�(���6�s��6̛{��	� ��p��4�U���=󳥗�F#c6~�5\����F�4ĩZ�p�ܴ:ƴ�a�5�_
�H˴ܻ��j�O�/�5~Ti5���;6P�p5�4�4�ޅ6�6��j�[7_����5@[�3�~�r�6HF�5HlI� _3;�E�ܲ�4���6�}��e%�305'���짐��U4���u4�˳�z�V��5|�����ɵ;6q�ٵ<�60W����5  �4k�"�#�	6
����|6�d�5H�n�ی����4ܼ��:�6 ġ���>6t~�U���y�6�P�5,6� ��ƍ�4lF5F6���6@�`5q��6�VC6ӑ��I��qr�5�jc6@�$�L�Q��J6|9�4a��t&�6;�6�l�6�f}��/5@ɿ2*�6T�4�'������5΀5�P�57$�5�ˍ5U64a36���/�.6�:궵mV���X���z6�z�5 �b6_� 5r؇6�!v5�K�P��30�U4Eq��n����:65O�4ࠐ5��Y4 -���
6���5D55���5�Vr�j�M4bK7�6��5:N����öo{�5\!���g洰r�6�T6�EF� �^���!������Ք3eK$�256lP�Cn�����;6���6A��D��5��e6��5�@���s�Ѷ�vѴe��5Õ6-��L������5�g�v��4L�9�`l��q���_5x��5�5���n��!E�6o��&��5��2��յ2 �6,�Ķ�⊶a�s��8��ذX���5��ε�j�4����6�D��Ou����`����6v����(� p24A�6�r�5��Ե2�R��I���е�$�����S�^�'��ٱ�U���j�5�*�3 �6ܕR6oG���࿶�?��߁�ަ��}�5l>����6Ś�&���a̶��=6C�6}ؽ��;6;�)����6��n�В�6���3�;I�@��3�Q�4�"�P�5Z�6��6���5O6�7� �5�h����6 �J�Tv�^�6r� ��6�������5��絡g���6f6��N�d��{@ε�ֵ36i �5^�7�1���W�4�7M6kX��>�5�$���,5P<5�.m5`��4��5j>?�$d6v{���/�2�l��v\���5T腶67��ej)6 Dr2B�6����$'7$�)���6ն�����&�K6�=��a��6�a�5`�o��_26�t^6��k��k5�O�53���E�C%���3����5�C�5��ٶ	6]n7���4�2qh��v��8�=��W~6���5H3�D��4b�6�ϒ��K�����P���$�t
!6Y�X�d��5����iu5��ж������|���N�X�5�K�5\��5��ζp3�5u�P6���6��5 a�22s����k5�{�����6�ͅ�d$;�6�`6�de�ַ�E׏5*��1���5ܹk5N[6���_�K6fv����5:Qm6+����5
�����r��4�?�5n�������g���"5�c�5t��5ȵ���4ؖc�B3�6`�&�Ϙc6��6��5�N�6�5X�3����=6��6�	�6�Ev�xt��
�L��j�3w���
5\�
��𕵄������൘��55By6H�4*1���A�`��d%������G<���6r�G6���/+��q5���6Q�6��?4(��� 5;�5*gc5ho(��ɶ�x
43�6���b6([5&�L��r-6ʳ�թ�::6�6P�P�4�4�6�?�6(�t�)6̲ٴ@���z�"6s@5\ˀ��<���T�w�6��7�h�>��5��6E{g���*6�䵾���X;�5'1�6�m^�h��X!Y6Cg�6��f�߭675��3K`��X'���g6�ʹ6�Q�vG���t�j���&r��q�)��55��6���e��
,���N��$�v6]�6͟�6H6�8���,N��p�ߵc*�6nS���.���2�v��>�S��Ǡ6����B6���5A�޶���� ݵ�����5�T�5�)l�x�*�"�6<�N6[�e�L6i}�5��57�S5� ��
E���>�5��5���5x�5�e�����5�i�:h~� �5�l���O�6*],��T�5肋5��2��9��D�C44'5
�ٶL�86���:�6Z(6�C�6����d5�����>��l$��i����04�\6*ѵx:B�'66Ox�6�u�c��4���%X5��+��hI���s�p�6�6��26���5~#Ƶ�ٵ��5�6����@�3��4<����9�X�x�&�5p�� �3l?�4669�;6 �0�n��wJx6�.���P��{��1��YJ���4{��5N�Ӷ�@6̌C��h?���е�����"�.����q5Zp0� ^6�	2��?S6}(v5F�J�.��2�5���E������vû���6f6�P�6?���o�����4��4r���gc�4x6Y�J*��ϵ,Q
7���5�Ԣ6*�65��c� �� �!6�!6��c�>!16誶�@�6 ���u���xG���=�6�l�����I5�e�5���3�z���+76��X6O�U6��5��`5��i63۴��9��(�5Ɔ���y�5���z��6 �W4V�� �~�Μb�������B6���3d?U�
/5�|-5�J0��=T5��䵂��5J{ɵ��6ә�6�-j6�f�AY��X��4eD>�h���-T6�㪵��P�3�ֵ�ђ���j����5�!v��I����5�2�R�
66%6X�x�6`訵:϶P�J5{�(���״1u{6|z���ΰ5ߴ�tɵ�*�,A�5���h�>L�1%6`�¶����lP�4���5t86������6.8����4J��5��5�z���|5Nc4cO���9t���76Xg��"n 6��:�@�"�L�3����6�v�5
�4�I�5µ���}���76
B���L�4(�5ʛ��OL6QK�T�57�;6eM�C(�5�aٴpN����5Nҵ}u޵�ވ�*�6z��6��"'5'��6����(���ݴ���+��œ��۵�lM6N�6�ޤ�Δ۵Չ�6��M6DL5�HF�*i��~O#�a�5`��3��C��QK�^sN6v�6��4�0��ݯ���26*Z6���5�y"����5 ���6qhV6��6��6����5����� #��[���+5��6�t��=<65�6 (�5�޶�d�5-H�6!$��f�_�	6̶���
6H���z��+{6�N�����3b�Ҷ0�ڵe<m6��	��RD�jˬ�ǹ�����`_o6gJF�U�5v謵��@�nl���eɶ�)�5�gO68
�6;��5(��3��6�����>I6�Y�6u��6Ɉ6F�O6K%L5\��4b�6�}|��B���8�6�,����>��h7�����d���6�׵�6&Ä���&6�.6��L���5dx5���4/���/��WW4 FV��}��p�5Y�f�`6`.ڵ�6������r�5��56����H�n�c&���C6�z7P��5��5K���j�5�%V4��,6���6V���(h6r��������5ݓ��6�y�6;��6��'�T�-�iF�5��5n�����6迕����x�4��w�Pڃ���E5 ס���5GĴm�B6���64f1��76D�öo�]6�ϐ4<�D�FBr6,�6� m���V6�H��k5FX06�O56'�ӵ=��6�5��"���L�6�r_�8�6b�6V6������QS5cS�0�5��6�xԵE!۵\2�6BTq6���6�H�3)ʶ���5%ݶ��촲P�6�)66���6��G6e	6^W�5�1$��d5Ϩ06�w5j�V��A16�ݖ�7�l6�ˡ�',86�&�5�X�6��6Tt����������{c���6�@
����)���.5 _�5n�����6�����a���*=6��X5�X	��97u�S���5Z����h��4$n�5����K\�c�5�L����6b�����6Ђ��"�?6m|�6� &5r���Ѥ5� ����*68�d�;Ku� ���*{�6 TF�F��6�f+6�6�5�$6����^6 о�dle52�6�'��8X�5^k0�Z�
6\z�4Q�684ִ��d�`Q�4P����t6^�	�v�9� g��+�4�`��<Ѷ��ٳ �d3��7bJS6E��� �6����Ly6O�൶�6�K�P���$���s���t5�~+5�!�5V�Ҷ�6��>56��7��5��6Lf���?�6M~6�ڈ5_#6x���216p�05�6�8=���S��5�_�6������.6!sc�����#����m=6�_�6~ �6�S����[��觵�g�3��40O5��6�ݵ�nB4@O����4�z�6Й���~0�
��7�`FB5���B��`f���)�5
���5��9��@Q��┵�w�(^�4���5��>��bõ�0��кǵ\�굷϶�bE55�pi���)4�L�5����+0�*F�pm���5�dԵ@�3t��H��5�S4���0�n����52~66&��6hT)6�E5đ)�P	R6���B���V����h$J�<
6�ε�a/��]�4{b�6f�06��&T����6`�3iWY5�Y4�[Ŷ�R�56�;6�l��c=�E�52�5�|�f�6��]�5�(6F 6�H�l&�����5tm�52++�n��6,ʈ5��ܵ?Ԯ�X�����5���6m�5��k4Z3��0Ѵ��3,����x�7�l��6_��/�e6�W��UO6�^�6���5�"r5�M��颵�	��S 5�ހ�v�.5,��4����N۱5���5h�4�ʴ������3�����6X4�L6� �5j�5�9�����ݵD5�)�5�s�5�B6�K�6�4�5��*6dSI�<���t�6�Op4��6��@~5 �#��s6D�5�ð6d�����6�@6x65����e*p5��d4�b84�a
6PW]4f\�6����#Li6V��6L]�5�����4�L5Ƽ�6pK61����	$5�Q��O�ĵ ��3Z�6`�3p���D������G�J�[���<��Y58P��Z�6�ǫ���� 1�!ٓ��'
���xmU6V%�5�G������ �6^Tn6@P�5�p����G�給�H�� ��`s��X���(��*�0�Q1���͔6|j��x�ô]X�6�Lk��b5���
M5U6�/���+���J	��G.����40Rn��K6""�Z�z60�X�|6b6T�Y�l{�6\Aõ��b6d_�4�45Y��6wE�5���5��=��yG6�e��14Lp)5��&6Tw�5e��4P�!�H�̴�,K�@�4��Q5��3�O 6�	�P�4���6��5jBE6�!�6 �?4��ѵ�ݵ�}5j�x������IJ�� (�F������3�.��z#d�L1�6�X6��{50�6� h���%�g�5 ��5�����6��X6񪊵>5�Wj62QB6�B��p����N�8�E��6����p�׵Qnζ��i�����^��q�R6�X(6L-_�b�`�x���66d�3�������͵����de6B� TV2jf|5��
��fR6@�����6��3���t����6.�����5�$%��4^0��q6�R}��ĵZ!<�g� 6�|8����5�(4��6�e4w�Զ:^�N��5�a�6Ҋ6���5�a���?�N|c6x\���M�6Z�6�6�v;6gj���=z�4�F6e	6`��5>(�6���6�{��Ɩ�7b6��(6Jګ6�]`6Rtl5g�6h���и��X46裵�64�6�M��W�54��5�A�6O'75��5�,���浂����h�z��6:����5Љ��J��6T�ɴ�ق6>bq6��5��3跻�  7����$�6�/6[�ȵ �b�嘛�&v&6V��5C˵U����-���>�6�L�5:���O�6�DZ6�b��Ժ��\O�4o�5��g��Z�<� 6b�u5�ݵ�MG��]�|��4�����>5�Ƕ��,���(����5ȣ1�y����|�6�T-�4�k�Rg*��(K���6�Mk55�õ�3Q���p6$P�4gQ��p�5h�F5�����^��PP�4��6ૉ�p��5�wg����^�5��5�um�x�C���8��5�,�86�m�6�B�6�(�5&�A��qG���c��c���h��Ԇ�s �J��5 � �x�b��+6hx���6'H|�%S5�@���56쩏6�Ԍ5Pm�4��N�Zh(6\�Z�Y�A7x�.5IP���޵Xnc� 
	�7W!���t���|5e����6M5��76�(K�δٴ,�
6a_�nm6��5��
��O+6���5�+�o��� *�>�5R��-�4�����X4Ҡ �Y#��~N�6�a����&�$5�I6 �\��J6F�5�˶�ʅ5�k�2�d�4p�����$�te�EB�5H��4m�I6�?�4����w=���m5�56ZT�3��5��Uމ5�}�ƶ����g6�L�4<���=6|P^4@X%�@�����6ƣ�6O��5"�]���?5�pI�@S�5��J���6��5�R
6�K�5����1�K��I������U4�����x66n��Ԯе�͙59�6آ�x���(K��5�5贵�	�4��6��5���8�4��v�46�|�5�u6�26H{õ�?���G6���5����6Y��') 6�܆�bv�6��Ͳ���6#:f��õ��yo5ƨ6/0ĵ.Ik6���������5.f�����6�w�5u��X	�h�*6�S5�说�RG6	_K�ҩ5�(�&���¦�5i%��.2�5�E�5T�$6�&��0�J39g�9�����4��?�@���ҷm��S4(� 5@��4
������5>��^O�4�
��@E60�5�J�b�/6�
5��5l��4��F�U6ھ������r��5�zn�-�95���E6�H4R�
�rc��"ᵣ쵦��hO_6�C%6������c�Z�������t<�_/�y8��
��4Li�߇����961')40���6�6�8j�!�/6+䡴�5�/�5QSϵv���f8�6�h5�#4�z�5��%�>�)6B�O6q�5��ײd�,�ak�5�06������[5����̨6:��50��58=a�V��
E66 Th6�Uc��QD6�I���24\��5��Z�f�5R�5͍õu�k�"d��ﴴ6K5�V{�=�6k>6Y�5���0�F��!6���5���5��6|õXy3��k���i5�!6���4#n�5���548�5��,55B5Nǝ��o��A�5�m�6PU5�%J�?�6�����t��K��5P��5yi��������D4��5?w5��;������&︴�����q6m����Qq�~a���������*�<A85�<���'�5ņ5x��R70������_������5CݵF6B_5�(������R5;��6r:U���6��4 g23�j�5��W���o�p���$d�r�T5�8�6\�5b?�4n3��a\6?��.��Au�e��6`��3��=5c	Ƕ"Yɵ��j6�5 �1�p*6<�;4�����6�d�5h���q��5�a�5R��. �4К�3O�6�kV6`,���e6N�˶���5�:���w�4�b��p�'���6l�O�6�!�6��4����@�h���/6Ln�5��5h��<��5hy�4<6]و��ٶ�����V6�r���5�8qm������X5��56w����68�!��r�2�w6|.�5~�C6�{�5�p�`, �����Jǵ0�F6<I����F�P�X�D��5#��>Ј�2�U6�f�4�|�5��7�B��\ن���5�ͪ��P6d�L�
�P5��(�h9��𤵴�)\6�J�5O�W��a�xZ�┏��S4T�75�$v6VLj��^��0�Z�ﱇ�"�5xM5����5#�)�z�6��ث��\���5��5K�Y5*R��06õ����n�4=�׶��F��rK5��H��,�5�����O���q}5�~f�H�h�5�V7��V5�"$5m�3��-6��(��}�5R���F�~��64V�5T��W���
�HM�6�R[�p����C8�`C,�|6y3�PHI4
�G6��p5/MM� �7�ʵ���5�6ɔ��ܶ��d��o��5�>6�F'6 �(�\�������G�:�A�B�t6�^��<T����%������޵��F6��6�z��cԶ�7��}�6�����W�x���~�Q�a?\�w�[�M�z�p�µU������6`�t�~��5��=��qr�����lө�(u.��1��R4��C�l���D��� ��3V�{6^�p��#�5��6���6X�x6�����0���G5pv�6 ��4��4o쒶�G���v	5@s��Ai62] 6�8�6��6>��5�ƚ5H�66�7��1��m��ȍ5�մ��6<���#�5+P4�������5��6�T6�vY6Z�)��}M5��W��`�6�~�5������5ض�Gg���빵�!6'g� C��w��+5�� 6,����m6�[��{��5D{$5�⚵_ⴶ�U6��ε.���yA6o1�.�5p'���6ӟ��L��Y�)`�tI�5�q,��Ӝ5�܏5I�0�pZ~3����<q�43�T� &.����Rˆ6
ֿ4����d��á6(x��[;�씶��\6�5�r�4�Զ@����61_6���6�������5+6b�D�6�.���5�|6�P�62g����5��5�55�ҵ�ω�^2z��:5��5���5_�6$���Di�~6��4aE5�䫶s�y���6ǽ6PL6�`"6sƵ�ڨ�{+����;6�V��<_y57!N6d�J5�r62?6V�?��!U6�=55>���t5f���5����4���4����EQ���ԲNo�mf!����6��5�"�6�����׵5�6�5�`c3Ā�m>��D�5�X;�:�ܶm�4\�\��ՠ5��5p��3��䵨'�5S�6�(	�����,��X�4̺�5�����5:�Z5ԅ�u-^�dV����E6��6<0P��#q3��H6�w!5��r������5O�6P{>�����lE6�Ay6�5���5�l�h���`�56,�� d��4���P▵�5Ӷ���4N�6����U��5������6�+�!6�j�3��%6����Z~�0�5׵����F6��H�:7�6��
6;�^6��g6�a���k���g���6��D�KM16�3B��R�4��5r�"����85��	6R�5��g6t�h�A���ۂ*6�����6���gۮ5V��}�e6*�5��6@�3j��5��b���[�1��6ҧ��At)6 �D6i�6�YRX��]_6�LJ�F��5�86>�ܵ\�6�٪��*26H��5���*�	� )L��&��}�p{M�R��6\F�6l0���.�69=s�� ��\��r)����6�,��K6��?7c�64�����x��6��7�����vU���5$���P�5Q��6v좶/�Զ�y�F��6�Qd��J6��d5@�]�g7�GJ�fõO(����r�ܰ���z�������"5�ח6�!� v��-S���L6���6�!6�k��E�4x��5�#��f붗�16p���V��Ә���6�T�qx!�7�����F7��56���6��_6{8o��]#��g��8�=6|H�6I7����hC�`(!�l�N�4�E���7���5B;���Ke76�65hh`6]�Y���y7��O�8���I�-�d�z5��@��ʱ6H��6H<�5<P �Je���e���� T\�#��5wp�6�&���j�ڽ���5.*%6�"���"�"����7���dӾ�H�����6޶S6�)���[17$Uy6B៵��6$�����5�j�2M�6�������lX;5WK&7�n���6�A\����3��� ��\'�5�yd5����7D7{{6$���P6�6����p��5d�a4Tӊ6���6p��4� -6e 6�T"�m�27L��6]
�N� ��D6�1���Dw6�r�6�%
���7�r�6^!)���d6�C�5��%�dh�5p�5l�0�Ǵ6۩�6�<ƴB��6�i�������2�6<i��ؐ�6��p6(�377K�B��6E��b��5@q�3tܵ�,�`�z4�-;7`|	�6U{�w��@\�6����H˵�C�4ؐ���U�5���6�<2��E6f�ĶV�?���^6�7ȶG��*�6���[ʤ64@������[�4���������[�5���=��6�L�������Q6 +��?�d6�Z6Qi���&��e�����x7w�7�?b6�P4�4Q�@?Ӷ`�$5q ���86����:�|��4��`7�˺(6fL´x7��7�)ֵP� 5R��@yo3����5��h�յ�d�5��5n�#�h����<���o���6砵��5paH�����t�7�7��@���7xu	77G�6:��6:po5�A�NN$����6�PI6������16�pc4k�U�)(�6�B�6Y!�� �6�X�<�����?��Ő6��6���49��56k�5 n4@�� "�4�it�i�O5�b�5��4n�{5 GW�ɾ��69�4 6�X4�g����6q�E�Y�5,�-5��v6:��Ȁ)�8�4��д|R�Dʯ5��5^Μ�*G�6v&%�Ћ4ν6n�����w�
��5"*6z��6���m��6���5bT����?4�q���j6 ��4���T��5��.�.�6�M:�.:|6�6_��5x�Ƕ>�r�����X[൬��5�Q�6�Ԍ� k%4���5�'K�@v�#�[6�����g6V�p�U0�5G{�`�y5�u�5��6�ʭ���6̸���c6�]��MC��\6jE�Z�H�%�6��=� $L6V���x��Y4^`��A 6V�-6&�t6R�7	+�e��5v��5����(��΁x6�����UZ��j��Ʒ��{6:ߒ�dJ�5�	д@��� qZ�h�6B�v6���4�C�5��ܳ�Vε��#���P� ��1�8N���x5�n;�W��0+4��^6�6@Ck4ވ�����ff6��O�<ӵ���4v�f�6��5'��������6��e6I96,]"��C;���64�Z6�)y5d@����M#�@��i^K��E�5���� 
���4�&�J�g����6��5��=�6!�6,�6.�ӶXTM��ٵ�T����9�A6V���dV�l�6�f�<��5���ʛ}��7!6��5����3��\fi6�!�5Q�5��M��\�6�����&����y5���S6܆�SY�6�aQ6��5���6�h1����6�36θ��ΐ�� �`�+5.�v��M�6
���X��l�?6 �m�l ����6㔶��6�����8�h�9������6w�Q�5�JY6�3(�j�4�8�5���:E�5Z���J�?6��36���4�sX6���4�'�6,6�?~������ک6�v�6��P��(u6��ǴOǞ6x� ��h��l7��5q5p�Pza6d[�Ԑ�:@����&6,:5X-ն�ѓ��	'��6�����|���O6�Iö8U=6a��bmQ7�F�6��6�&͵��8����6�̫6DIW��8�6:��6ț��Z�;�YP���6@��6�/�5�>��K+��l6�sU�,䐶���5S|6'	p6#��N�&6�PI�R�6ԝ�6xU��U�5��M�"l��|��5�v����̶�B�6�+6xN�5��{�>�f��a�5��z6<�*5��6�ø��g�~��66b6���֔p��6�6_��LX���9#�@���Z5p�l5�M�4Z;�5��!��[t6��7B�*6�8���j38=�6��~�9"��'�6}���ڋ�9�9��Ys����6�Y�6��!�l����l8��,��27��׵�Z54i�6�#¶��)�DM����(6b�<6��7�W�&.5ʶ'n�V�06 ځ��n6n	�5��ϵĢ�����8�7h��42�!�fS65���6�&�����5�ގ5%�f6�0�6�)��wPC�_E�� g�6�?&���+6<��6> �=�6=��Y"��,�6�{6�	����6p�m���6����(�����j�6�27�4/�`�Q�<�$7�W��CV5A�P�$��6��4�@笴����^�8�@������
���m�6���6PW7rH��}���fzm�.����7���b.&���߶_f 7�y���qZ��)��p 7�=�5NvS�]������"�l_8��ꁷ�/�6���.F��X6F�_�6�76}W��>7ϡ+6�46��9��*�53��N���3����M{���x6���4�V����5�е�0*7�>�6�,�6��H��;�5	����Oz6���5��5vM>7~O�5�J���O�6!� 6�c>6�_��Fq�6�Y�6܄���b���;y�.8�@.X�vwF5���4����M/\6呎6  �6'�5��O���6��6�;D7�U��.31��jC6I��jrڵ���54ێ�p��4�����5�%r5��˶@;�� �絫�|6�����q���u�@(�+F�6O[��Z��6��N��G�L��6�f*�h�y�@?��v ���6������� ��l�4zl6;&�����6\n@7l�5f�:�jU$�`�4t�N���5D�7�/7̵�Z&��Bn86��6�8(���k��6q,�Zh��(�ߵ�dI6"��.0�k"7v(
60+����6�T!��;s6��7�V6**a7�OԶ�|� @�2Z��̰�66F7�u�65�6�,7�SI�4#�5j�F7��N����6`J�U��p��5 %�3�8�8��5��m�x�6�6�p�4�-�6<�Jq�5�_���M;6�m��V%�6$+f��.˶���6���6�Q�vqQ��E6s���!���|]�	+��r��6� ���{���K�6�7g�4{����{6�+����6���(�
7@��p)��"'6y��6��4�O��rz�S�6����P/[5�����`�(����5p�#���5H ����� �֯��h-e4h�46}�6���X��4<36��ϴ#�]˶����J�6\�mP)�B5�6D�h5�{�6��7��A-7�P�6�^67_K$�K�1�X�M6�������~�7 �5P�%��%i6��׶$T���,���ڶ��M"5�E)���46S�6�h68�6�T	���6�&7����8�öE��8`�5���Ka6���t��6Z�(���&���� �6�cG6Z����a�6��5-�����5@i�5�̚����6�[����5vꨶ;�76���6�}�68-	6"\O6y@#���ᶦ�F6�Ā6�O7�!6��5�
7 �ζ-7h�l5��޵f\U�񋳶 ��L�6�$����K7�����BK6�Cy6��,s���c�0�f6g֟��9/6D�޶����4��6 i=5B��5��ն`�m4��ӵJ^1�|�����5�?�6� 6���34�7�&�5��3�H���㮶�r�6$�߶�7�88ӵ�x���n�6���6���5�2�6._�� j��R97��ݶڵ<��R�5D6������P�&��щ6
�7��L62u2��':60b��7�\h�:	ݶ��q��9V��M����6s�6tU�5�/˶h�[�x� �Ӷ�MH6�߱�;,��I�6i{$6�=���6�FC�����ʮ+����6@L>4����5��+4�7���5
�7g�����8Q�6��H6$�6���4�=_6h� ��0�47p46.#6pQ�����5��!�*�7W6�9J6���5�����Ґ��D�� l�4f,ﵹ}-6���5@kG��0&6僰6Ļ�7Y�X���6~]������ 6p8�6b�+6sH7*�B�X6^�����-�6t�o6	7H��`]������>}���6�-6N�b� \B2���{0�6ɝƶ������L�h�H5��96x�Զ�6�c���6��w5�'��2���.6��Q�p���l�6�t�d��8����q��i*7��6�r¶p���p7�>�5�q��?�j��p���u최:�6�-6ؙڵ�~�5���իA6�ǎ5J�6�
2���5�MC7��Y��Rt6v��6%�6�$���5*H��!�@B67h)5
�5�z7��\69Ŷ"��6����?��� ���z6�����9���,��_�� 7+8�6��J����6�M�5�U6�1%6�T�6�A,7:0@��a�3|"�����4�a���v�6���5gy6>uu6�6#Ԋ6��7�:�6�i�z� 6�%�`���Xﯶ��ѵ<ױ51TO6Ь�	�� �ð�ި��(�M  6�����6���5��&�6bN�5� @6`�i�@!95F0"���6����T��6 }4*����4h�6��6���,�5�;�>0���S6C���}��|�T���6�ܥ��4)�2�6��5�u16g�N4��>
�6"��6�4E�������6���ڇڵ3ǰ6 ��3��ӶPe|4�{������&���5̄6�k�5d�U莶�>4�{?�hl���'96&E7|
�6.N46�X�A�Ͷ���5pb͵r ����6�.6�{
� ��6 �g�?�T6~�봴162/��оv�7����q
��ˋ5������)6����¶w�6�ص	��6N��,�W6���4H6]��6�o��&ۆ6�B�%Y��P36�T�4�^ζn�7�7!6�0B�F��6�y(6p�H��5@�������b�6�n��0ɵ6HX�4Z#�r�L�Ή6����^G�6|�
�8+���'�\� 7T`@67�,�>zѶd�Ѷ0�E���?�~�M6 �5�f#5f;a6&e�*�4��Ա96*�6��7`yҶxe2�0&W4�2�}����Ƕ�}��)�5:��Y�7�q��8]�6�Z�5�(�5��6�ͮ6�D�|�*�v���5HŶ���*�#�7�5�H�еy|d�����&"7�)�4��6~/��mlŶ �6��5��B׎�j�h��UI���b6����F�6���.z�6͎�6\Ͷ>3׵���5 �O606"~F6�d���w6eQ�5X14�7�6�6J�i�𞐴Jၶ��b4���6ݯ}�����z��*�ҵ�_Ķ6�}6��v�XE��������5�	��ȵ��6x����m�5@Q�3�a��H�H��b�����[�6VѶ��*64�\�j����5��H4�h�6Fy�6�"��.�o5���̓6L�6x�6��*6Z$&6��5^֝5o�5�+��"g5�c�k"$����k���}��k�^�J6��6*�67�7pë�H�4�jD6�~���gr6����Vi� �;6�j16�K6�9O����5@6���5p5�5"6��/�8�51�^�c5��A6�볶P8�����,Z6�*6���5�U��d�5�8@4����<l��\� �0�3 ÷�G�e����v���Xo6O&n5�Q�5.���Q��+r�]�:6��/��g�3򹵶���6��=N�5DRX���\ʵ�d6vYD� +���N5V���O`7��p44l�!O¶켅6��m5V��5�k�6�_���ҵ4��50��5��k5D"*�F#c5���6_�����N67�'5���5�	R60��2p�6�u���҇��R'6^(:��(ĵX��6�a6�3� Js4�X��vo�&a>�dǶw����6�5�>)5�Y���p5gL�5��4/S��#-���͵�/6k
�����6�S�5S�6&�4�Z/7�P׵�)G5�>Q�*߶�>e5�"��@���``H5^? 5 £���6��-���w�\y�n�ڶ�"M6v�L�|(D�Ω�6"F�����5���5�/Q�e�S��6	S��)���N6mz�5@���J6X�#�j���{�����6�ɵyw57�u5��b�V�ʵ4��5�A�5hyU�r6暻5���QΒ�cʟ�i��%c}6k����3B^�6Bz�5����� �g"���2��6~��5l/?���,�vCʵ�ǵt6�Q��S�5�z���O�i*"����n���D4�o+6��`5�w��&.�"���ϡ5,����3��("�H@P3��� ����M.� 3x6*ל�HkH��76&�r�b��5wg���R�|vʶv��w��0�J�4O,6[	P�2 ͵�b6��l�0Ņ��\6|H�6ȂW6٠3vҳ��\鶴E������oJk��芵�*�Gn.�i6��5��o5�"��Ð�6y�d��p���#�5NC6pQ�4�`������(6��0p�5��ֳ�6���4�f�7�R��^�� 	2��5��6$�N���E��5߳�sĶRŶ�v6H��6pv��B5��5�B%6��6��04 t�1O۶L��6�o6��y����z62'�59v�3�Ɏ5j��$��5"b�~r���>5����_��V��6->���f�5�5�5�17��T'6�#�5�P�5Бu3�I�4 OD�t̴D�6���ʂ6���5>Ց�<�?6_����+�4��5�C쵬�3�8z�6蟫��׵.���M��M:�5��7��6N|�B��5��6��r���܊L6f"���96h�ϴ�2*5x�K63�?��Є� ����浪�[���6��W6p���c����T:4p|�4��_6�ԙ�dˮ���Q��=���X!6��5R����cF4l5v6,��� �t��}ֵ6�l� XJ��I6�֍��H��h036��&�Ld���+���E� �2�5�Ƥ��u�b��,j�4��O��U�2#
e5�-'��ͭ6Nɪ�)�ٶ�)�:�,��%6�J�4��6��(6�FF��-�5�l�5?��D��5�b��m ��2�5�u5-������B���y��&Ӷ����ƿ�6rs6��ŶN�k��'N;6��� ܶVQX���v��o:��5���
��"#p����4�P5Q3�6�l���*����5.��5��6��u��1#6v������������5���5�R�8�Q�6�A�6+�;��,��^�;6�F�H;ɴ\&涄}5��6�Vr)��(\�.B�5���[qz�pqi�n��T�嵠�:�j�#������6D�4z!����W6�f��h�J�ؾ����o2�?���3� T�2�`�6�oD6�s��:b�*��5�z_�1�`5"KT6� ��5~9Z�o%�ࡴ�dc�5�(6VS���/5���5|x}�5BI6&P6*7��Ƶ ����Т�E�96���5��޵��5�6�5��4l#6ZK6d�L5~���cƵ`~��~��5�Z/��ܞ5�|�5�!6����=6��i5��4��6�hӵ��k"�h�e���s�$�5��5����r�y:,6�y�6�'���5h�A6Z�66�
���BB��H���ŵ���4F.6����9ƶP�6RYʵ�h�3_��5�B|���<���5�74�{����tz6�E6w����5�jo6��@6�H��!.�6��l6�2�5�ȶ���у��èB4p�2p4���#�p���[����c5��G9�4v6ВL6� ���F5��6�T{6��������蠗4�y߶t�+��-m�Z����ҵx��5<�P�p�ĵ� (�
9�6]E�6,�����b6v�i�?�M6�����6�~$�wPµ@t�5^OR6_�����D.5 A���5!lL��4�60�s�T�c�^���+D5���6���v6�O6r]�6�TS6���5'~�)-{4l���D1��x�j6��6Jw5�M6E6�	B5��C��W�6]��|�5�����m޵��p5���5Ǆ��z9��`4��5�)���O�(
"6t)�۲6#l|�'x�5�k6l�ǵ6;�JƵ�~16�дN���R���N�5
�5�(	�ȥD5u�M6�@A5�R۵���6��_4Ȇ"��]4Ń�'4�6D�g�.�V��fе콶X�_6��V��;ϴ��+6��5j-��jW6�/��a��������6#��0s3�Ɇ�ȡ���->5�@�4��i6��Y���0��h���*6l�~�Ip��k����v���3����o�D����6:�E6��6v��ͷ�69���(#6�M5h,5 "J2Г"6P�l���g5�}%��+g�p�w6f%h6N/#���5�e6N~�4'�y5r���rT�6Dl�5� ��a��XT5�z��o��˩��>� 5Y��6Nie5��v6���OJ{6��5D6(?�5 �вm�6t��5T����;L�`�|�:��5��5��5�b�����4��N��B5��Ե�Q�57wz5 x����� �M�bb�5P��40~�� ��2�LV�cXW���6riR���p6:�[�A�8�Yy7�x���G��K�¶���6ϧ�5L�����9�5��64�붞�Z��{�5,G�5 z2 r���W�6��y�K��5l��4d%��ྪ6h	��Z����"��}.4?ۮ5af54f�dt�֨�� �m�o�6DM�69���[�6�6A��蔩�t�5+��5@��������(�,M_�H�˶�76ǵ;�W;�5ȁ���郶y.��p�6��5DG�%v�P�3"CH6��a��:v�6N̩�!U6��4����S��s����|�5�#5606�� �E��56�ά4
��5'�5â�5N�5�F�@�5Y赀ր6���6.��إ��0�a5.E��"���2$5^�F� R<6ގ�5u�[�w+��@7�3{�3޶�,�f47 �5���� O�21���35'6�Q*�Q0ʵ Q�oH6L�6���6�1�4/�6�|5�6�̵T�~6˅�6�Ņ5�H�5�7#5�6�5����ZM6�sZ6�	6�Us5�{|�f��576-'6�'�5�sC��е2zX�p��#>�לq�z]4����5h3k6\�6��&6S�6�ƛ5�� 6
���>i���"�@�,65T��[5e��6m�������t6zlo6��74��ܳ� ��%6�o�5�È��g�6�5��5��6r�ö�1�d
6x!�6� �lC��A��҈6�J�6��_��$�����-N���5�&6'�4И߶�'6!ĸ���,�pW4�#ƶ%������5P	5�]ɶrH`5��P� 4|�5B�����6J��õ�3�v5��䵠R�����5	R�p��5,���j�6�8�5�(K6��6ԑ-��r����4-��2�G6@|7�\E����6�NN����6O�E6|��f-��l�5�!G7������6L� ��6�궙d�e�5�^����ѵ� 6���3�7�5�����6 ��0�:L3u��?��62,Զu#��e�5Ml7R�i6)�z6�2�5x<�O��6�O��q"붠�3��6���6����!��4�t�5xޤ��^�4�5�5.��25׍��h��Z{���5�i˵�/����6�� �l�S����6�o��t1��v�6<�(6:�%�DW��I+�6�Զ@B6�g㶰p�6p,�2��5b�867��6z���$�5&�6X@ݶ
}�6�W�e����ϵ��o�D{�64�G�i	�6p������|6�2 �f���YA4��j�%]��Ώ7q۪��Q�6޶�5p��4T������^�v�Clc�s1�5���3��g5vt��$�`6����� ���a���5 e�6��.�&{����97�o�6j�5��v�6�4���5g��6&k�U��i���Ф�6��6�Ɵ� ��٠V6�e{5�1g�VG6�O4�^� ���5�6���6�,97^��5� 	����������'7�G6�@^6�6w��r�6��$5<�6h�ʹ Zp7��n����:�g6?�?�\ǚ5�9�6�,A6C�1� P7�~6��6�͙����58ȗ��7(��5�����V�6_�5%����
��<���6��6դ����7��{�$��6EBa�IY6:+�64+6�����������,� �;�W�6^3��""�6(z�6���6,�ݶ%ݶt�6p'�5�6�D�������;6�D6��]6���6�E�6(̠���ö��L5yS7DZ¶�v�6S儷�������7�B�����6׮���5��~6l�����_5�k�f�6-��6�$I�`�@7��ζx�L���1�j�`��;4�Uk ��$ж�Ԁ5F��#�6D�5���0�7�I7�g�@����)�e̶�:E��X����j����t��1tS6��h��6�UM4 t�5��6���[�(6h�崐#6�Qt6�$��H�6*J�@,ԳV��5>��6��54�5�a�6��6N^/�@����Bw5�=2�@J�
��M ���m�&O4ؼ\6 ��5 ��6v7	���M��W�6�7��1����v�'7ϵD:5x�����V���s6�� ����}ܶ@��2��6�˶W6�6��3om�5 �����5DP�5N�,6����T�[5d����6I'�68E�@��
�<6$a�5��Y�����ϵ^��a##6�rѵ ����@�L�|63�>:�6���5�t!6v��5�i����4�#�6���6�.��AU6�چ���5�	L6�Z��ֶ�n76��5HZn�`��#�޵�%6"��2���p�h5|�5��ʴK��5XsI����@e���%�A6���,�5J۵�����5��H��Bk�p�g�6Uc �+��p��5�[6>�35��65aU5a+�6�g�zVF���+5ϑ�4�w6$1Ӵ<�u��%���6���3�7��
��CE�WVk5$�f5(.��D�4���5��u�la��iܙ5�����5|�:��,�4�o�6��_�v��6pvu�������T� 68�95��w� M����5��l5@
��,M�4݈�9��z7J���7����5�^6�@��\(��`oR�@�B5�B�5]�5�J�5��l���g����u87�437s���>�6��5���5�6g�<����:6�x�6�M5 �f�V�5z�5J^A��s�6�Z�5��k�@��6��e�`��4⟶
��6��68a5"�D����\�6��5Ԙ���Y6)2��P�D4�6*5�4���O��p54P/�4�4X���.��b�T��5�S͵0�4��248��� �t�C�����|�_���86I{ε@�v4�&&� U��u���-ȶ����@5����\\��$ڴ��7�^층`���ҕ��ӵ��5���6R��6��O���(6�Ъ��9�����Jj�5�B
6��5�)H�LE'6[;�5��+5 y��چ95�76S<�4	_�5�}(5	����5���4Z}X�Ċ���}�2ڌ����6��5_���"��5�Ǧ�X6�+<��K������j�-�����д 7Q5kY۵�
���4S6���(4�ʞ5;�˵lHV�NSB�ٕ�0B'5�V�5�x6�2�i0���_�5���+6�p;6�C}���\��4����v�)ݵ𵹴h�`�-�������6����pG5Eȵ6���s��"��Pu6��!62۴5iw�5�Y�5��͵��X�h7f�bq���4�5�O´t�E�(ݵ����%����)�6���(i�+�25���4�/6`s�C�3*L]5�n>6��)�N8ٵ�̅4�j5|��5\���d5���5}��N����W	�6S6��f6�y�5/k�� �5�7}6.v�50Z8��Xl5�.}5*�ӵ0�4��5�wS6f�5ziC6�r85�	���I�)����df� pz���5g���t06�8���fU��� �4�M��k*6�y�5*��5"�����5�#5����p��ZS5�0�iԁ52��5�˵�H&6 H����6Q(#�M�V5��5�
^2w�ڵUf����=��{����5�p6��6s~�ɽC5C؝� �^����N�洬/$��Ǻ���5N��5�Y��A	<��.0��4΃@6d͵��#n��a5�W.�V7�5�6$b��hE�5f �rjh5t� 5J��<I����+���0����v�CE�����=�#���6B���S(5�[�N�!6�]�5&S�5�> 6��5��5Эʹ�{�4ݨ5z~���06>rC5Ĳ6)H�u8�5��>6�Q�p��4�[��a�b��>�.෵��p5�����*5@��4_6T6�V4@����4t��5 ���9��u���9����6�F_����5��R����4�P�6��Ӵ�F�6���x�O4�����:���V�6�)�v��5�@6��е^gr6�<5�z6�*�6� 86`M��V�o6�!�N	6T3���<��������6zi>�^_x6�|�6.T6��۶ �дDނ6)�5�>7���5.<�5�se6Zz��xpF���:7?B��i�6J�r5.6V�7�� 6)L!5|���S6Cҹ��c�6@�F4ⱐ��w�4Q���H�?^��r�5��� �a4:���I�յ�q�Z�۶g8�]	�6�-�6 <��lŶ����9��p�#4���5W&��u��5��6�n'�r�s�+�}�.d���6lӵ��}�����]��]��(��4��O�4�7��/�H�5
6s6 ���>���K⚶��6�7����E��h��0�5 �������f���j 5�Köt������Xa����25GaǶ�X�6��Ӷl}��q6
����:��>L6̛c5��5��Tܵ��㵜T&��*6������ 7�S(��A/�IS��(=��p
�6N>�6t8V6ꚿ�P���X6uv��L�5�➶@���G�6,Iõުd6�h�����6��:6���6�8z3'-�>�55� ��*�5 	��`K��6�h�5���(Xŵ1C�5������b��P��v���Z�5�b\6��0�fU/5ă�����5>�7�����l��9.��7&���B@�_m7`��q��(���¾��\6t�O6=:#�̕�6����5}���:��#� �{3�"�6+Ե:�6�d�� ܲ��[51��6|�:��e������O66E��6�<�4- �5��,��>��H��b���ң���6c��[h1�E���|�p� 5r�I7@�5r�7bG���A��N6���#5d�U5(S|�KY�3@7M����6ҠH65�6�6Ӻ�� dv���$��M*�$��5Ž6K����O7Oֵ���o�6�H�5�Ff��5¶�:9�^ն����A6�0붬q�Y�̶�(H�h�7xȣ���f6Aə� �R3
�6�}.�w\���]� �N��6ҳݶ�06�E6/k&�w׆5�6*i7���5�G��/���*7 ��3d�̶X׶d��jr#��V�6J;6��)6�c�6!�Զ~Ҝ6 �1/�����6@.�63��6�~͵46���b6
����+�6��5��6TN��T5��X�J��l�7��8\L���۶��$���"4:�T6}}�6� 6����'��vB�����)[;7��5T%z7�陶���x��4w㿶���4���6Nx������*聶 �7������6Ҩ�5x�4K�A6�A6��޶f"6�J$7�\b6��6)�Ե��6�;���6=�6>R|6u'�5C炵�H62x���� 7�?G5���h�6G�������n�68r78:��C6���54�ҵLv����6�R�5��5�IƵ 6Y���@�6��!�a�� �6�ö[{6��37��=�q�(6 �!����x&�6v/��6P6@�-7h��^	7QƂ�ߤ��5�*6b�� hW4x1���Ҷ���&g���C9�Qu_6C�6T�-7bY��Ǖ��Ԋ�\�g5�ݞ6��;7d��5;'�6�k72���\D���|�6�i���W .�����Tе��6�ӳ��	5�I 5�t�6W4��8�49s�5��45u���6���0� o5>��h�.5�S�)����p@����5t�_5�kx��0	�
�6�8�9��`F���х6��6^ē�X6R������8J����M6{���~�5|7�a���7қ5�+���� 6�U961���I�5o�:6��5����05� ��4y�5^�5!����W�aF6$�6���)5��N��4�x
��N�	7t��5��5�El�6!v�3��6,6Q�{�&��6�4�Ƕ�6�0L۳)85��26�a�����P�F6I��5Hb�5�vo��%�6�s�@7��pۗ�,w6��6�,�6�]�5�L69�5p��8����:;46Ud۶��|��W�4��ϳ���5xp�4|�37ǥ�6<��N#S��_60���#�Q���5� �5x�!�~�6�R�#:�J�86ʢ.5�h��B�~N���@_5��u6./P�)�ض2��5�9�3��>����PΪ4�V,�We���G�Ӫ�6o+�6�ճ���ŵ�Y���d��r׶�Ƣ5�[b���6	u�6��5�-�5 �n5�6B6tߘ6?�6����>�B6�5y��5��*6ٹ5:��F�,�6��5������{�yI6��_6��65G�86r�U����4��6쵖6a�5� �P�l�g�	6l%0��n�6�{4@.=5���6Ɂ �B����5$����Г6��5+öO�6.��6i�!7 pU4��6������P<�������|�6^�A6�r5䠔�.���*����-6�k�4x�6̆����z�5�B6������>�Je|�A��6\?�5���i����쪶��6cv�5����elW6�Ң��?����|�ƶ����͠5��5x��6Jp����c���4�k����6��`5Q��6�v�5d~�5�����.6|5 ���M6�d��^6U顶�E5�x�5�˙����4�6:5�6�յ���5a�6�{�J(6�⵶�u���6�n���A6�$R�:���J�6��5���6P�+5U�;6�׵�>ضy�I6��6rg7�>���ȵ��u���6�\[6X�I6�%/� ��2+N��SS6$���E��ڊȵ"L��6 ��6F���\��oW6:��5z��4lkY�� ��ؙ6��5`Vյ��e4�@���#56ံ7������6F �4�ܮ5�����3/��[5�(۵��	7��6�	2L�6a�&�L��3�4xb�3\��5`�[57���ǲ����6�w�6  Ӷ���5�7ɶ�`6�&�$����a6���6XO���dY�F�ζ��6���52�S�a��=�,�?�6K�^�ZT��� 7������)�X�6<�Y���%6�`ɶ��5�^6
��5U�¶:y����5��W6p�85���|N����6	!�H젳����Ȧg�zo�5P�D5��6�e<��w�5񭤵o�����>���eL
6��C6�-��>6��o6�O�5�I_�S/X60D5�7�(���E�� 7���6���z�ٶ�?�6Zŏ�'��v�۶����>-�5��!7z��54Q��d
L��	g��"ض1����F6$;��\eq���t��r�5��5-X��S�5����������6~:��p�?��︻��6exl�d�7Kl�Ȣ'5x�6�7��vLx6�	t�'d 7�?�6��붂`�5���6�~�5H�d�VFd�
��5�T�6/�6���6�H[6��3�+�r86ۍ�4lR�5�j6}ȃ5r��6��I6�9F6�t�5Į��In�K��5.�7h�4�U�6�`���]6�և��ﶜ�ĵ�����+9�\`.6F�U�Ѯx6J�ٵS��6DM6$0�6Ob��b�¶��4�G�V[�6R�A64��5��Ӷ�/6Tm��Ž�:�D�j���|+�a�������\��5�q�5*a�5\�6u��5�����y��6 j5@�G4q���x�9���e6�6��ڴ�~��g�3��
�5�߱��x6�I�>�D6��%���O5�M�K�����
�6fY4��3C6R��R�J�@�F6���6�۟5�p�5���6�vP6��|;�J��6XG�����5�ƶI6��[�2����Jj�N���_�5K6�_K6�;���tr5�^h5ق'��n\6%��5Ee6�o��an�6Ǫz5R�6�����5*�z5���60?�6�lV5�z�6�c5��^�m�6�̶ �6K�k�Ĵ�5���6��=��6��U6�[�xPr6DW��<�&���}5c����?=�68��5H��5�"��#r{��F�5���6����2V��6����f�������.�����5�I56h?6��Ͷ�T�5������W6�u6WR��.6�y@5zX�4L�6�M7˻�`�6a뢵� 5�R�6!��5(���)���Rs�����3l5�I���Ա6j�6�nE��\��6������ɵ`�d�I��5
K���=5�ͯ6��N5 �4�8�e��}�&��4-:5����յ�6�[�68+�5L��5Č�e�5B��4�&���:� ����P�6(�Z���5؟6��4+��4��5�k?"6,��6��5?�5�7u���x�/��5E,5����5j�U4`�6�'60�µeɼ4M6,���|��5(�>�E%�5�D{6J���xY�5~l�5\���Ǻ5>���J4ڐ�5�h�E @6.ٴ5�[Y��"�5��2����5U�ѵ�����f���g6�Ո4:�:��6�9��y5���u���@60?�5� �V��%�5�����ℶ���6X0?3�&J5 ��6\��e���N"5RW޴T��55�,ƶ?�J����(65��5,~T��}�6��V�+�6
��6T��53�c5��5E�5q��4����wĠ5,�:��&"6���3�%���h�����5M޵x#�Ns6u�E6�2��������|b��Y_6�֬��z��d%b�w��6O���^�5��$5c�=6�6n�S����5�=o6GAZ6Gl��o6!��6����-�l5������6Jx$����4p��6�C05#5��G��C6�0%�;�6�u�6� �6��44��6X�=5�>`5�F6�H�Nu!6�f6 �(�7��6��7�|굆�
6�⇵�s��g�E5�$൰:����"���/6`���F۵��~�~&浡`\�����fH6R��5J�5&i6����� ��˳�5�׶U�G6JB��m�M��='6u6�0�5�5b"��	�5��5*6u[X6{�5ξ����ҶEH,��tZ�h�\5�I���mj���L6�.6.�6c;6��Ƶ��6ۧ76����FH(7;Lֶ,�O6Ծն� )�S%5���6pŤ6i�1�mm��M5xFd7��޶r|�{�6t˵��O6|0������fSE6R.7� 7�L7Ld���Mϳ�~7��5�N�ܗM�:�g6@���dX4#�#6��ش>$�X����p�5k�6w��6�N��6�6��E�4�6 ζ����*� �H7Q��!��Z4��O��5ab�6Fة6L�5^V���M��h�!�
$���*��v�6*6�{���2��x��[�?7�C8�!�5�l5����5�����6�l�4r1y6��A��ܬ�D�]6�	��2��.#�6FXs5�Џ6��5-�C5�#?�觴5ah�����6ɓ����4��>���˳ ����:6N�;�Z�6/Y�5P�5�R�T"5��6��+�n�9�X��		K��K��y7ε��i6����U]��I�5B�U6*�ŵz��5�hZ6�ZR�猍����6���)966�b���g��}�6�&���M60�t6��6(�!6��
@����J5�y�\�6����>�>�y5�:6�C��dd�N�-�R�'=�D��5�ö� 6K�6�Ĭ��Ӷ�E6�6,4�o7v��6D.Ƶr<���mX��h~6CʶV�6��o�
>ٵ.LU��1ݶu86��d4�74���p6 �޳�n�6C˶t�K5��16��5���Z�f����%����p��f�<6Y0��� 6#��5�L�6�Z"�E���i�Yl��d�6�~6F3�5<<��g�/6n�b�F�6��:�xd6��������5FY55��" 6H7\���Ա��:5���5R�5�D/6��5��鴶x��	Ȥ6��5��26$~��&h�{��5DL66w��y5 P�5g)6{�6����@�A�I�p����i.7b��r\� ��3�ô���6�،��6�a��lOd�L�5�w�4cxj����5`����d5z�V6�նzO=6Q�6䄒��2�`W۵�V	�јJ6�ô��XBҶ��(*�4�Eb�0گ�f-�5��6��#��h�6CJb�:�M���6�c�ȡ��@z�y��6��g��u�6�vz�:>k6���V6H
W��^6c9&���5����̶�6�G6���k�!��6�v�ۃY�3t6��5 "0�@0�5�R��m�T|6"ʤ��)��^��6����D'絖7�}C6�%�2��P�5��3��۵�}��@�}5w�4#�6Hȴ�J@�5�[��9�36
|69J�*��`k[5I�/�<S�5n}ɵ�����)�4xI`��Gv6$-y6L۠�w@�-����5�Zߵ�4���8�������6����?��5ų���R4p�S��ԃ5t4lj��5��6�_�)�ٶv,��,OT��$����9�����nx��i��� ��2�gW5�:�5	6��ҷR���y5H<�4gq6i������5ˤ�6�y��:����"n���/6�2�69�.����$�F�^z��5p
J�k3N6��Ҷ �c�#�6B�7�;��K�)���h64�ֵ��6F
Z��7 � ����J�4�2�������56�5�u	�@٫6p�W6���5�6�-�IO�6���6I�V-$�����.��6B���R5�Q���'��\�7�Gᵸ̜�\��x�&4����ޠ6�g���6 �"��S�4���6m,���]6Ս�68y�z-Y�#vQ6��k6�S���6�v}�2,����Z61�7�+����6��ҵ�����?����54ąh�Â��F�5����6�j6�ꚴD�16��	��_*�Ĳ�5���6���5 �6Rǘ�h��h��4��6H�6�	T��OK6l�2�'U��]6%2��i45�O6��5����J6�vX��'�.�4���5�|�3I�61�^^Y6.�7;�����6��f5��5��W6�U��5е��O�Zk666�]�4�7�4!1v6�&7LY6�+�5r�u��X6� �4�z�5ē��滶�6!%6�r���R6Pv642�5'̄6�LB6�8����6�#6�. �pD���jR5x%�]!7�#����S6�'׵�W�4��7LP&�o%�d���T�����M��6AT6�ӂ4��ȶ�h�6���5�b��F��U\6ȡs4q�|5d�G5x[v��3�� �5�(�&�׃�4~��l���m��4�n46J5`�f�n����5o76�d86
s��T���vp6�M���E5BVön������$�d�Zp�5�M���Y��RX�N	�5յ�C+��c6c����5�p�E 5��6Z�5�?�\P�3"���b�嶿�;6R�������9���<�%������666-I��,�6���6�ﷶ��I��Cص[�6��#6t�5�S��D6���5��J����5�h6K͏��4W�J��.�l5=5��=6'����16��[� ��3~9Ǵ;������,U6�5�!6e8��{���0�6��6;�8�4_�/�)��4�U5�Q�RD6�L�4�A14�<���*��55�n���c/��%���<5Ǝ�5I��4 s����6"�5�
T�]}��{K=�M���|�6p�����a6*#>6�����5t%L6�.#6�E���6r��5�S����6}�+ku5y�P�x7�4CI��c�g6�d+��ض�b���c��q�4�F���*���i��Ѷ��L����5�}��}-�5=��?ᐶ��5�P������nw��`6����x6[�4���6��@�����ɵ��Ե_�+6qi?����'s�$s3$�Y5L;�5�<�����b��Oi!7l6��������0����%	6 ��������W��L߳�˶��$���6Ѕ:����n��u�$�8�,6nm�5�9�����5fy�g5`�e�|�F���6Q0a���w6��ԴR�ʵ�sI5��m�8��5Xc7��T5�yߵ��<6��\6D��Pb�4�����#?���6Sћ�d	�5��5=�=�6H/u6��	�ph�5�҃�^�S6 V>��ཱུc��Hp4���ڳ4�ĵ�7�6������h6��˵ ���$A��HX�/�� �3�4����G������K���5��6�ڀ�i=������b�����Qȵ�3����6���6^�T6�~)�����u㵻I�6�"o7��L릵f��=�5�6���P���*ڀ6o6�6N36�< ��"Եh 6�*�r�-6b~�6p+���4e�6'���>�[�`;��Z'��hp��1ѵ����:%������+6�c66͖���ƴ��´�� �?{���yc��S@4����be6�ε2�)6�J�5��P�~���i��6	��rڔ�@ q�0�86�մ���ҵ
��6H^6�O600�6Bh쵛��46�ݯ�<]26zn��:)�L�˵�M~6e6���r���>;��'\6<�5�A�؋6��$6�o5Nж ɠ3��*�x�N5.��5`a,3�1��&6M�U6	�;���'6D��5˸�6Z}��1q���6fl;6^�"�v�6ɐ�64ۏ�,�E��vx6z/�4}�5��B��UD��.A5��J^5 �n6=6t{�mQ�4N�Ե�|=6|jB6�?�6�F86�l]4[("�.��6F�6$�6tv��;5�7�6ĵT�.6��g6�3�'л6|�5�浵�o��>�V6���60����5S�G6@���A#4����~Hʹ�a�D�	���5NEa6�I�60W��/�5z 736�;4��5��ζ1I26`�B5�*�6pӵ,4���$���`6\�!�@��3�H6�9�p*@�f6�5��6���6fN6��C5�.r���Զx"�5���4�5��������7�ʴ���<*6��ȵ�026���4�z��4�%5���6����37�U��@~�d7-r6����� w�2��6p��6fz䶚��5�ʶ�����,�����4;�6�A�6�d16�E}5�K���Yx��w����57��x
7����5C����(�G'͵x��6��Ƶ������7��@Qf3 l���S6�E�5���4x����6(/��e8��x�6�l���� ��=�6pxK7L�g�\#Z6����u����@�7��eԶ|��̭���r�\׳6�C���|��V$5t��6s˘5`Og6�m6TrQ��p����?Y�6����zu�@\���b�ʖ���:��0��p��+`��uI)6���"��2�5\�]6�	�6h!� <ɴ��7��t�^�U� _��Z;6�>,6�/5���}��V��l�f7�=���Rr�����'27���DPn6~�o6�Ӽ���3~6ا�� �����5@�`��\���C�6�e�6���6LE�6J=�6~.6��B�`�5���4��D��4vp%7��W�>O�6U�6�5��+������ߵ���4T�)�h��5����#ڶ¥��zM�5��6�:��>�6�6�F�5��75o:	���6�fG����6�Zɵ�4���<+��yR���U=��A�4,���hJ�{��5��6(�A4)�Y�@�H�@�6�����6�	W���9��b��r 76�7�6�~��F	涻�68'�6V�5D"�xQϵzZ��H�i���6��K�Gܮ�h8�5��/6	��6�	���A�6�d�6Y&�6h�J������Q}5^�����6jW46tH��ܭ��ی6c*���9��S���_�Fc�5�\���Z�
J�6J^�6�ʎ���7�y��L�5�7��޶�d16�x�5`�'� :���5�2��i(�J^]�ڲ�6��6$�S����6��O�19̶�Ec5�I��e؇6>S|�"!ѵ:y#6�)x6�.��v*��9�r5�5h� �����5U7��6�H�R�=��6�Yf5��T�=�+.6��b����05LH6�<7�Y쬶5�g6�4�6����v]�50Л�NE ��+�<<G�Jʄ�PL"�ZA`6��O66)�X8����6��(c����6�N �m&�����7�����$Υ5ߘ6(������Sa����36�����
6@��4z;67��TY��ֵ�4o6�76�D��z�� �6`Q��k����6���\>Y��aܶZ,X�J���������㶦=6��5��5d�x�ͫ ��v6l_[4��a6)ǵؒ�6�5F�i�b�5a�5�µ�x������"Z�)꠵$����6��"3�1��<��g��5�\Y�S�b6�o�b�6<�7��HS�(������[�5����6M���>	��_6�v"54�O6��5��~��.3��
6�j+5Q޵���R*�*UZ���6��5��F5��I6.����t5�i�5�xb5�++5� 6L�6�1��m519M6e>7��:���7�(�4��m6�g�5n����m����4.�]6�J���f�5�˵�6�a4!_�6�.6���5�����Z���δ}�"�PD�5߃60�4_!�4
�ٶ��n�һP��K�0��3ĝC��5�΂6�6\X5�ʿ4��E6rN^���6�8G5�^�4s>�(��5�5PE�����{2�5�s�5`�-5,⤶��6�q,��p�����L�6�1-��r�5����u����ĕ�����6������5 ��
��6��7XA�4�������m���G愵�m�� �3���H^7w)�5�F6�6����������6���b$���@�6jD�5uN�5Kص�36�W�6!�:68A�3j�5l�6�Ă��! �}k6F6�횶���@��B+�5eĶ���5��_�1�5��:�;6�J ����5:�06��g�"�5�@6�,���cX�}�6���6N�5�/�%(	7�e�5\��6EM��>����,6��`�$E6XDW6��+2��6rRJ6�Zq69�5�V��6Q�L�g�6��j�Pל��I�P�����>6E����+7�7����4s��6�Y�6qɵ�x�6!p5�\��*�6�Y�5~�`�`6���V����zW�6t�͵7/�6�yh�Jh6�HY64T�6�?,��H����+5���@�X3��6|6k#���u6�,��l6vd����j5�<����+67�D�4�i�6��6z���]5^}�qPʵPtO�#��5�{6 �5l���P�6ݛ�5�}���뜶� 6��5 `��meW6�-���5��6١��C��, 6�̉�\��4����2�6�(0�v����l9��j6�0b6W�h�Q��6oކ�`lϕ6��6 %���[6��8�KfY��)6r䞴\�6O</6�4�w���s�5`��3��6��>6	ϵv=���0?��r�F�6<�e�pr��\l16�SQ6�6��V5�%�4�N;��?j�eT�B�
61 �*Et5��6 �T��vG��5ֆ5��5^�6���4.Z�p:�L����&x���$��|��|v?6������5�����5��w6fs����6���4p�36&�Ĵ`8��Ѽ5eM6���v�B>O�ә�����Y=�$	6�j�6�5�
��.S6�K3��d-�`g,����7��@D�D�6��25�`�5��6)�����5,�86?,E���S�H?�6�ۼ6�G�6�_	�#an7���6#�6��7�e�6�H6�6`�7�f��&M-7%eе]��5�`7
�	5[da�dʴ6H'�����x������x�+����5�=5�\µ-��6xb5 d��6Dy����5bc�5]�5:��6a�6��2��Ͷ$W=6`��3�w��j��6/����W6�X�6#��5D{���oZ7(CȵjD���赺�y6���Ӈ�L���yǵT�ߵJ!M���5TU��~m5h��Zyϵ�q3&�"5 (4����6�]�4\� ��
�Y`�6�T=6b����Q�5 ��4��5�����5�3�� Fd��x<�u	��/���ޜ4x=��~��4A�6�6�SG��u�6,��6+���v65j��5v����U5�N6��6���6|F\5�(�5H[6Zp�6pD���i6��Z3�tӵ j�5P^6��G6�K�'���5��5�.T�����M5�Am��M�p�25�-赦07���6PAs�P��4�H�00\6LT15J�t6�Y��|��5d�6sԚ����8��5��ȶY�=�?����6RW:6L6��`6dj��L��|���/6D�4W@�5�Kյ�bJ�DoI��d6�f5��4�Je6*#24^��!�3x�����5���s����8����95QT7U3�(�n56V-6������3��������6Lp6�`��, ҵ�j�4xZ���F�5���B���$$ �h�Q�M� 6�bӵR66}��6
f6J@?��u��S"6��6�%��v	!����6����;��)�5���5��Q���5��f��o0��l6�u����5�:=�N˼4�-6�M��= _6� 7��b3kH6.��5�׶z�:501�5�Wɵ`�:� �1Z=8�$�3v��R�e62u��Ɉ�6���59	����6����.A��$�6<1M��:��9*�ʄX��:6V42@.�HGT5��^�(�6��6��6�Kn�&/9�`���굱�5A�66`�]��i��B>6�5͵��&50�5�-������i�5�?��O֜����lZ�H�K�̬66����9�5��4ާ͵�4 �8ݵ����J�6`�����Z6)6.�ϧl5w��B6���y��� 0�0ֽ4��6xK���L6Z�6�����?7����5E�Ѷ���5W������d*����b3�5����x�5`
�5�]�d���T'�8綩t�6=�E���X�X1����6я5?�׵�ְ6#쐶b�
6dz�4xa	��j6�@��	��(�6X.60-�	��z07��6n�6f�ŵ��`�秠6��<�6�A�4�ʧ�@�(36M]�Tn�5�G��c#߶h]ص�
�x��@X�6�/Q6�Q����50?ض�l+$��3�����f�6�����68�5�W6fet��L��B'7x+s6�� 62O����6,�A6䁼6�m�6�Ͷ Y�X6ޔe�4�.z�5�AC5Y��6�j"��ص8R�S���m'��6Q5��1]�5��[��z5�|K��;����5n�7��l��4h����u�5/���ι��{N6L79���6�����cG7vA�5$�7��ɵ�^��ԣi5=����7ԥ}6���S���D�6��ܶ,�36��6.B�z�5+ ����5��06�Cu6Lw��]�60ܵ��6z77�AֵK����hi5~;t������6�ν6�m%���������}�6㩵�`�6]g�B="6WX6nx36̺�Keض8����:7 �i6����u3�6�6�E76�Z���5bD�5R>��A6�MI�
�:6��Ķ�P/7��ڶ0bӵ<�N�{��N������r{4&���v�6�E�q��6�w��rB6�}r6�l���}��H6�U���P����`6�I4�83�w�\q;���69����6� l�226��b�5����
1������]�6��04����C���!�h�96�R-��\U��^
�N)�kŶ�v�63�6�73Y6��:��1�5w�+���ȶx�˴ ��6?Ŷ�lE�A�^6�i�5%��-�\5R����8L�]�X6�L>�5�P�z�s4~��5�W�#�I6	�����H��T&���7�G6@�9��{:�<I䴆��~�!6�4�*��L?�5H@)5��G��ؐ��j��4-5@C 4�er6N2���_��60�h�$>�5�x��#�l6J��6�F5�����%4ϓN6�np6E�o6�d�5��K6�/r6����a1�ҕ��^��6�̌6m]%6��I��-ǵ@��41�P6h15�1��5+6x�6��
7,";�u����K�4V��6|13���k�t���x94�j���5F�w�f�Ķ��,6���6�fw��5�o6��6�B6t�2�k0��a�60�?���T	�ȓ�6 �63�a�44�D6]�6�]����j��=f���;6�J5�5����6�5�?�5X�2�
�R6"�d6N 76<�E6��0���a�V6hC�4d�6�9�5��s4��������2ٶ�� �β�䊶�G6Ng>��\��~�㴆�����4CΞ5�����w���������&��@�����������5�t|����d�@�x�6xTb6�=����]�&���8��5(xM5�~���1/6�r_5��6���4 o�4ǰ6ҠR7*���8>#5��5�֚�R��61u6�ef��h�6 k6M�h�2�� �ZtM��mF6���5���42�Q5'��r�����~�5�����'���56�R����d5S�6
���������r���%/�5��*�V�{��tX��v�J^���n53,/��80�Fui��dB��+7&�ʶ NT����B�p=6y��6��5Q8y��ң� �S��s��t�L6��6Z�:6/�ʵF�5�I-6���-Y��
�Ѷ|�	6�N�6n����5z1R�0�4���f�7�ڶ�g¶�]T6�')6XѰ6�����Z6��R9����y����6|j5����v�66�X�4N67���6�7d6���4dSW6�+	� �ҶLp@6��+�l_�6�&M6ਃ3D$6N�5;S6��$���6�tx6�ۨ6@�5n�9�P͠��=5��*��P�"5N�εԇ����D�=�6��="H6�g6N��6a�55k�� �3��3����705ă 6�o(6�M��*����6�S4��s5$��Rw��8E�4�[��d�ĴB{<6<�z�.�����4�?N6ȏ���	���>�6��J�$8�4�x�ZZo�,��6i�W6��6����<�3�T�5)���n�$�5��6�iݶ�f6�$���ߖ��2L6̎���N6�&�6řD�@��3��6��z5��4��\6^���h8��'ҵ��~5�95�����=5j7�J;�6c���P�55����R6޵68�5���04�6��������V�;��Ck�w�6�Bյ�6,	�5)�'�vA(�r�#�5��4�zʵ�
4ߺ@�}�2�PƵ�86 ����Oq��sѴs��6���V���cM6�DX6ώF6�Q�*w6�!�4��5�6�Z��(ؔ6���6��5�{6��6t6�q6��5�(�6`�5�P��k6��k4�9�ǁ�Z6�ޜ6Vѵ~�w�����HS��[���}'��N�3@?7�?s�"�6zrZ��G"�@6��G���ؔ�5i��4X745�����^�5� ����4�ZI�8;a�
�6P�^5�5��6 �@�ҟ>6�6��p�3��5��'5+d!5n��5���%�6��߶ ?�G��ݼ�5�O�� �3�Z4:����㤵J}�5�G6�b�6D�
6��Z5@nM5xko6n>��P�l4����r�s��b�2��'3h���Z�6n�ɶ�ݛ4��6�hX�
3�5X@������pf6 Kl5�r��E'��Ҧ� �1u�"��X6��$�}5���,Ó6A�G5��ƴ��O6 ?ʴ��d6j�5(5��31{�6v����zA�5�:��B
6��ǵ�e���6�B~3��f��3�6n"��h,j4�<���5�a�r9@6���������)�4���6�ق4�@]5���H
����h~���D6��6���]G�65��\9�� ��3i�5`U
�������\�5�Ub�*�D������������X�H�eP�����m�5k� ��� Tt4E���,6��=�l��p��;5��޵Y�@6�� 6,�
6:�6~4���	7�O��D����z��&6(7e5H��6P��3�,,6r����̂5L�6(������5��5N��5�H�6�q���*R5���6C8[6�c_6�6�w�r"6��7R��5N)��Bm���Z6�P^���K6(M�6��93̒�����5	w&�^�,6�`޶A
6��6�'�5�"Z� \w���I6��4`����"�t�k:���7J����ڬ5�z��ru�<H6{0��P�T�ٴ�=S68R6�Tݴ�߶�����U�4i�j�۶&�)7r�]�����zO4|杴BI6��i��Uڵ�y��e6mu�6l��>�7>��@N�66{�6���ܬ�!7ZQ�6'��5�RS��*��:����6:=���Ѷ��6��5G"W�E��M��66��T��\8r�.&�6�����7��7v֗��x�̯��t�w�r�M��{,6�^	6=n���A�6��p��}��:�5J)ٶ:Զ��6����ko64S6��_��'��L<�6���n�B��O44��=5�6��6��7������3r�e6��3<᮶n�5�'6������5���3���5�u�6}������]�6P2Z6�2�X	5�
"�F�%�$���l�6,���96y���0%�|~7T���0����6��4���l6<YT6�3)�v�����5^�o6X��A����5t�P����9$�5��J�X�6��-�U{�6Lu5�%͵��6p�!6�G�5*��`����?�3��\�77� �����66�G6�.7�܊6^��p�$4�Ŷ���6Zeg���>5�7x6ݞ����#6�iB5�?q5�e����������"\�HW�6�l����!���7薶���4n�R6(Y��1�6�x�ˌ�xNQ5Bֆ5H�5`�4��s6O֠�Y	�����6�,6Ŕ�6�Q�6�x�5�xٶE�6
��3�؟���6!�~���6��6wx���O
6�;"���)6�D|��OK����vw-�F��5�"ĳ�v�6(G�LnI�R��6"�6�yS6@G6��5�,%�5�6�TY4�Q48�5G�˵���N�6���7��6����㥳�ba6�r6EL��8�ӵ������i�螶5��Y6�ߵ5k���NB6 lϵ���Ō�����9��j�ֵ�_6N5:6���6ô5��5:6F�u���c6�|�
����.6)5�)����6C�F��Y�5��5�8 6�[�4Za��І���6qt����6�Y��f��5�Z6@U�Ӿ�4��W5��6f��6����o�~��5I�<6�z6��ǵ�(�t×5�r5(L6:~a���6b�5�2е ��4�Ҩ6}#)6,5s�[a�4u���!��6�*|���5%�5o�\��z��U��5����p�6��5��3 �p�a5}�6�6ۥ�52W�5��յ΀]6q^���S��lf6���4U�p5]�nƓ��e54&�4^�6�=5Jy1�j6��>C�5b6�Ү�,Y06��M�OG6�g�5�!R5�/��$��4[y��*#����6b�36�x� �3�| 4".p��K�5��5wG���-���*��L�4`�+��J� 6�M#����"D�5�~4�]�5B.)5����/{�6TB���zڵj�{6`��3B:�6��5��l6t���b赚�B�6}�,6W�6���4�
�6n�68PҵB��6��64ŵR�*5�n�5�g3��6rD8���G6���6�
�Wd����5P�6�7)�I����6���j�6J�'6�&j6� 6��5��B�76^�+��
E�ad6(3B6f6��출�O��⳵��v5�2h���/6�創pf�5-~6�(6�٫�8O67�W6��"� ���4֙�@���H��#�4P}�5L#�5g��N��5"F6���]9�<=�5س4mT4/_��=	���!6N���T<�����軄6�L6���"}y5�kJ�s=���$���G56	I5�,���!�,5��:�^��R�5�⎴$4Lۭ���� �VwN��-ɵ*��4�?6*V���� �Ry'�F����e16�^��w26@��4�Y��p�54i$���5 h�3����^)6,)6�:�"�5ZG5%1�5B���{<�Y�Q���5Fa}���@6:��5P�۳U�Ҵ�M4�9�5t|	�DO6����n�R5Z���u056r�5Xܬ5<�5�@6���˵h�?�� b��4x�	5���5���ʟ3���5Зݳ�<6/�]6�H5�&�4�����5�F󴺭(����5:e����5��\�m4��m5
|86T��4������i�*�6�6�5ȿE4ۢ�~�����T�׵������5 �a��s��$Z��,5�l5����k �$�r���fm�4b� 6�z�4"т5�>˵�V�5D,7��96���;D� ��4ɏ?5�/W6���5 ���֘5�r?3F��5P�B6�ƽ��	���&c2$��4/x5���������H5j6��3z���L��oʹ�*�� �5�56�3���5�Y96 ��5��b6���5��4�3w����ĵ�θ4;��0�6�s"6�3&�܃5���5HP��s,6]�5��4���5��J�<5���w6�iq3�*���f5Q� �:��58�,5��5�͵�<�5z�6�˴�ŵ��&5�$�:벀R����4>�4^��5��	5(<4ŕ#6^��o 6y��5���5JY;���45��!6I��5��B��g;3G8����52��4���?�4�>������6m?:5�5n�b�ު���5@4m���l6Ub�5п�4M�]6���4rq4/=�5:ӹ5dH�5�	϶�q8�\�6*'ϵFE��F6>sG�>26L�'6�����6�E5�s��X*4�;2�6 *94	Ƕ��5#6N����8P���5{6=�6�!�6�n{�yt���Ѵ6u���)�.�^��4ʕ6�҈���5&&�6 3Y4 f��
��5u{l6i�p�2��5(ٚ�J����6�.�EJ\�)D6ޛﶔ�_6s�ܶ�[�5�l������u��O��-����'��@=�6��P6����V�]�F9�����4v�(5[���?��������5>�е��p��<�Y�6�Wȵ@�e6�}51v55�`2���6f��4��˵r�3����}{6�~ֵJ���r�3�\�q�ȵ*:j64�5��c�6�X���ɵ<�y�|���i*�,��l��5�hg55e˵y¥6��5U06wȉ���S��u��k3����Pp��� :�����BtM5
�e��bi�8��4�&m4�s]��2)�����s$6�լ55Ķ^d6��46��$�s��5��3\c�5ظ6� ���5W�\68�����%3����(6b�G6�6�6ֶk� A�5`��5�y���ʵ_�4~2'����5ZN6y�5�DB6,E���5�~���N6��6�y�:�Y���)���i�`�����6�(J�C��5��&��|�6@O��T�5�5���4���6&�u��6{�5��z6Pa4��:��{6"�5�����L5С
5����o�6L�_5��G��LH6n�S���)��8W6'���8c���P���7����5T`1���6�G� 	6I�ζ`.6*Z	�
��5T���2�S�{S�N�/�P�'��;�4�2���\���z6p�L����4
�58�������������5G���C��
5�+5�s�6�2ൎ�6��5���'5<K�5[-���5 zV48��5��5"��5e�6��h�/���d�ĳʶH4Z
�D����3H6��5`R"4���5i�߶e>c6`�ȶJ弶�gg5p���9�6@Iг"�5^\x�����L�9�`����j���\6B�,�)��56����@��v6��50^�4��0���6��Q��l�4�f���U�4$H�6tR���H�5@�P42�_��Kp6p��5���5N�06`��3��)58��6��2��=�6IV���g�X�}��(f�:s�5?�﵍�6 ��8n�5e�6bɬ���4v����6�E150I�4���6D��ʚ86[��6��>��� �D�4߳��QZ0���_�� ���!:7`� 4PD�4�k�n��5,�6��5�P��Tؑ���6� ��B�L��1[�J�r6�%�6�I)�p�l5X�Vp6�򐶒�e6�
��5���y�6��~5`⺳��nk���%�6e��6z���{��,4���4 5
WL6�Ҷ�D�4[6��6�
��A����Y6�P�Ȍ���-5B���<�5�%d��0M����60:�F6���X�p���������@��3ʆ6Δ�5 ���`��!�ⵜ8�6�n66�ͬ�e듶��{��i�v�_��z,6П���X���/6��P5�T���Q���g6�[[�PUK7�X��J˶� >�$9�5@�#6�Z���O6�k�4�L����6�E6�����5�"�5U=p6��x�\�Ӷ���q��r%�b�ѶZ����e�5�O�6@�����Ե2$�6eJ�������M��"����6q�H� Ve4��S��2b�bV6�bf�Y	�6$!���9��k7�O�����6��w��ep6���5��6��6�K16"T$6�56�S37��h7�`6�.�X"L�,,����=���7�\�6�ז�*�6��H6w�1�� 7����a��5���U�7X6��6Y�16����CT5Γ6 �4���5V�+6�S�6 ����ɵS��6�Z��#5
ݭ��3^�ᶃX�6m>��G� �m��6�?7-�5&�76�6�f���j�6�0P6������4��6��,6!r�6١6�s�6��������ڵ��X�"ܵ��:6\u5r��X/72|f�y�5ݺ�6bS�5tu�5q>�ʒ�46\�����6l����ٺ��^�686<�[�/6>3�6�2C6�h7g_q�_ɴ��
6�R��6z		�@�6Z�5�� 7R痵��378�T4� 66l�7s�޵_؛��t5�JR�����5^�5��G6���5q���|��5�#��G_E6�G�6����6��͵➆�i5�m��&<�R�6J✵,j�5�=�4�,���n�����4���4�[����O��l4�+�6/]x���l��hq�N%X������5D�7Z����*�4$�161	��9�6܍�6p��6��ڶʿ5�ᓵ�݀���|��"�k�����B��6��	�v�-5�"�����n���q+h5�Ŷ~����&6�oδ�6��J�)�6Z=M5����������6�յa�����ߵ<ke�΁��첵�I�5���6�T
��	6���6:Jy6����y��6����)H)�����3��V��gE6G>���H��G��6%�d���G66�6B:7�A�6-��6����C�?G��݄�6��Եx���	7;㶜����2/���ѵ3|6��5XG"��L��N6;��6������7��`6�&�5�2x�q�P�.w6�"��������X5 J��[C6�SO6r�M���:�6r_�Ka��z�\���3�)�5��v�*�ߵ���n6_V��6ܵ>�P��fݶ�|Q�v_�5ظ�4� 6���5�8C6Dۣ������𛵋�6%�6M}��i,�(�5iu�����*����Sĵ�u�-2;6Cs�2��5��C��
�5��U6C	ݵT�5�"絇�0�
�l���o�"��4n��5�t����5��4�016ГD���6�5���5kW36c�65�i&6D�ʵ�,�6Έ��<�7�o-��甴1e��'�5�B#7`�#5@_���"��9�6B���S�Z6^s6XV�5Ẍ6"�6��36�7�5��85`�e��k6��C6T��R�6H�v5l�k5v�5?�5���*����0�6��/�p�ʴ<x4i��p��4�:��c�`�;4�6�a�6���s�@H#����5d s5X&�:a� �7�-��4
ҫ���6�$�6���6Ѿ6�����56d~*��P����5{K����\�6p�A��6�
7R)�H���y���6�
7d��5�p�� 8S���o������(!5��F6�#���/5(�6�:��N�5�|6aG�����ľ̶�X�6�Y-�`)�3=3��.��5�iR� ����DM��\�5f�u�8`$��A4�	V6ƨT�z1��H��5��6��6>�	6����5�X%^5�r4��'6��50�	7-ִI�6��6`�͵\�T��5��D��Q�s"� �ƴ(�6L��6��5k>�64�z��z(6�;6$[���|45qG�5�VC5�e�6�b�������7K��60Vc5���5~�޵�[���5���#85����p9B5�l�5 G!4�6(���7��p��4՛�6���5�:�5KG5��Q�u,��c���!��m�Z��;�k6_q�x�
�P��6hf@6�Lr5  7���Y7$�%��E��!ض$�5}�}6d�7���:�Tx�5>���2p=�@��5�ڇ��L��b��"��6@6@���M���
6��6� �����Rx5��6�6�f6�&����ҴL���:���6�V��"6x�´>6{�l��6GbJ�>7dk�lQ6������5��2�t��6�AT6W85��#�|�Ŵz�>�25�l2��)���V6*���V�D5�OI���	��P��Ӽ6�aX5�����5lg�5Q]{5��"6Nq� I94��	���5��Ƶ�7�Pn~6bn�l9?�Z�������'E5d6�P���Kϴq����D5���6hGq5?:�5����2��6��v6��4�b5�E:��Nc6�{a6����6p���(�4p�6xLx5&����6oյl�Q��Nf6�R:��86 ���8����v5`0u4l 5��6va5��B�D̵������tԣ���4�����䵒\�6?&67�}y5�*-�&G�^��+6�TW60{R����5R�/�У�6���]�6�9)5񌃶Aק�l��6�)���m16�~���v�y����5X^�5���5�x6ؿ�pk�6P(���횵�Gy��~�4�j�6��k�6��4�b�4ga7^g�5�ŵ⮧���X��,��X�^G�5�6$�����6��/�p�ʴ��D��(���Y5�Ǆ5~�5�,�6O�5m�M6�%5�c��E5U�5ӊ��P����6d�U6��5��z���B��yy��)6fLw���3 亴oF�� �64ZO��p6LW�3P2��c6j��5r�;5�	�*����'�$;6��^6 �_6�����ޔ��Ut6`5"
�5�؅5��x���6��5�L/�p_ǳS6F:�5�xĵ�P6����1-6z��5��6A��5���j�36�е�Y���س�@���;>��&�Եn�۵�,&��)5��#6P��6Hr-6RO�t��6�f����5

�5`�l�]NC64q6ʤ���J�52N{5^�ε��V6E�ߵk��4(�ش�:&76�)�,��5dB�TV6���6\���Vv���M�|�V6�쒳Y=׶��6���n:Ӵ���5,G+�2�X6�e�h�U�rd}�lGе��6� �6~z5�Hz�iyZ��s16pv�5��6��h3"ϵ��S�5�6�R{�ף�Y��l� �B16zA����5�$�6�U���G6��H�
/�6�&�� 2�4�"6��T��o5��B5�'ﴰ�v�CG�hC_�L���6�t�5���\�5I<#�4��`�%7����^��ɨ�l"�6T��6 ������4�&`6�ߑ5�J����5��6�H6������!��FyN��E�4�
�� �6��7�27�X.�"$�6�H)�d�o5���z9%70�#��t4e�n5Ӳ��pP�е��#6�3+:3�����\�6$X8�b�J6�k����+6�ȵ5�.o7g5J6�����P�6����V���Lr�68�����6�p�4�46,��6n��5����6X���k覶b#��}
�ѠU���A7���6�95�=X�|�6���5#7b�Ƕ(�Q���ѵ@IM����_8���6hh�6��53�6F�����,b�b�5�n�6�.����5:�Զ�� 5�)"�`��2rk968`�6�ߴ�U���\� q-��#�� �m6*�6�t6��Ƕ7ε.;�6����(�6�̯�5`v�NB����K�2�j6���6 �S	d6h����/k5�1��d�A��a4�eM���,��@�6�,�����ĸA6�W6�5	7馴k�G��P�5��N��V�6��O6�����I5�6�n��$d60[5��K�g��544}��J5� �6��5���5<��X��Ҿq5�7���=6se���i�6���33���F�6�<�6���6�f���	��gF6V[�5x��I�<6��5���6$M*6��.��C0�����}Dh6��m�?�6R��5�^6���5iK���z6,�a��6����t���5��6>�U�����ʵ��7v��6��ڵR����)6+!5�ӵ��X5%:"6���4�%��E̾6V�z�O��6c��h����-4�r#�=�6PYk6�65\
�@ґ��k(����4?F����5
��5��5�5\̢5UvR�<��6��6�Q�6�L&�x������6��5���5��Ŵ���6�^L6�U6�s��%?��o�5^�4�D���U6L\|�#;���p!���󵨧�4P>��f�6�k�����5��6�� ��l�5���;i�5�77`&�4���6y���CP6�G6 0��>86|ڀ6��647�64(��s52�#6 �v2ǚ��yI6x�t68��6)�^���`�z5��۵+�1l����p�J� ��kb�5࿕��j6�?�5�:06�N�63؆6��Ҵl����6�gY���5�B5	�;�j6��6j���|����0������ 5g(�5<�z�<i15_|��&���2����69����8��<y�6�x��l����6ȃ��=���Q6�1��\��&4�5$x6\��4�s�����`��f,е $޲�T���6K3��@�.4�< 6j��5��h�6F����6 v���4����ޞk6�;�5�,�����8�x5)6�c��26/0��6
¶�
���<6�b�6�Gp6;�5Ȫ�6�u�l&���5.����s�6`�P6A����5VGk6덿�q��6�5�!��f~����2H*�5�}J6�.�4L/5�I�=�5��b5.�,��|*����4q��+J~6�o��`	F6��E6��6��v�<H���ִG+5�����G6��(6~�8�/\%���5V�'5|ѷ5���5��ԓ̶$Ρ63ﵢY65�2�e�;����5�f���t6�r*��0�6��5 N�3��q���F6b��6��{��@����6�Ă��PԶk������5&�6o�F��Y�5/�j��U�xO#5Qdඕ.���,6@җ6�$���*�M�5#��6
�7C�J� �,s�6�Q6�[>5�����t�6��-�W5\-f6�%��8��5�j(� ߮5�05Pn�6<	��6���Ц���}�p�84l2x�e¶���6�ӏ6k̂64����O�6�X�6E�6�W�ĵ|Y�T��`�5�'��0���A��w��)ݵi؟���	5a�ѵ�&��s4�P���OS6�wT5 �=����5��m4��Z�x2��E����ݵf���!Q����t��$6�3�6ld�6L�l5��t5&!�53<6�� 5�<6��}��h6>��4oɴ���T~���ԕ���ڵb0k5_��CU6.@�6dP$6M�6-Z"���p'2so��~*�+���E���\�6�$�D@���	#6 g,��I1���6/�X6�5�5�ڳE�o6~�6BS�6$�ŵز�79+7ث�4�"-�>����i��	�60-��E���&+�Z�w�� m�6��!6���5�!V�K`f6 �I�f�m���Ŷ������f��ݤ�<t8�%:��!!Ӷ� �˓˵n~j6�h35{�5]UV6t��6�q���Z��u5eU�5燶���5\�k��w!�5��5�a(6��/5�^�����m<v��v��+2��c�5��4J�4q��6|k61b����6�m�6�9�d(25bQP��5f)�6.Z6gX$�|�����z��/��U���'�J�F�>@��OV��N�5���3���6>X`6w�������b��4��5x���M9�6�`6�6&�6��Z6
(�5a�_5q�1��9��x��4�k�66��6��E6~Kb�/��5�/D���5,��5�aT�?5���?6�6>@�5b9ĴB_w�SZ5�66�b~�fZ[6�6�j�6z4.��XX��1�69��6�?,�-@�ԁڳ`Iy5 �5T��[��:��Ü��}�6LI�2_b6BgF6��J�f����l�ն�6������5R��R2)����5T�6�j�6���6�� 7>��6�`��i�y��� ��&�5�4]4�͵�l[5@���	66�tN�n���ᶥ�b�3+5 ��6kr'��J6���5�a6E6�5�/�5d=��T�m�^�$�f���`��4�OǶƎ�5(y�4�bm�ū�5Ȝ�5B��5
�ϵg�{���6,G/�lh�5rOk�<R6���Q9����7���1�!`*�ɪ�6]��6!�6���"絣���'ܟ6�����6�Ǵڌ��b��Hɵ�6ʱo�>#�`_K�/Hϵ��S5�Lʵ ؉����6�L�(��/N����6dFP5��;6 ��4Jh68�ò�4����a�@���<�*�\h�6B��6���5�߂�9�5 �)�Pεt�z�i�=5�� 6]�� __5�s�5���5���q�����"W5���6d��[5���58�W���l��U�6 ���X�5����bY�Nth6�
{�96�Եp�<��J����5��Q6�v<6 ����5��N�8��5X���rc��ϥ5�1�4�k6�-�4�wZ�3P�52���=�3`G?4���5;�6���3z��5��a���r(`6`�]�&����D�R-�5��56�_�P���2�5��5��&�lr��C5�2C���$�.5t��60ȅ��7���%��2��޷��!q�pr�5 �3t�;5�^���*�5�s�5@R��n���P	�t��5�g	6�6�*�5�2��S�5L�`���6>�h��9�$�#�@gE3��ζy@���u�5�:6\3�5��5i6�6�x�>��5_m��ԫ�5��A5�4%ȋ����6`�7���ҳ�L��>����F�߫󵀶�5���3@��3Fg�� ?�4`���k�����5�R
5&Ø5S����ֵ�j�5��?6R*����?6z�G�TC66�vB4�
j5�*����4 j 3|����~�@��4h�M�s������5B�6��|��i�6���v��I��4�
1�B}����5G��5���6X�b��b46�A	���5.��5��5��54I�����5G�5��>�0Rj4$ka�{�B6�R���5P7/5 �д���6�L�4�F5�<�5$�%���j�3X6�����?��&*6T��Q=�6��6�]�5���5$�6���>|6���5�N�5mo�5M~m6�w68�@�3 ������J6�;S� $a5<�鵆b\�66��6�25�o6�>��| Z�Xz"�GD�<����J\�1H$�!�5��m?6���9Lȶ#��5�WK��zN5��쵰.L��m����5���6 �F4� �5D5|���s����'5�{��݉��5L��� �˴�(o4J�M� ��J���i��I����v5�a�b9(6?YY5��L6 5̳8��4���[�6���6ȕ�5x�;5`�������/6�0�-�tp���X��d�5@�k�>0W�@h�4>X�6�z���Yo�tW6`75�Zݴk��5i�����5%�t6륶�<38���q����5LUf5uZT�<��5b7�5.�#��4S6�g�6|{�6�����(3L�Υ5f6ѕ�5�������(�5��J5��� '@4��\�� ���h]3YS6o6H槴6��6�վ5��K5Տ�Lͺ�5��e����2�])�!v� HC50,����� �m2z��5���5�8� Ru��6�15T�����5̲/��d5t�R6�ѣ����d�s��\5Jc�6"�o6��55��d�o^\�"�*�صZG��&�5�E��e#}5'�^6
��6xū5(��p��4�������@��|쇵�{S�:ʉ�x���Q�3�F=����5SO�5�J�6�"͵�	@6�壶��[��h5�v�x�y5�U6�; 6�L��DJ�ϕ�6;е��
6�L^��*�5�ŵd �祹6��5��#6���Eܓ����5�,�8�hٵ4nK6���8"6�i.6>��5���3m��������5�^V���� ޡ�B,%�I1�&��6��Ǵ�k�D�f5�5�����:4��c5�*����ڴp�%6��m5���6��76�P6A�5�i��q�36<5|��6(Ŧ68�v4�j�6��5��3��5�h�3���;�_�E�6pV�X�5Ӡ�5��e5/M6.0#6hXO�4�6PϘ5?�#5F��516�=P6�r¶�O��Kô�p�܌�5L�[5=���av6ː�4j&6ʣ�5V��6����X�5T��5�5֥�4��5�'�5��ݴ�5r5J� 6�`P���2� �ɳ�M\6�t��u�5Nt�6�9}�*1�5�Ų�/�-5*��5�C�5+��ԭL6Z%6������Y��y6��͵t��5��X��4�7��[���Z5n�R�X�׵����⟇6�4��`6�"��x_:�I�6�-E��]������5����Os{��U\�����1�u5�6�εr  6j�5+��f�5��W������K5�;6�o���C5�*�5܃��(s=4s*�5,�����h���(��5֦5�@V60K6q-�b�688���M4t['6����q52m6��4&�p��cb�B�ʶ�6��5��|���D68oo6�'��Skk�v��5L$�4��e��V6�p"��#���66E�6��h6 9����p���}�5H~5��v�%���Ph�N�͵N׷��q4~�W6��4,�?�N���M��ʵd����5Z��6+F�6�������6.�&6�� 6ڈ���ҵdk%6<�F��i�5�_	65��L&���T:6���5X� �T����a
��D���b!60O/4to4�8�3��!��e�^J�5@�v5�&M5��O5T�Y5�F�4"?��06��>�?���0k6�����5���i�5I���5b58���:��6�i�5^LڶI�H���+�F�i�&�a6В>4��>�@��6p�K3�������J6Co2�N�6��0� >6���!���6#�@��6�ϋ����fɣ5s�S�s 6�V6�f���'��b�����5�B�4�&F���KI��V$����J5�����L|5�8����5�Gn��5��,�W���50�~5{������Q��m�R�؅6��Te�6`j۴ .O� 6(P��5�m6�kE�\.�4�W� �6c�6+6P�P6Ei�/��E�3���L��5~� ��nd�g�k6�<%�@�14P!05�Q��	�5�0K� ���#v6��5L�˵�ɗ��k5,�5B<5�k6 �6�� 4�}�4�Y4�N�5;�h5&�ߵ��M�T��6 �5x������6����c@��ȶV�%�r�q6�Q�a`I7RT��-g׶� w��k� �C��k35�'��CZ����6�(���ε�A��6�k7|��6�[}6ú���/��H�kr	7�y��e&��
7f5��|��6lB5_ ������I6�5*7:&���t��R1�t� 7�^׶-���X�_5B+�5r
൸8�6 W>��ö�k]6H&��3}7�5����/6���*M7��z6�B���z;6$�6�`%�d�7�J5�=��v~׵{e�Ě�| �4����[6��5qм�p�6ɩ�6K��6Ѭ���ĶސZ���F�1�6$��6$��6QH��T�5�(�y��6ض�5j킶d��604 S̲Xϓ6`mW5��	7FL0�*�5�s�6��?4����ho!��r�5j��XTJ�%��&$�6�f�6P��5�M�6C�����68+�47W6����.�5��6K6u6n�6gǵ�0{U�ldG�����=6G�!���Y��s���	�6��G��	6��)6q-��Sp6�w���6�A6m7�¢�6 K�<�i�R��5u�4� I�LB�6t8ڵ<��m/�6�e��c%�T�f7��5H��5�"�9��s�6ދ5����M��h��69�7߉���� 6��L���6���3L�h�\�Y�ֈ�5��5ruK6;��Ơ��Hq�Lj�6>�ضJ�w�� {��%��+B5�ҵ��6h;��ʀ�6rs�5
��6�� 6�.�5Ρ��T�Z6��6�Ι4/Y=6�c~6�=���6�޽�ӌ�6�.7�I�6��6���68-��@豶@�6��%7��5^�46��6�w6H5u5Bf�6|J`6���6�:B�ΰ�5�?ڶ�Ɖ����6$_��h���NN7�Q���`����7�++�>��6p�5����~<G6��ѵ���5f�a٦���r���6�x����߶��t�x�v6X>��hv.����6D C��X�6�aD�����*��!��$��(*���6G66��o41�j6`_j6�s�6���.�5�����4��ܵ��.�R�n�Ķk6�6�6��4^���(	H����dW� 
����4bv�D�8�V17�?�ѶX¶1c��J�6<
7�=6��{�z�y;�6�:���F6D��5F���Ĝ�6�9�5��L5��5�50�dD)6��6B��40GU4Ͽ�6�-��֨��0�iP#6�ʵ^65��{6���5u6\�5�W��M#62i�������4�\��5dK�5V��6,*�=06�8���%c�|F�5;�:6�I��F}�'S(�\`$��,�6gv���6���^o:�m���_�57�����5H�i6�KN��E&�pc6lwz6��s�ԩ�6y&��a�6�J_52Y���i.�e�5��4<��V�6 �5Rf6ȿG4[����K6�[����6R����>d6Y�x��m��i�� �T1q1B6�� ��N��D�5�B��4���w6G�*5��^�6@Մ6DvI6CJ�4Ț�4&��lAŵ�]����_?�t���-�L5���6��e�t~E�v�ǵ�6��������������� 6�xݵ�/��ǔ3 �48���7�R�2A�5�[6�Ò6m�6��)5:+(��
�6(S��3$޶�뵟����6Q��59Q5��6C&M68%�j����E�6��g�4P���Q���C7����5��I�.�6��Qr�3�6h�ܶ�-�����ަ)�� ��v��H�SQ��0�6ƀr�b�m5�	�6�|��ʤ�64�?66�жY��}����������Y�PN�5�6X��ޣ5�T�4�r���õ0�75��x�;�6�+,���ƨ��6�6��5���@r�3�y|5�q�rA6�@������fa 6�IV���60�ŵ�a����	�������}�DA"���6?�Ƕ�p6Pv��56�>^���۴��Z�Ȱ�6pH\��5�u��6Yr�6�-6U˴����4�550����6��]����3��56:��5�6�c��n���p���l�6���#���	0 6�J_6D��4p��4Z���<����6�6��5�e�6�µ�Q!6P�0�4�6J��6B�&6%r6�:�@x6����Z�:��ʶ�(6��� ��4X��5L�f5��7��͵��M�d��5��Ŷ� ��Jhs6P��3/��~��~|#6HZ�6uA76d��5�.���3���4�%��no)��Xq��X6���� [մ�B�h�{$� �)�Ч6bpn6�R���r����d���aO��h6Pn]��Ȇ���������z�6�O6|0�5�Ӌ4��76�y^6w1�Ř6`EA6�:A6��5J�g� �d6��J6z⌵"�[�T��5>�6�춶�~���^����6z�ǵ5��&�7,�5<L�5�� ����d�J���.6{6�rX6}~�6���lZ6H��5��p6���x�e5F�6Y�6��µ�/�0����5&6�̉5@S�,]P6X3��o6�wq�@�#��JY5��6ob6wѶ��!�tꤵJ;�6�i%�����n�6(�6��:���5���$k��&������C	�"�6�!�:T����3#8����ǐ�� ��2���6��fZ��> ��$����}�6:VR�7��6 ��5��(5�I66��6��5$�1�P�"6¤���ȏ3@��4��T�')c6+(�6��v���[�`��4��6��P���"6�L�6]�۶D�������7ȵնt��5 �w4�Ǝ4kG,6���4N(69A77-B%6=
7�%�6�zж+�l�,��5���5Z^�����5:d�6�4�5����W����F�5H�n���w�ю6��4<�^b�5b^ض0$�3^g���6�;6�6l�b�,�6�O6�]��5�Q�5�����*5v�*�6 ����O�ꔆ��������ht�5(�	�ܩ�@�3���c��6�"��5>��60�}��'�6ַJ�LQ�6�Δ6(�6�D�6B�Z6L�O�3�6O]6J�6������5eq26 fM�y�ʵͶb��6>�,6�Zض@�D�G,L7�b���s�O946ݬ;�HiN���5�j��Y��6h�Z6��͵��ݴ{��Ԯ���6��5���>6�Sܶ�	���6(��5��5�+�6#6r"9��{�6L�5����o�6rC��ԙ�b,��T>�6�n5r�x6<�"�&�#6�@̨4J��6�j7��7q�s��Am5u��6�p�T��6.�(�\��5���5��5꾫6�a$689K5���5D�5�!6�[6�ꇵ�jj5Dee� �X4@[�.�6F�6���5�:6���}�06b ���S5ұ968�e�I6b6���5~����=d6�Ю6��%�{�!�\՟4*q5�Y�����r�57!������4	�69x�&*��P<�@�3�^��^�͵�b�5\�6^;�6��7�������6ȹ�4�q6GŶ��6"�������+��Q$6!�G6��ȶ�-{6���\ "��=���3w5�s�6�[)�8;K��D�6Z�(�6�A
�h�i5(�Ѷ��g��sƵC*j6�g�5�K��rV��w7�^̶��7ذu5��o6�D(�ה��0�6R� 7���a�68P�j�'77L��O�6 �g��l�5F�P7�9�6��D�k�ʶR�5���6�8j7^�������'6��86� -3���5�*��[)��`X6H;����`U�6��6s����7{�6��6,#H6���6�Յ���b6�<%4�ɶ@�?3����r�5''���q5lp�$x5�h.����6p%|�p��"¶kd&����5�����L�6>+6<����ڜ6�vJ�Jp5�M6����"#5l��4@�m� ׵G35$&&5H�"5�{�5��}��ε0(���tͶ.�����Q4$�@��L���a�5�Y走�>4$�M����5��7�D/�6>���Y���N�'6���xx�6B|��P�Ķ9&ҵ�I���6���J6` X6��}�6�g7�6�Y6Ǹh6��C3;p6� U4�(:���3� B�6��6��D�ş�܀3j��6�C5�-n6"�E�R�p6ڎ��fo�ڠ�6�6�,�"�4�P�-6�fN���6���5���Y�t#w6f��6�4¶� ��T7�O�5�m��>q� U�"d�6C@��s9�6r��5�o6��
v�5�P�{�?68�49�Z6���|l6A�V��k��pE��29���ȵ��C5X
�4��S�6@�3 o޴P�p5�����<��5��4(��8�\���/��a�?x[�,u�ʵ��>4��5�t]�VV�5�� �8���µV�����T�������^Xk6<PW6���`�4|J6��5 L���"-6pVV4�A5G����/��ݵ4&7-�!5�g6 �Nn���?g�(�45�4��H[/�{ᒶ tV4\���a�P��M��V�5����2屖r(��+�67��5t&ܵ�;���Z���6΃��)'5�R����62����-�4�T׵���Dͨ��Ș6}���Sg���!̶��w���5�q6�/5\�7������!�Xl�5ZC���:��&6��Ԍ��
?����5��7d��X�6,ȶ��6��66����"ٞ��
�DQ��ضd�O���S�<85X{�6!��>��65��^�06 +��(�!������(�;PڵY��0�}6�`^��N���õ���4F�4�H�|���ܟ�5�l�4��I6��s�nL5��\�8�6���5x��5V � ��5��<5g0�6�4 m4�w����4�B���v6�D`��~�5`�w6���5 o�5"���[���F׵���5�6��x�A��(�4*ʵ
����ԯ��	b�v�5Pk�nA�5�� �f�;66���j�5�f6��������n6j�㶰G@�`u�6|�X5
Z�6.�5����J6V�����w�1��6���6��U6L�5q�W6��6���h2ʵNhe6��\6@�<������z���Ŷ �������� ����4��@c���j��yy5o���J�϶*�66N-жUm62�N6[:���5�S�^���t:��|'����59A���?!7��\�
cŵ0�k5]��5E�Z6�jƵ>�86¢���M���5ŵ��6�@�6u&R�ŭ5��?4�\�6���6��6��D6�n58��4_;_6����F�5��6�W�n�^� 6\�G5`�O��ڶ8��O5�N��`&�HX�3F�'.?�J��5ֶ����cP5��6�XL��!�����Y�6���4HԜ6KQ@�8@z���@�H4����u���j6�h�5�;�`�+�N6T6�V�����6��T�vb6Զ,�_5�Ȳ�֮ⶬ��6|A}���`��S�6�l���0/��*�6��_�6��5l��5�(����h�Ⓥ�6�>��+�6�,�5p�4�o�0V�4��R��vI6:��6���5��5�s�5��,6��4{'��N��$y�5du|��k�5�DL5~\T6LPV��
�̓26`i�4�R7UM����6���!�ֶ�O_����6`�l�F_*�N���1nK6`�(�x���5֡��Lk5�S�5U�5|x.6������5pEI5�	N7��������ߋ�6ޤ�64y5⍵���4F�Zfd6iZ7|�*5�^�6��ȳ��f6&Hȵݼ�丆�7]6 ��5B
65Y��NC�Xw|5��6�df�����Vs��TF6�x(��ǵ=F6�,��^h5�:G4v6��$�q�	�6��5ȁ@6���f�x�^$n6��Եt)�� �O�j �<Z��li5l�K��]�5߽6�d'5��<6���2�۵^��6��6Q36W$6��Z6d1�5�����6Dm6�����D�<t)5�����˵�ͳ��;6�`7�y���p6��	68�6����o�>�!���zL��D�5vR�-�)�����*�ѵ_�5@��@̂3W\?6/������6�o���p7R��C��63g�6�g�66�ɜ3��E�6�7S�6p`�6� �6�m44�S5��X7W=(6>)��_7܏(6�
��o�O7��o��5�k6ϵ�6&����C6���6X��D�p��c�����ȱ6<1�6����KL��w�57*�54�x5��5�ƶ#��6��#�f�5�r�� a�4�&�5�@6/�5��,��� 6#6�����5�B˵A-]6c��I@6�v�8n�� �_5R����m�6[W��D����5)��6$���:����m�q��6r66��������ɵ2/��Ǯ�BA]�ģ�6_�6;�ƶh���@6��5b��KU��U67���6�-96bS��6�������6Ek����5��D6B�O6y^��p+Y�8<7�K�6�r���Y5�������!�]�bU���q�4F!6j ն�!����$6lP�����6,�p6b�4��>6@6���5��޶�_�jᵆ3�6��63;��8���L7�eȴ&+7YP׵��6o�5&1ֵ�Qж��5�k�6W���o�6�
D6jtf�J,7��6�=���(ڵ��i�G��A�^y�6��� ��b�6;��̏�����5��|6y�t7B�Ҷ�l� F����H5^��q�*`6��g�P� �{��6�;6\��4�q(5o��6�B���?7,�ڴ
А��c6����׶������wqL��,J�CZ�6Y�)5�6-6��5�i�� w�
��5v�{6�h����2�:�>�3O����V���1	�1��6��	�y�3�B���6 v��q� H:4�e~�۵굫R96��43q}6��1��5�*6���hn�����6!�&6�S6ך/�(3��i��5L� 6|��޿S��~T6��6�N��M#��g/6#o����5�DI����5$�p��*�3��N5XO�ފ5�6 ̅�om��*�26����~��5f��4�U��7�50r%��5��(�5^�5��a�t�5����|�4�^67&/6뉶��N�X����?5B:۵��6V�ĵP�H�b�]6t��Sz{�<#6�i��ꈴq���c��烵a����w��,`��~�5;w1��rö�����5���X6����9���>6vc�5V��5�i��X�2���5��5�ъ�D!G���.6����5"��5OR6 �05`���s5�46c^16w�/�@�ǳϫ6�ڣ5��5��5�̰4Y_&�7�5��t4��Ե���5��6�h1��(�6��:6r8��g�b6��Դ澞���ǵ�(�$~!�BT6_�����V��K浒쯵b��5*�m.w����5!��5<�p6 �3����m6 �r6H��4	Ӌ�"Z�ʛ{5,&���#>6��a���ڵ �E��y6b��DT����N��@[���N481�5ҳ�51�6|YZ���V�@₴��5 ��<UP5�y�4�n6a|5���5��y6��5�2��4X�60��4IX����(f����6��O���5P�5*k%�{��5Fd���5�?�55�̵$!�5L�06J���5�I�5��Y���ڴ�WM6�A_5�l(�8�6�35C�l6_�4L��4w ��$�XÍ5T&6}<�6�o�5�l�5�M�588;��e6ڹ�6\x86�DD��js5���53f+�8V�5,8�4����!�@6�6��)5��`6Al���)����4��k5��ʴpm�/�3�Т3�.:5F�6�vt6!�6�F;����� ���!���v5x#�5�����6@W�4�(6��5(7�5�MO5��е}x���]76������g��!���}6�I�2r����6�Ѹ���F4e���J6�5�y��Ҏk�&@�6��H��05�	K�����]ᵀC�4�Ѷ�o��&)�_U�6X�M�7��@��(<7���6���џ�6K5�,5�ӵv�������Q�6��z6ܣ�~�6���5�6�o[5�`$�z0�R�96�汶.�6�WQ6����h�5R�6�O��pI5ݤ�6 �3���lI��Q�6��]6����f 6Ԕ�h˴��2�P�����7DI6(��[��6p�/58%�6B�6ӼD7aS����ǵM䥶���6rnu6l{�3 ��1 �\4L���� �Hf��U��&�4��6�zJ6�T�6�.:�$b��Ȫ56e�6}��rj��Z�50��4˦+���5�讵��6B�6���� ���76 �յ_��6d�6�M���@6��6$Z>68��6@H"��(����4	*�ی|�9G�5 }�6(0�6��4�ܮ���˵ -���6�W4�y6d�/�������6���5� �6��!�B�/6e/ӵ�V�6����t*9��^����4���6ʆ6�Ͷ`N5w�x6�>�6�`7D���
����U6T�l�w�6Dȇ��{u5�o�6�Ķ��7�:k�A�6��;6��K6~���:27Ѐ�5���5� A4y�167��6�����M5վ�6~�����65܍��,�X��4��+6��7��5�����	6#�`W��36���L�|��6�q��WK��TN�B>�������6����F���o/����6��6��A�Ei�6w��6�Z̵�<6H�6w���P�;��6��f3�5�-5>�7�l�6��7d�-7��{6*��r��1�o6(��4.O���6�.{�@q���#>6#��6$���}��5��ڵ��!�5��6B��5Y�6)�������%6��v5�޾6��U56E���s��BJִX-��~'��v6�Z{6T��5�;S6���z�~5��jʹ��'6�>[4��5zu*6J���쐚4��5��84n��5J��5 *�5��ٵf�ĵ�546��C5K�G��-��ԗ6o��.V6��5>��5b�0��GصP�����N�7����26�'<6p�76����GMi�'�6L<
5Р58��4��Y6;|�5 �ĵF�=��+,4��6�����R6�aе�<����;6�I5�j6��7���	6fJ�ؙ�lW60��������4��eR�6���g�>��.K�:L75!r:���g6@�{5�&ʹ�(���7d|�4h�5�~���ʊ6���3B����u���56U�5L����l|5�ya5:q�50���!4Nͩ��:?��u~6�/��"5K^(�(d���z6���5�K5���������V3��6N�/�G������4ȉ+����5����U�2������6ܼ3���8�=��g5l_�H.�!o��}6v�Y6'uӵ6�6�k�4���PBs6��ҲȻ6x��50���U�5�6|�d5��4h ��zWx5�W5���5�4c��f�����3r:���~06{�>5  ��	����������������G<��:L6���5Xé�@������a�5a鄶��T���5�`V�Ī��@��58�e4�&X6�l4�k�6�#�$�F5��n�赨#5�U������5��166,n6�S]�����5�=5�W��.�5>�c6�7�5�7���=����?��4����39m����0~�3����&6X5��t�Z6ݲ;� �A�p񨳀m�4{��5:�M6
�.5�赝p�5r���T��6J�96cu�5-��5���� �Ƶ��5�%�6��~��6�%�5�ȁ���)6h�$6�5!4�<���6ܬ��X��5p߲��O���5��4:��5�I�42E�5"�6F��5�z5 ;A3��R����4T�h�Ж3�ʉ���j5,�4\�5��V6ֹ5���5iE�6t�̴�V6�6y+4�������y����"���W��A�6�Wi�b�!��?���j6��5t��5�16�r��
�p���<'��m��ÿ}�Va6�#����4@�6y)����5N�n6�6�6[��5����?	d�6�4#�Զ�jA���}5k���^<ٶ81�6СK�l��bp�5%Sz4���\�-6D����(�5w���#��6�,���&6���5��V�"7��%6և'��uC�8�������I
z6�ϵ���?���B�5�\b�x#�5>L��<�5"+t6�6X�X�������6���6h�~6~D�ܓA�����{�S�/-����4���Z�5L-�5e���v��V��GS6�+�5<��5�06���5�����j@6A��49�5�[5˅W6��65V��5LÒ6S��5σ��J��]�� ��2x�5�s6bֈ6J��5�{�e��5�q6���6d�J�|�6O�G���>5!���k*�`b�6���6�4�d���PS�����5�8(3�Q����N_0���a�?۝5n�x5�W�3s/��6n�w�xڥ�S�R6�"Z��޵Y�E6<� 5�a�5�D�5@G9�B@96��6�Z6���5������=��"�5l����I6C� T,��6I6����N����g6^,y6x�(5q��T66�62��5DZB�0l�6�lֲ%��6WI��"��_���� �F�´*�R6��ȶ`505����d6��7�q�.4_WͶl��;�6)������j9�5�&���R�5hb�6R��5��y6`е3���ɤ�5$"�4<��4�ͽ6������5��5$3?6o�6S�Ե��40��5�g�6����إ	�t	���U���V6:i�5\��6b�5-5��o�d\;6- �5G�9��45�o��.AD��@�d�a���4���� ��Q�6��9� ��%���+4��̶=��6��64.�����6�'4��d5�6^K�5o��4��5M
k���9�W��6D�4���6���bmߵm9��Q6;жZ�6�46���@��5��5<:�>�$#!�}.6��� Ͷh5Z�6F��5�7�J
���5��26�8�t�Ӷ�Ͷ�6��/�6/�6�6N�������?C"7�l�5�ڏ�p��xJ�4)�#�\�x�� �5�x�3F(�6��68^5�m��񵠵B6�~6��>3�6ve�����>�/6�q�5Y%y�����Pw�(4�5��28��4��I6wX��j
��W�'��ð6�"6� ��|_�45n��5�2��-m7Q,6��l��uF�����y6$H���6���6t7Ͷ�2�Ǻ������05�{�56G`�l�5�ǝ���M��u5�g76�+3�)J�+����X�f���;���6V�����5�Fȴ]�e��N���r��Py�6��c��Z}6_4:��w6��J��w8��˶��5�4r6 �2�L�6К޴�y�6��/5�*/6�`-7��J��B��n&.6G���0��6��6��Y5����ц���D5(g|����R�5b�۵��6���L���x�� �r2IK�5춉6��`��#U6��4�\ݶ=f쵾�7�:����6XDz�㷔6�����q��}t��{6ؠI6�ǫ�%�6��
���8�I5�Q�e�5"&X�w.6h1ɶԍ46��7'�7�(�ز�6� �U#�6�)���5^�78{j5�1��x6�*6��S6�6)�~6�Ჵ2U,6�%.�.�>6.뙶���Iƴ��H\�����X�X�����t��2��-�(|�5ؙҶx�5���6�{�5c���d_�lU��w�64�N5� �62e�6�cc����5ȱ�6h��e
�5���5� � �y��������6X�4��6� q]��@�6���6&�6(���4�5��̵�]�6��6f�%�Ol��a� 6�r���0+6T&�5lQ^���[6()95�4��J�4�J�����*�-�eu�0̖�P����4H*6hX�� �y���X6�Z���$4� E�#������@�5�;�΃6����&��pᵨ6�5���4X9�^�'6�����[���46��4��!6~�׵��C��
��� 6��q6�H%��5}�?6��A6X>&5}�(�������5����4�s5�8J�p�۳��@�4{95��A6[�5� �6�-���$!6@��y|@��p�6���5Y`��	����SM6d�3Bğ6,� �pb5	��6���4�c�P�5<�~5�65�`U��;��6�6�W�3��N*�6ZS6p��c,6�E��c�4|�b6� 0�zm���+� �K�\ж�g6+�M5h5�5a?6d�v6v����f5��'F6j!6�Ҍ6���5��]�R�>5�`~�4�Ɨ5��2<��4���5.:Q�c
�6x�_6'	��-� �6������;�5N����n4�P6��6 7߲u�61cU��,�62-p6|7�5�5K6W4�5�ZF6p"�5;�6!�51�;� 8!��5�5�06 ݭ4���6�*Q5֬5>6~��5<�ǵ��g60��5d`��0�p5��U��p�5F_�����5�#�4�.I��L�"u�6��5�}~���8^-6��6�p���3&���69�[6�� 6�|�5�;�5�ô�t3�������^�3��� 6N�6z�6Y�ٶI^5xk�����5X�l� 	���R�6���5\ ����6Ø��ܵ���5��<�`DK5��6���ƅ6|��Á6t�뵮J����Jg5Z�6MO�6�l�5�~�����5+j��2�׵d����5̔�5���Z��6\��v?�6�<����A6��/5�]~6.	���b�4Ri���ZE6���5"��Ɖ6�%5FUm6D���v6o���D6���:���:�x���-���6�2��$�5xm5��i5��n��1�5�S���K� �Ǳ�=��4]��M��� ��L��*صx�4$!!6H�5 67����̵��6���5���5)}�����?�5 �e�p`�5|>���%5���jp���5V��/6?�$���3�T��5�i���8���� �2l�����6ty�r	"���4֛-���R6m�_�VA5�<�6k"#�Z��5K?�5H�R5��k3!'��z�!�w�06��9���5���5 z<5޾ô&$��8�64���n����4�@�6����D��4��5����6�}��(�����`�B�!xO5r��4ZU7���5� ��������õ�C������(��6lZ��D���g:x6|xA6�d��~�� .K3���II:�Pv��q�B�ܲ�5��6��$�䵀A�5������3S_/��R6�I���K�鴵��6d�{6��68^��޵�x�H��6�?c6f��6+�5`Ӹ�����h5h����6�������.������4�.$6��5��r4����,�!�$�j5�% �9%���5������ֵ�1	��°5���5|Yv4|��5yX��$�t�3�ݐ6;�95�a�5��$6����hi� ����sg�8� ��!6c�|���<�'I��H )�[o�5�5�I�5zD6�+ε�U	6��4��[���}5���d��5�&5^��5��F�Z��7��E6�5���fMڵO�� �²���5P�ӵ����D�5���4�H5��6���dq׵��S�$j�4�C+���J6�d�6`��3}�6������6H�ĴR�Q�荵(X1��u�5[27�+�����6��;���6'��65L�5�>�Z)6t3t� �ѳ6»?�@P�iG�5R��R5�q�6�M6�b6�ɰ5��96?7-6<Rq���W��䜶Aϋ6��5��o���)6�R5�ހ�T\5 d4�/b6HJ~�X��(�/5�I�"l��@�4x�V4�mL5?�G6&�6M6X�$�L?q5Pil�4�5���5��5��㵈5V�y����)W6 ֙�q�16��58䶵�����#�=����5>�p��@1� /�}0�5ؾ޵�E� 8T2�.��i�4Je
�r~�5��S�5��5��ȵ��k���U������6X� ���4�u�(�5mj4��d5H�L��
��&�6H�U6�g���\��C��
��EY5P6T���2�5@���X���j�5�t0�}6u*u��[5�ާ6�� �i�Ӷ#�5�-������̻F6�U��8���,p66:;69s�C|6Q�5M�^���5 �4F�����ӵ�ɍ5����1���8�6U����p����ϵ�5�|K���ܹ���Q4�`A�NA6E ��Ncݵs�w5~�76�Y�5�AѵXM(��f3�m5���Cd�5삵	Nε\`��h�F5�����Xx5 伴Ҵ�k��X�D��
����Ȉ6� ��G�x�Ñ6�ب������4�P5�c���9?6��H���Y5�@4���4�Ǿ5�R���wb�!&b5ݣϵo ;5x4x��m�5��6��6��I��ǵ|t
���5��$����3����^�����4-6���5�R쵼��6" �
�5B����?���5�h!��64}r6����&#5j16�ϓ��N5몊5군�G�õV�"�|��5\^���<62wU5��j6�����<�5���5@z����<�� =��4�5��߳g��5" �5 

4����^���}�5B͵�%6
��d�5Ԑ9��J�5�õ씺�����H��4��G���o5ӵ<F��h��5|��:m�5�4����	�@$|5;S���|6�Mܴ�E6(�M4�/�4jH-6f�3�n� �*�Py��q然���fq�ֺ$��Q�46�^�6 ����8i����5P_4H�^�p���Sѵ�X5Hh86�(�5ؒm6��3�,���9���ߴ��|�X�>6��
5(�d5s�5y�	�H���m5����6��v6�Ԝ�Y҄6�\���6�ت�Ĉ;�1^G6��76�FX�� 	�0w=5��6F�W6М��C�ĕ6�6����@�q��=�6�{6n���N��6��^6;�s6�`2�О��۳6��O�&��6��F��������$6��n� �58b6JS���9(�C�����a6�F��֜�6<[�6�eJ�p�4��>5Ry6���� �t��5#����m5�G6�����t���S���@���om6��:5:��5
�5��?6��54���B����3.�=6����f��,���#6�@f6���!5(帵�A%6���5�$���1�Ģ�5^@��4ե�T6�4���5�Y6Ă4�rֵT7���g³�լ���5h6�伶ӭ������񊵺՛�Wk����tg"��6.[�u�<6 ̟���T�I��5Dv�=��5Q�U6��V��>��6ĸ��昵@Un4���6��5gt�� No��ㅵ�x���?6�O���v��H�S6F�Եϵk6����ز>�¿�6z��6
�����4��/6��~�6q6�w�h��X6b�x-Ĵ�l4b��~D���RV5~��@�6XW�6�]�wc`5�¶Y�*Bt6��H�`]�6��̶�,��z�7�e5���[�6`��4��Q��h�5k�I5�Cϵ�68�����U6}��5d�5F2��Y�6*3Z�hԃ���ص��Þ5xk6�3��Q�5 �@�U� ��fÀ5TsĴVR7�I�����l̄� ^Y4D����#5h���E��5 6�3���315��:6"k�5F���6E�R:��������}�6� �|_���6�e�]M�L�+6�s��%E��/�6�d6���S6���U�6AZ 6��70;�5�%5��~6�Ҷ�O�5ֆ6j�5�<:6X��4v�1��*ɴ:�����J6��H�p��3�'K���̵���50�[5�	�|��6R�[�@�/�H~:������L���ŵ ��5�q��Ç5
�6R���9�6"�
�pj��H$�4(�5�� 6H�C5]�-6��+6��d���46!U���1���\5eM��P�6�6�bO�^�(��6pA7��̵�6r6	���w�5���K�4��"�❑� d����6�?$5�f�V&-6XB6�K��пA4hN 7�'1��6^����D5��6�
4�#贈vr���6�U6�εxA���;��5H�O6\}������v?6��5��]5��'6,�}6~k���C��B ����61*�x�D�h�!���Ѷz�6�a��g�'6m���VM̵�.~��}6Q���n.�@����y�5$I]��-�*�6\˴�"7�(�i5�����T����ڼ��[��6Pr����2!d ��Y6��6�;��]6�}�dR�5hh�5�u�5��|5xƵ tz�z�4����n4�6:P�6�&6D�5ܓ��LH66�w�5�R*���k��6`!�3{'C��;m�hLn6���5V����<��Qn6��T����5�%36���4���Yd6�U���}��R�m6�Oz6�Ao4H(6��'6�iG�P?�i�v�f��5���6��6�F�3`�ö5�6HyL5Cõ�U���^��yA�l�y�N6�F�5p86@R��{68Q�dQz6�V+�5TQ��\B5�3��o���r�tIc�@}|3�f��#66�����6����
��6�]�������E6,��T�E5��H���G6$j\5�����X�5�r,681 6��s5 炴(�ȵ�w69��5���6�f���?	3h�6O�׶c��R8���O��Pd4�ܽ���`6�ɶ�X6���4@O�H6�5�����k�*W75�E��Hô50�W��8f4?!B6F�6 �2�⾶0�Y6����F��^�����8⯵���4�'�����#(�
�4E��6�4h�5�z6�*��=��q����̵X��4�5��6��6�E�5h�ѶZ�D��[������4�#("�r�66;�J���g��(O��[�5��6�*�:J��۸�6��n���F�p�P�����4xݶ�l��L���	�5p���������4Ͼm6hf7�3M6���w�#�`{�6��<�������^c�=A:����6�(۶����1�bYJ51�5&5�6��.�$��U�����6���2����r�H�ZZ6� �5 @�/�tI6i�"�̜T�<��5Ou�6ˈ�6MG��5��5`�ʶ�銵�0"5v��5L�t��W�6��6=,61^���x5iY�5���53�"7�A��ۏ��J�5�g���C�2/g���7�\j�5*e6V�s���J6�����5���6�ko��#5]��64ڙ6�y6���6.!���E�6��I�61�6���5^�5Dt����d�"���FI�6�X6y��6�
7�営 L#4���6FW7�7L���6�̊5��6痶H��~g6��7��m�X�����N�4x���NC���6�o���еE+'���i����6�=��l��gԌ6��b���6D��6W�9���	7<3�� C6t.�52Dc�`�A5Wu#�Z?��p�x�ն���:�F6�H�e�7O �5B3ȶ�'��_��5_�� U6Z��5щ6���-xp�q =5cB�6�pH�ٜ浚za6Y�6�E���(�Je6������@6�,������C���X�y���6�B�06�3a���.R���6 Y�����^'�6�a@��|�6V_6�=��6.�R6>ʼ�M�q�@��vE�4�7�¸�;P��o����6�Eų�z6TGK�;�4g蹶�&�6����c6�<|���f5;�T6�l�6�W6z�a5$��4��6��r�M�u�;�T,S�����66z�d��4���: 7�G����]:6!W6�R|6����}���5_qH3l�>6�u5 �G��D�6�C�5 �5&�54�	�ҿ6�5�HG5�t4b]P�I-n5Cv����4PS�FTߵ@�3��˵��5m����f�����4T�3�[d�Zz5�]<5��4`��2r�^���i���%��7��C���$����5@�(5Z�@6�9�4�r�4Nm�o�5x����!�hm���|5p&4ޭ�5X�Z�M�3�6.9P�2�Ե"5ce6��۵t������"�h�Y�MG���;6�-���q6̩h�x�0��H��R���y~���C� �^���6�zB�'�5��l6(��rx6}t��g���Q����P�5^C6�tz����4���4̐¶B��F�J�'"��4�6q�$����5@�ô�?c5�lS5�MƵ`-�5��	6��̴���в�5`�W�>u�5��u5ζ �ٰ<�:0���Y6#G��G�4�S�5Vg58O���k5����ς���[5�̮��l�5�����wk6�68�&6y#�5�9���t5|��58f�6��u��񊶠�$4'Y�����ɍ�-R�6�^�X�͵��
�t�-�녵AN���"��?�+{6И����˵Ơk� $5ꏐ�����	��6Q��5V��51�5�w 5��6�J)5�W��/`	�r�6�[�4�jV�@,ʹ΀��ﵴ�nM���5K?����A44�����5Y��h����3���fH5(Ӡ��T)��9���`�06���4w�U��4ĵ�tϴ�b5�1�6=`26�x)��� ��)6� յd��4��6+u������g������	�Z65�5�3�5�QG��'%�n�E�R�������=�Fy�5�_�>6�WݵL!6�K���6�6T�=5����~��x!�4М��J6�z'�RZ���D�@�8��:-�Ѹ9�a�:�6�4o5�[�lc<6�!��-�L5.��4�P.�,8G6@����&�z+�&;6|�J��B�4�?�����S��5����ø5��{6hxR6��,4��-� 2�2�4��5z$絃v�6˦6 `���!��?�6��5mKo�T�P��¶��;6}�0��54�6`�Z���u5-�6�������6�z�_\��D�6����b��
����6��t6���^��6���GC7<M7�fx�J)6�_l��^F6��!�t���r��4��Å,�6	7ꃩ�D��^�5T�@��>�
�7����oa�6�%�����6�~��\$���6�ص6vB6hc6���6i���e�����<:��,>7F�86�¶�{\��:7��?6D�6\ʒ6rQ̶8Z17.�/6�-��Ƕ̯i6�b)�b�`7`��[[��|�d�9
a����H@m�`��4�<2��#����,_��6��6+"�5vc�6P�����G4�i6�Q�X¼�ty7c�h�6O�6~��h�
7C	7H�n7���5QV����6[ 7���%7��j6��%6 ���$�6��ǶpE7 ��6;��J�_6`k������,e�6�	6��F6�#ප���$Iq6If�M<��U�5�s�����~6�ݝ�~�P�*��������̵��
�j]*7�#�p�ϳ�gص�6��n��5)D���G6���6 X�1�H�5��50� �P0���{6���60�4pd5�\��e@[6F[��6�\� �~�T�Ŷܩ75�8/��N���;Q�6Z����#���[7�O����Tm����5\�t5��G68Z5���5o	�5tj���r�6ڂ�50;j��'U���6���6����$�7ѵ�6�6o��6hOd���n����.���Ly��Y�Ѷ��=��,�9�;�n���+��j3�մ!��-@��9�5���4�a6H-7e+Ƕ�b��	!��5�V�aHt6:� 7J������6�X6�_��6�m"�K�G��Jյ�(O5X<]6^&=��J�6^l��@�4�ᠵxd�5�˦4���l�6�%�����6߳��K7��� ����%	7�W�yߪ�Z�6��@��#����˶q�n��2��cb�6�<�2�N��	7#���T�l�5RK5 �6�������@ٵ,�(c�5`�Ĵ�T�5|��[Ͷnr���ʹ�q�#�5SP�WS7�xP�Ɗ��Oֶ��C6��R6���t-�6M?����5��_6�-�4Qy6��5��x��,3���s6�5`=�3@N~5j��p�����5޻?6�?�6H�'6l  �ۉ�9��5�>6�/+6�`6�36�,�؁o����6�@�7��޶M��6��5� $��Ln�5A���	����6��%7�X*��U�8H��_�6c�
�b�X7j0���L��끖69e9��/�6&J�L�5�S�6R����T85끎5�d5v<
6��¶��5�:.6���|X>��y��O�aπ6�ȼ��9���6{���ȴ��c5(�(��06,�5�����F�5ߴ���N��\���u6��6��>�v^R6$�t5���)6uӵ�.�𷁴!ؚ�����Xߵ�z�56��L�׵���4���6��Z6V/\6�Z�6�G�6eq�6[���Q�5���R6�ץ���6|u�6��A���t�:�8��y��a�6�Q�h��4���.���>�6%�ֶ$�5p2õ?��n͹6޽���%2�6�hֵ���6:-���dd�d�k�`\q48�Q6�Q#�fQ7+m*60�O�tD�D �6��J����6S�������#��r���.6zO&6g�=7����F�V6=�5>v+��546m&�69\ȶ�m�6�f��{����6�V��L�'�un`�*��6�W����s��5C�6L�P�����O��6�To���o6zC���(6 �6$~ζ�B5x*��g����w��\X6�
,���6�˥6�Y�P�6|h�ަz6�1�6���5*�6����pwY�~�7��V�}6�5n��5�N��>7A�,6��6Z_��|6�L�4Y3�d,7�߃�^�V6F�c6��aW��6�0G5M�6>!�Py:�ە����60�Z5��0�p5XH����6��A��15"v6�35������S5v6pJS5$��4^��5y#�6faҵP<2����4��60-�6G9�� �3���6>6<���nD��t�\/�5_@�6��~6�1q6ʙ�6��6�+�6�����6]�6���6�U7��A)�0�����6�Ax����6B����]b��N�5b�� ��6�1���H�55��k��6���4��{6@��{0���Z6u=����4 vص�<�6,`���3�3�l˴���yq��6"ά��6�6�X�}5�6��״�d6t��SS�3���6p�� ��5X�b��s����6o/5���5`�5[��,0(�M���
Q�5��
�H���U�4��<�&���<�5�z{6x`�4��t6�;d�_�j��֟5_�dC6��4d��ƶɑ6�6f���R�.%(��+�?��� a6��5��|6ql�6�lb�Ͷ۶_��������6����"{�f�.6PJ]�n!����4�ʘ6��	�^ ���t��*�
5D������4Bh�k��5�1���cӵ�k��nM��h}�?I6�����6:�� �3�M�4&�C6ǡ���"6(�d�D ������a�|���S5�)�6�<6l���q�4�gY6��UQ��ɶ?���x��5��%�7Aj6�(5tC��f5s�6��2y5&�)6�6���6�o+��ҵ�"��i6��5�����*76<�H6��L�@�K�Vdܵ]�6f��\� ���;�6����6  5@A5q�ȶD�Q5'���h6h:"����\��� �����y�6 �|5"�ٶ�?�6|e5fq8�O��6�\�M�C5�4�F�O^P�����떵�Ki6^�5&7��ܵ$�q�Pq�4F�]���J�86�vB��mҴVt[�.�7��)6��c6��6�X��
�\-�6�wж��6�]������s�z6��϶�[6�<�5�?�5��ȶ��6������y���Ɲ����5߈�5����H4��6X�6f<���R���Z6��
��?:���~����(w����?6��v�֩y�f�G5�`�_"?6�Yi62Ty6�[T5�!ŶZ�¶$�m�\Bs�@��^���Q���
��(�5��0�	7
6M`���5h��5K��6Y6�궨�S��6�`����=���&j6\�6��_6��5$����ƛ6>C�6�ô7�����W6B���  ��i�6y'/6�`�p�
�-� 7 �±�����A�5�O� �)6^*
7���L4��r�Ą�Lm����6�"��I���E96��Z6FR�5f�j����4�낶O(#7�攵���5�Y�6e@6�+�����:eҶ!u�6z��4��?7ML6��6$����L��첊6N�϶�>7\v�6���5�X�5:(����ҵ_�5�C�6�{�C`16Q�J6��!6�Qi��6��c��t�68��ȓȶ�h4��57m�d��4�����V���ŴPr�6n�����=�"�&�P�����L���5#Jܴrb6��^��`6H/����\6q��4��R5<6���5�_�6�����ֶV6?#4���X6��ᵚ#Q��=6x�6Nl��4�=7��v5��x�l�@5^�Զ߆6���50�Ƕ��εHKR� 6��6f<06�m:6��ζn�%6��6��`�D�"6<�,�N��6�%6�ɵ	���-ٵ[6�%�5��[5 ���8�=5V�f� ��3���5zv5�hZ5a�Zn��T�R�u6��5��H���4 �#��˸4�6$J�5�O��kx��&��:����g��l��=��53S�66֊46���6Oy&6�l�������z��x����d�&6���7,�5���6a/�9vX��Q5`_Q��W5�]�6��%6Xf�5��5ل6�5�ehu6 bT6r�g6<f���d�6ɡ�e��5��=��NO5z�5@j��3�q�������51�5�N� tA���5xy6F�%�nȌ5���5�H�4��*�k&6�Bĳ�>6�	�����m��Q�h��u��*J5�I�3@ֳ�2�(�ݧ$��< �^v5@�I3uW6��68Jo6	������6�X6G�6��i���6���5ܱ5n%�6ܵ��2���5�LS��6?����qs5GK�5v-ݵ�B�5?nX�L�6�d�4G��#6Y3�5Rw��x�6��m5�W��3�Z���m����5J:�v�:6���5�A�L�� ��5F�
��+
6.�[6Ĉ@�$K���gT5K=69*����3{�����<6-S5	�6�\'5��9�
y6��b5����h@̴)�O�5��a6p=��[5���V/T68�7���45��5'���4~��4�6E���a5jU58'v�T۵kȵֻ���+5�<6k-�����������F�`�6�_5dZ��H�ݳ䰎5gB��\�4k�65t��5�ϵ�7�A�4 g��1�_6Z�����5ZKB6vO6N����D����5U<)��&Z5��5��&���T����V�q�`�N�b;��y���I�J5�q6$L��WŴ�ɇ�>oU���<������M��
"��6j��4�
�5�66�´F6h�C�М�VM6E��4 �N2(p��R��5�q~���M�LZӵr�5�&6�%v5x;@�\~K5��5ύ�5��I�a]5TJ��2��h�_�%��(���b�4 ��5�gL5��R������v�ѵܦ�5SF5���5�R6`'�8�H��ܮ5z/U�W�5�3�4&y5̸浊��� ��4��t�㏴c'�5�����G���5��#��O�P#��H+6@�����4��8�s��W�5�u�5
F6�\ش�Ə5�Ћ��`���=�:�Me;6��65�I��!� $�3ѮB6�>�����5,Ë5�|s5�+�`������q�(���/��CJ6{=5 g6�&H�p��5�)&�e�6�� ��}Ƕ�A64���@6�H��.��6D5yp�6���5dJ55����?>�����M�PwӴ���5r���6��V���L� ǖ4l�16:#�6�I�52@�6� ��\�Ӷq~��������K��-16M���L�5��K���0656��7���/ܵ�)�H
�5�L[���7����x����50�����6@�Y���ضP�͵����c7c"ζYa����8�l&7��A��b6�ä�	6�ib6� 6Ս����*��5�{6�"76�(�6��#���57�9�5pSֶ��6�
n6h���g�]6�i�/�!��r
5	\����-��,�76P�6�E׶%|��u7eU6˜�5�zr�R*���_5�05^r]7���6��7���<��6�#ֵ�j�6�a�6�k6��6�#�6��n�f�6Vh66�S6�+��I���o6ʤ�5;�6�?���e�6�Qy��W!�`.ҳ.
�4��.6�X�5�U�6���Hv��xƙ�l���;'5�ݏ6 �(6���5
��66p'5^�6�
���1���l��R�5�b��Aöp�Ӵ}A7���p6�6�6n��dF��~�5���5��D7�16�󵡸e�T�0��ĆY6ȼ̶Kj�6�r^�F0j6PWb6���ĹZ6��=7�g�5X���q6�u�L��6�T6��%�<%5���5Ƹ�6��� 60�W�9���<G��c9�̓���7
	��L�\6�<��x�5ǩ��x�54��5��C�:� 6�r϶@�`7xfC�kW�6*���56��66���5f$I5�(�6 sF�HF96��6�(��%6�h4��д�w�6����3�5���6�X�6Ȇ�5�m�6<f�z)	�w��,�6��V4�!"�,��6�N*4\�V���f6ƈ;�b	C62L)�؛n5��*���m����6"~��A&�榍6S{�(i�41��6�\�+�l6>PZ���γ�2�5+�)+6G����5n��*�6r\� T�4���dE6��4�kM3/��,��5��?�_���㋴�;���o4͢A��Ė�̎��"��5��6e����06�TB����6�~�6���5Xt�5�@��T�I���6:B���\6��������67�Q65Ȕ�@S5��6�}�6��J����Ձ6� 7��䴺6�f�R7w��5�Q6�ڴ����S/6��7c��6Z�T6P�1��9�5�x3��7�6�36�T6FX�6 �'7Ȑf�����AE��h�5��6���5�8�.����6��6�
{4;�0`M5���2�5���6�(7�5��6Y%�6�#�T駵빍6�g�5�Q�6R%�5�3	�+0��62=6dY�5�E�58ˍ64}�5�G��n�׶�l�|�45x�ȴP3����6�&�3�5������R�n`�9��6�d6���a��4Q���5J��$����6���pI2�`�f�z6=Ժ64D�5�M鴰�ֵ�V��7��5��ζ-�X�(�4��5w�5�.7d�b�!�񶹫V6x�<6��6(\r6���4��6���0�T4�n66�-!5a�$��[[6@>�3.�~6r��6�9�� yA6��(6tz5�5�؁5���l��at��Y�5��6�Y66��5 P��{7��մ�������jյUԵ,��6R������4�7���6x���uٵ�87 �5ǇP�,zǶ�C����646�Q���{6��J� ��2��7\�e��C�x׆��?e5�&�6[k������Q�6^��4@����f�5
��5�F��vH��o6@؅��9�6�\v6��ɵKz�6��L�\�j�N����ص��I�!���5V^m�7G��w���7�C�7N������5�"��ʋ��J�6��0�`x�3x�.�|��5�? �0{d�_޸6�b2�@c�3e�� �5��X�3$'��8W5P�3�3�&����
5Fzv���Ŷ0Q!�=���>��6US��m1�6�՜��^��XK�p�R���P6T�6��64�5���r~�6莂��?y�� �5��2�((�.�5\�60����3�6�t�� l6fF��@�5`�H4�;:����㱛����c���
� ��2�w�6@ؼ�=�,���ܵ�&7�j�4�C�[�6�#�5�e�X{|�p�]51D6�ъ6��F6\�:50��3������'�#76D)�6o넶(��6o�x�U6]7�6I��
�5��t�|0�6������"��8��5lX6�S�6�������6���p6�5�65��(�j�}��#6�XO6VӴ6R���=%���+�P��4�@����5$�o6\6 ���� �vV�5�ƶ@@y4��⵬y6��5z��l�l6�Tȵ\g��fA���7U@�5x(66X)6��W��6��5�_϶�4�6�y�6�W���A5��6ւ�Hq�4�L5�̶̕3��<\6e���2�R6�jh�����*@��(5�vD�$��6�5�I5ʾ��]�|��Hд�
��к-3j��pq�5 �W4�{6�fN6fҢ�5ˊ�����B�6���5����࿵CW��������봸Ѱ6��5L�Ե�U��ę6d�5�3��e�8;�6���� ���ׅ��{r3��G�<&{6G|o6P̑4tz�6d�Ƕ�Y6��6�� �f�7�c��l6���6F�����F^1��`����*6�됶��5?!�6U�a6�>��n�#�C�c6`�#�7�M5�jg���6�o5�Ӎ6�6}.l��1�������6��_5���6�)����q��8n��b�6n����y�5\૶����5�Օ6b4O6��x6�Fh�N��5p��� � 6|���7^��^�6D_�'´6�ص0<6v��6u�5oR��4�5�I�5\q�5�Ph���6�Z�5Kђ�D�#5�c�6njL5�Y�.ޛ6 ��5���5���428���95$B1��96��(6d�5 L��@��T8m6�MD�D�G5��F�� ���ͣ����̺�6��� W����5�u6�{������6XJ_6�`,�H��4*3367?�5���5�p9�[F��a�6�p�6�8���#��Pp8�¡%6
�����5Dc}5�.�Љ3pH����4p��pyԵ��6Eq.6 T	5��A��U�����62��6�^��H��`$i3�2����6(R�:{�6��D���X�d;6g�6��h�|6P'l��q��vǵjW�5r6X=7���5K��Y�ʹj�6O�5�26襑5Г&���c6����v�5t.-��6���=@+�'��`[N4v	7�:�5 ,��t�6짶@����6��w�������(�25�A��*���0p��5�����6е�j5�.�Һ��N�6H8�6�w��66�16$����5��5B���!״�Y/��;˵uKK6b�C_96�	x���ǳ�۔�L/۵��,�u�$�6�-�5M��P������63�6n���*.4��p"B�m�'�K��6�������#6�E5Չ��Lb����5���6�N����5�$�5�6�)��6ܶIF�����ܵ���58�5�,��x.a�����@嵀">5` ��86=}55�%6~�K6�[@�/�6���5���6rݍ��.6�]������k�6�$]��9\4�6��s�>��O�6�5�6��t��\�6��m6��/6g��6 a���_�6\�P5qj�f�ʵ�6��6�x6z㼵��7pǌ5�}�4h�ٴX�5������6:52߱�>_�6&q7�
6��7}��6�>6�M7Q6�n���ٶ�Ǭ6�	�� `4/�1�1P6�	78J����5y>���c�5�Ij6��J��YE6��5�t���S�/6�h�5m��ȷx6��Ƕ��e6x��6`ɶ������7��R�e.�6��U�\66��oo6�*��i��ҽ�2��5�6P5�����F��"6�Ox�ԠI5��T�ا�4� ,�l������6���6�§��Z\�J��ε⤤5'<�6l�5��6�QԵ$Y��C�6�8ĵ�����P�l�x��p���:��M��/G676Xݕ��a�4��3�z�41�6��}6�=5 �*�<���5�n�5��'5r����y6t�96Y�������6�o�6\еу��\Y��
�474ĩ5p�6*��5�u
5���D�,�Y��L��4���5��ʵ�x��-���d6 �6�Yʵ|�{5k�"���ٵ�� �h!���$�60��c<�5|#����յ��q6u�s�7S���D5�*9��+���;ߵn�ŵ�-�6F>6��5�C6�q�5��۵�/�5X4i��h�\6v�4��@�>}���z6մ���� ���5Y}C����6{�5�ɓ����F$�6�>ݵ�0����y��p�x����B=�h6���5�擶��D��i����4Jߙ4g^��,ߵ�/��p�Z5 867 �3�!5����6`6kY5�L6��6 !��P��6���
r��c6H��6F�t6�S� t6��5��ŵ-��6����T��|8�4�"�5�?�n�$��4ڵjy,6f���#6t�5���3|]I��5���LW�n����zܵ%�N6 ܕ6M�]6h���@,7&�$�"����(�:�ҵ�cD6��4���(5S����`K%6MH6�A6G����Ե6*6��$��N�fhZ6 �z4��НL�C+�5��M��k�4�#���rʵ����U�������b|�����艀5�Q���e��j�6�¶��5l@	�n�ֵX�]�H��>�N� �94�ǘ5�I�5=]��V6^.��:����aj5�t�Tz&���E��5X?G60�#6<)6��[��D*��z�5�e�
�Q6��Z��4�6AFµa�B6�5xt�5 暴��6@�M3�\~��]�\C6<F�4\~S5�I��6(o�5 �W5 &41�#�++M6v���㧶4��b}ֵ������5�A5A:%��W����5��l5�36�(��c+� R6�;��`�\�_V����:��d=a�ǻi��o.5p�5��e�&ᆵ��T6�>�b4JH05�1��C&I��044?P�4P]������N�/�f6Ҁ6�?44:�5�P6�k66�삶,_Y6xJ6T^_6Q��m����i6�'6*���xx����4o�����޶N��p+#5bXV6�:�5_�=6�.�xq����[�`���w���R4`rԵ���� �S3���_a6��9�T��D�6�w��d��5�6�s%�n���ޟ��`K���6�]��x7�6���6�����~Ƕt�5�A��k7�k6�"!�l�۵�	)6�O��I���6&T��p�r���=�*�N5P�h��Pu6f�HlC62�3E���6�4���4A�5{�e]_�#C5��5D��5P*	�ҳ
��>&6vDm5(�W6��� �M�bͷ� ��ě$6� ε��5��9�6ƒ�5>+6@ַ�#{/6�)���S���46d��5连5�)�����5}5�B�5�2õ�5�6o$��,���Me!������50�4�Y%P�� �GP6��϶l�h5�`���5�5���8
���NR5��y� ��0��xt�5���㷅�DD��i��`��3�l岾B6ꌛ�։6���fLI���@4���w�D���3 �x��gε�����jI��`6d�-��3xz���]��d��4��R6�/5h��4�7�<E�drq��ZX�����Do�(\��<��5�O���~@��}5Ҳ<�z�ڵ_�6>����5k}��u��aB�58 "5aM���85�KF����	���ش�6��|6���5W�U64C�7R�8�6wFz�$6#�XҴg�+5o ���6��64~�5V�6��N�et���`X4�V߶H��;��6@~��Ȑ�}�H>�5$�H6�s �`�M7Zö����A,\��%ɶ=�)��	�?$�� <N4��56��5r�ڶ�Z��0�5	��6sa�6��嶫��6�҄�9�x6���6ܘ�4��[���P��� �D�PА������#6��w6X7��y��6=+���(7��54\��ֶ��ܛ�5J��6|��~ �6��M�c◶n�4X��6
�7*纵�+6����m���󵬵�6P�
5�7�6� 7��}6���!O�)�6��P5��6bT�5���� �c�R��t�33@�� q���b���6�67p�L��P05�������6����+`6�ʂ���\6@L�4�}6UJ�6 Ke�۴�4h�N��>�6�Q��)`��1����\6N���sdǶ*[�6b�6Eo�6d��5d���\�`;N3�9�6J`5�x�6�>�58�5��6��N6 �X6HGT6����h��*ʶ8N��|�5o��5�\}6���4�憶E�K���6'�6��5$H��s�5�Y���D7ό����$�t6�}6,W�5�1�6efW���F6`̴P�O�O%�����δ�����5V4�6 &�6 �,�b�5xn�6ƹ̶���6'���� �5������58���j3�Q6<t5ې�=Q\7<����6���5h���k�6֪���	ζ�y�

<6��d�P*m��t�  '����-�6���53������ ۷5�.������{�$I�6 z6�\ 6��h�*�;6��H��!7�E6ꕽ�"��4b�Ҷ���5J~൘��64��@�+�@�77!��6�,6�x_6Q�$7c�H�1��6�q(����|@�5��}5�96���5�ff6���5����6g��.4�9���?7̠���~�6^�*�G6O6�6h�f��+E�ˏ�^S����u�֕�5����e�B72o�L�u�(�u5`�4u�7(?��Zh�Һ5d�4�X64��5��-5[��ڥ1��8�5q򢶊��8H}�ຟ5oي�	�!6CV���l-�'��"::�>7���!ҵ��4��f6E!����5�3Ե�����a5bz��Ml�4��W���T��m�6c �5��q�.���5D^��Qn��Z<&��l�6��7�� J��N.�)=�% �4��ѵ�Sn6�����53e�5���T3�6��6�x��M6�ǵ�#6����$��&k5 #�5Z���h�5��_5�ٯ5L�!6�5��
D�5ک6�U�4=�5��ʶ�6���T��6h5>�.u6ҧ�4���5�~<2N��5��6��26�%��HK�5�^��]�{酶�6n�6�p嵄iٵ�F5s��D�q6��6O���ð�6�M�5��3��Q�BA�6�E�X�s�b�D5->�5
�K
 ���6ՠ�4T�57炶���6���5�m����̶��6�x�Y,4��F�6����O6�E�q�X(��=Z�������⵨j�_��6�416L������ѵ'v�6V5�Ԝ5��ok�4����������5�1g���6����-�5*��l�4pݵ��4QLt� ~/3��x6z$76�dɵ��˵������6U6F��2��Z�5�]E���6�_�����5��6���`�6�6��t6�Mϵ�c7�,���e6��`6�8'�3J]�-[
7jR�5zph��0�6�'�5�Bd�L��6��i6¢6�J6��ĳ������5���6'�k;J���5T-6�J�6}F�5Pm�6Z�����Y6��G6�g�����4���$�h5B $5��Z�� 6���6L�m6���5�W6���췸6���6D^,6���5k��V��6�Sk6(Z������,$��7���!�6CV��4	!5A�5	����ڄ6/��6��N�&�赨=[4J=��k`�5�v�5����&�%7���5�K$6�.�[I(�^�G5�<T6@#�3�\��ve��G6 �6�Ǳ6�6���]-6�2�4w45G^6=�U����6 ]�dBJ6�ǳ`U�(�5�Ū4ַ5v�R��#�5�>�R��9�&�pn�6��g��,�5�g�5�Y��M3^��5N�F��4���4�̇�����!6֜M��5���4�F�CU��x�H6��6��4�և�4q�TO�4�&�6b�6\M�4/�5�e�Pi�)�6�����p�4<@,6�	k��	�ĂL5�B�$�?6Xo06ݕ 6&7������P6T6��8Ǘ4��3��C�IQ��lƴ5�52��5�l5٠�4/�c��]��G9�6|@�5Dᠵ|8�d��4�-x5f3�5b4
2��5�Pl����5 �Y6�Ӹ��c�5�V>6�z޵��5��4�P�5�X𵄞����5����G]�6_��5�7�쵾5��?4�,�6�n�6û���Ғ5�2"4�&P5�o6^³��8����5�5�� <y������u5F< ��06�j$6$D�}KI6zW� "��9�z6�����,�Xd���D=6�y�6��5��M6�6��6��z6��
3��56�(>�M�����5Dٵ�R�)�&�� ;�5�D��Թ=6�G����2�o��6oP�5�F�5��-506���}I69f5�|5��9���T�����6���5P�t�H��5[�5a��6�%�4�e�5n���"S�6&�r�����h5�����������57��6�"�6ZF��T6�m��(U6��6��	��k6d�%5��5`pm4�
6@��4�5��(�;�61XP6��4�;��3@���6�P	��]��6�y�61S��Pm"����5�786.6>5�t6��|��6�=K�V���;�5ȱ�4��y5���5���jB��0����|����
H���V4_���@�ٴ����q+��ftN�Ӹv5k$55P;]5x-�5:)�s�굁�������5a�5��d�۵ж%����1!6d8+������U6Z�6*��6�=05V61y7T�5)P�6X���|6p��4Ѹ�6jq6s�����6 �/��[5
����7,��5�u��Ln�5ȣ���<�en���6��6�Ķ� ���V�6�2�{8ܵ��5�&>6�t�4;��6� T4II��DA6��x���Z�*�a��5�F����7d�g�6�6WK��@��226b6�.��nŇ��NW6����\� �6��6��f6ܽ��F�(��ć5D|�"��6R�h�� ����5��}���d���Զ���5@�h�@�'�c����5T�Q�g6�'86�}3#��5����S06���6`CG�,���v��6:S0�ؠ�?&�P�y5lS��6�Qm�ϣ�r����V��͎6�ǵX^۳�A�6f&���Ⱦ��-˵'[���76��46�pŵ��9�;�ζ��6� �D����͘�P�����4v�ԵFs6�u���a�6��5����r������$�C��Tt6��46h�50V6��%�ge����6�L����^6�Ỷ�[j5�@6���6�9�6�ߵ�vE6�WS��Ȫ�23C��"�������6x��5��u����5������6�%�5�6e��6��0���6ܙ�ª���Å6���;����ի���s�6������ĵ �5�մ	 z�&��6uo��6��o5}��P-)�N�C6�ൕ�5|��5&�I�*X������f�@�6��7��ݶƸ6���5E�N����6����ҶE"�6>;ٶط��yv�\H�5��5(J������� 6pw�5 ��2È˶�3r5�p���(6|g6(o\4��жB0k� 0��G��{=����5�9��^�{���4�(k�*p�5b���q��6������61*4�� 6�6V̶��4���D62|��(_5��Ͷy��6j�6l�(6z)�6�ɕ����2t6Xv�s|6d���7��n��6�eS�,dq5 ��23�P�$4� 06�%������Wv!��(K6�U��A�4��5�-�5p�9��7X4�r���3NE6i��(�1�{�4X]!6�~�:W���6�5r�4o6��'���5ي͵�_z4��6H&5x,�5����Hwõ�y�nE�5�[r����-5�	�96悊������8���{6�6>�4�0�5X��5��ǵ𶱵 �B�������5~K6v��3R?E5��z6D��5���4�c$6l�����j6�E���ڵܪ�6�7Q4ඊ56˵7i�59��5U�3� i��"�P�x��d\�5�e�͎�6`����6/5��5�����59c5ßR6��I6���5�����A��,#�5T�]4*%�4%{�5�NX6�*�����5��\5�ߖ����Vx�4�*56�|�d�5]�W���!����4H��5� �3[~���\�5<�N6�5��%B��)@5"�&�b!$���C6�`��
a�5���5��5Z�Z5�������v}46`���U4%<�:G���5��h_(�]�5���� 6����-���dе��P�8Ѧ4XYx6V'�5�!5�����4σ.5�д��V�\3���N)5KU}��5�
x�baֵ�Y��l��s��5�_���洗 ?6u�"6�*۵4��5&+���E�5�o�5"���|%L5;����n5�e0����JS6�e6*�>5������d��4��Y�&�k6�i�4�Kz5;t��Q��Ȫ��i6d׵�c�6�1��^�׵16l^�5Jm_6X�ʳh�-6�o34ˮ�5Z����1�4_��5�8�5㪒5b��(~���������´�$յ�_��J�Q5�-��x�̵�V�4t�_���"}�4�l62a}646K6��[+��.i�5R��������ɵb\��_�5�_��FѴEg���ĺ������3��3(`�XȪ��)��fb�5^�5�8���H4�������4<��@��֜3J�O�	��v��5���F����C�j�C��~�H�`���i��6ֶ�U�6�@�&��50TF6Z��6��5���4\>T5(��45жd�K5F���:�6zzZ6
��m%�6���6D�]�H��5�wu5���3�Bq���9������'7pP5����L��f��'��DM�60�7�m��� 5`�3 麶��g����6��~5S�T7�
�6{O�5z?��ڰ5X,Q6�2,���7��S�%Ӗ6���5����z�6��6Pd����6G��et�����6<���z706����T��!���6���5�õ�S޶���6�2��U�6p�5u��@B�4�I�40��5���6��5����^/�6�������3Y�6Jŝ4x��4vi��պ���6"QM6v����ҵ� γ�XL�Ut~���D6�KE�(�����ᳳ4�6w��6Y
������GF�pz6?�:6C@����(6Ҟ�6񚎶(6���5�R����`�&��6�o6S;����s6��{�	B6�ɶf�뵕��6¤�q_�6�rR7FZĵ�G5�7ֶHm��e6�����5��}7�a�6y�b6�k��d7�6]��5\�k��\���6�lB�����"5p,:����5�;��0�e���t�E�;�w�S��Ҵg܄7rG��T�6ݯ��9/�6�!,��޺��7�5v��5�8�6f㉶��Z���;4�%6�ʵX�5F�h�\��5�̶�A7t>~5缏�
$5�"6�n	����68���t��6�27�O_Ŷp���6x�6�7=�������]5Cv07|kz��v^��6��P<�6>�Զ �ʹ$�b�TП�x�6��q��>����Y6����b���7@�.����x_5���5��6L�5�`
��b��;+�6Ԧ���s�6�1;6�Ԣ6�2��r���5\6mJ����r����5T넶���54+�?L�6h+����#6D:�6J�����5 �E6��`�����TK� +I��U����l��³��
��e5�B6ک5�5���6\�5N��6�{5���5h+R5W|R� ��� 194����Dȵ��6�p}��l6�P����5�5���5�$k6ȳ��)ͤ�Nex��7�68��4����? �i�4��?3���4q��6�oC6u�R6�L"6�֣6ض��26tT'��ot�:�0�����}��8h'������5���x̴��4l5845�`4�����K5�t6r�5�ٴH�Ӵ�?���c7�6¾�5~�� [ϵ@�׵�	d�p_Ƶ�5�	��R��*�5n�8���6p�~ܝ6�[����6��}��7�4hv�5�6��4nQ˵�A���`���6��j�%�4���I5(��4�[50��2ڶ��|4x�:��ͥ�J�5�SX� ��6���lp6\��4���?Ҡ�(�.�48�6�u4������5!)d6�򑶤�w��]�4����&#��R(�5�v 60gn5r��5Ż���v!6@�\6?]#5O�/7�W��M�����5���_6���5�*�5o�J6��6r-5L�.5��ֵ�Z�5D�����`?ڲ�`��[5��h_W�� �x)�4��4 {U3^�D�yY���j5�\�6(�ٵ �)4fR�����+�[6\���|�5��5�����鵱?�5H����k���g��е0`�4l�75Lj��N�5�%5�c�6�!��85e�����6ݷ���6f*�6Ԭ6��+��s�6|9c�T��y+�5�����Ӧ��b7	�B�Ӹ�5X��~ܩ���5*������T�6{�.6D�Y�`�ӳJG�5���Y6~O5����t��6��.5�1�4�iյ��4.)v6�"�\Je6v�u��2г�~6�[�6xu5�-޵ J����/5�r,�(L6��;6e2�S�@6N��2�6�a7�-�����5s^L����6���5�C)5"u�5s��������5��5:�F6��v�@�33���6����I�Z؜���P�+��W���7<�+5�97�-7Pݵ	�6&�5�jF5��6��Y�6ț96�T=�л�����5U7���d35z�m6�.�6L���G��6[M���AZ6䊸�̫ �_���9�h6j�6e����6�e�6 ��5��6�67�҄��S6+�6� *�o�^6����9��\�6�5%� x5��@�O���_������5���� ޴U���5j��5�I�5����J�Y��7 "ö�~ŵh�e׶X3<����5�jж�B�����(5�;��V�5�"M����[G6j�3L�5Ȑֳ	����]�5?B�6�>56�K����	�#��6H��5�
5jl�0Ӯ6 e5`e�i϶��16�v��z�D?t5��96ZL�5���Y#�6XH���4�wp5s-�6"�ͶF볶h?
�KL��5�9��v���
o68�s�s����e6�|�6K�5Ĝg5��a�������6��Y��7PE����6�0�6���*r|51��p��4=��6 ���4v�5"��6PW嵊�浏#ᶊ�(��`5��� 0��P]�5fQ�D��h��4H 6�FH4�q�6�7u�x�(�oǴ��&6P��D�Y���д�V9��趱#7���5>M��x�3��r6�����3^b��f.k�F�-����<�v�޵�k�5D#+�8��6'	�8c�5��7h�4�#h�5
����Er6G���q�6|�.6Z��u'�6|K6������5C���2׭��6��E#3��լ6&~�6��7��������ZX6ՠ5>�K5����`76`�O�߇j���36��X�v�ɶl�6>��������5�r��󦂶D�I5bcY�&�����5�Q��؅�𹫵(�6�_6N$��Q���Q�5�o���U�4�c15P=���x�@�b��6��H6���5�wP6:��`���6�ö䰳5��,�xڵ��a6��a�IM�6h�ص�Q��|ƶ �Y��
�6�˶ح�6��:�涖_A��l��iZ�6�;'7Ԭ��q�+74;���3���6�c6f���123@��}��6*K@�f�6 ����ȃ�� #ócR�8�3��5�6�&06��G�����吶8�5+�'�Zd6���4��&�6��5y���J�6\a�5��4�X4#�K�bö��6ء2�����r6�6����$>U�Rp�6��Bܩ�μ�6>��6�
���/6+�6�z��>�6G��6&󐶑ˤ� �+����(\}�R�6�
~�-܆�՚�5�t�5�q6�D6�Ӑ��޶�2�6W��6���3>X6RB6AAе3��5D��
�T5� �4�M���5`��4"�<�$��Ք�6�3�6�-6^��6�L����#7�We6`�G5�6���3F����m������N8�5N�6� 36�� 7�h6r�u��������n�6P�Ҷ��p��/7x{����5��?�A̶X��6����Y��!��>�4�����"�6� ���8�5�4C�3�ҵ�Z���YH�������`[�6v:>62E���X�6g���X����5�����M��Iට���ܧ]�px��r1�6 ��6MǵP= ��嵝^�6�X�5X��6V�6�\6*�26<�\�E�6�C6O� ��ύ6 �����6>I56l6z��֝7�ZW��P:6d�7����,����-7�k�����5`��4��d�?��6vü��v���J� �33��7`�(6K�7��E71�7��^��@͵^5�C�6�ザON���>6�՜���ն����M��5V�6���6q���{�
���#���ܶN� 7ĺ�4���Œl7r�7n�d����6�D<� �ܱ��G6Ȋֶ�h���R�x��69M��ZU�0��� ��!�Ӷ咔�Ƶ��H5/�Ϧ�M��6U4�6�Co�̐�6�����6Ȓ������.���m6	���b-��6�96 '6�������5֝�6���3.���@A�4��5�w�5���5@	>�۶�۬6LX��K�����ZH�6<��6��6܎j�tR85<�5������5 6s�����@���6Xa��G��t���� 6-h��,6����]��@\5LC�I6��,�<5�Ɖ��e��� 76zG��ҵ:m��(O�5�O�6c9u�jI���f@6��W� ��2��6��6*X�5Fe�B�6����Ј5z�δ���s,�p�3��5HF�6����+5X�?��<�5��v�G��5d�5���5�_���p�5ӝ�5�r���e��5�5��3�.6��&��}���|��6�e6���4��3��5�߽5�M�����bT{�j�c6Lbz�)�(���f6>}B���4L6i�����d�5;�1��EW�.]��0���R�5�7=���]C���c]6h�b���0��5�q����C�6�����Q�4c�?�@�ӳ�N���6�6T 䵝�V��Vz�RB52�5��s6`��4���(�j��6~ʼ5%�����@g6:�4���3��Ͷ3g6_�v�.}5�6��4��~�^���U6M}6�����,�5��A6D
�6a�=���>����4B��6��6�Fo5�j޵䤌��µ�u5t`��JT5�Z6Qs�5�h �/�6�ڞ5@ҏ�0e��X�h5��!���5�ϝ�J��6���5�Ѩ��x�6�5c5�wt6���50B�6�#�5��ĵ@Q*3��=���66w��o�k6r�5hU�4�ެ��'���55�}�	A� ���� 68����߈5/�55*c6�i�D��5w�V�����6ʵhZ�@lA�95��av6d�f6H�y�|2�6z3���O6�@r�7���|���vU̵}6��y����w4񡜵l��5�%��Iö�q��e�6��6a��5�R��Qm4��o���(4G
���4d����6o6t�;�G�;x��t�+��j�G��6�ĵ6/�>i�:�6̇:7���_gm6r���J�6���5%슶t�۵H�_5�����0�547/f6h��5�ia6O6ȅ&��=6��
����6t�76�i��F5����׵���6x&�R
�5U�h6�6���5�-�5r`�6jh��d�7&��6��5��5dx���\��P7 L����u6���Nl�6��o6ت��@"���;Y��]5-Qp�Hsn6�[6��>� �2�����ƈ5���5��6�t�@�I6�w���]�6>��:,�fHx�y$�6��5�E5�D��j(u�Uz�6r�	6���6��M�T�6@!���3h���6�75�:�5p/�4(�.���5�(�A3M�|ǐ��ϵpn�4oj9��5��8�63�,�`.�4��07�hն��Ӷ�7]��ߵ���[Z�6�s� r�c��_
��H��̡[��_�2/����6V�$k5���k�M07���ܠ�5R�Ŷ�~M6�=0�`Ȍ��_5��5+����C�*e15��T4�,ٵ
�\�7L�V's6g^�5��4^ȵ�Q\���-���5�D��6bp57��6v9�5��+�D��V� ��B鶬��5��6F�6e|a�\��6@	6Ȭ7Gƍ6�lN�g�^�l'60/6G�Cl5��6d����U�fa0�ǣ!6e�5e���,KA5�)H�^Ɯ6Ή5t��6 0�5l�5 C6ֲ
�?�4*�R��6V�8637�2��O*B6K��4�m��cض�:�6�d�������W6 �E��!6[�6oxV6��	���`u��b�v6�t���B�5��ɴP�q4A=�� �5�El�:��� �j�ْ76`�4���5�ƶ�v4�6�(������,��� %60���Z�����?6��*6�d660ó�Rs�6�Bu5�u5ض�6$C7Ϧ5����?r��Q?6�,�6O��ࡵ��Q�SV`��۴�^��"����6��g5�63S�6�y��n��5�4״4�z6��[6��z��ɇ5I.���b6@��4[ o�/��5Bح59��������wD�6v�6��U��]�����=�6����.̶�-�6;\������p6E6VMM��iJ5�@����5�ň6��6l��Z|�_@�6@v6J䴆�I���f56'6�����3r�95��ŵ�v5���<��6�-2������4<&޶�z/6��ڵ�c'6���4��P6@�p5�v6��$5�O^�Z����6_7�Fd5,貶䝺6�=�6������66@�T3��=6�
���Z%��Os�譄�Q�7jd���q6&V��wN��l  ���7�(6�����4ޱ��V��6/Ֆ�sĜ6PU"6$�y�<=����^5n�l�Hgյd�	��Kݵ��6ܸ��,V7Զ�`��6�O���ٴ!3��|T6y�?6pw�4�gR���A6��6����䘵d��4c���P�3)颶�) 6��6@�35��*��0�6�.�6�(f��"_6̢�X�5L��ִ86���5��#��%5��4�ߍ6 ��48�@�5^���3�v>5X���8C]5 7j3`J�3��Ƶ`�ϵ��/6���� 2�6�����4`�O���׵桷4 ���V�*6�b���� 㘳�ٖ�xѳ�W���g��5h�ĵb��5���Nڵ��2��|�5�l���;�����Q�5�[�5"n�6���5�6Ǣ�����Ƅ̵~��6�a ��[�4[���G�������Fx6YRC6��Q� ��2�?5״��!��f�5�yr6���6p�4<B�j� 6Fw�6��6`t��cG6�_��3H����5 7�5p毶���6\ζ��fK5�
6�ނ5f1ֶ�P�6*k�4ܪz�6N��PI��t/5%�5@�U5�AD6>�
����5�釵��	�����6�
J�|ݒ��d�5�]�h���5�5d(g6n������5wƵ4x����6�1�5~�6�Pw�64(���B��G��B�6�8��ܵ��6����á6�����xa��]�6�o���xI�?U�5���O6��������6��6n<�6@̳t�O6�p'6>pz�_ �9ǳ6a��6�'���|����O�͎��W�5�����2��6�t���56���EL6n9���o5z� 6�h�5��6�ѻ6��4@7�EI4�5�5���`��5߬16.�6��(`^5Pކ6��
6�6�w̍68�%���>6!��	����J55i6P��52v�4n���'6@��4�׻4NVY�$,�5 �	7�X4[L��H[J���|5V+Y6O�6y*��4.05b-���Έ4���4;�5d���;�5zZ8��vd��*:�_�%����*�5���5��6V�5!��n4�6������6fכ��>5o��5�����6+C����6׶Ҷ�֒�
�
7�� ��oԴ��3�@lp�����a�6�{�D�p�!�+6��V6xI����6��I�x{�54����f�6�tz��X|6�C4��q��A洈`�3��C�,�5BI���6�6���6�N�����5}����ʶ�1D4��s�6��6�W�|�6\:6�"�5za.6GtW7��x��'��⤵<.w��4�5|E�6췄�B)�4f1��\��6h�<��ɴ4@s�����5!�6�� ����5m�60V<�<�5T\��I�76�����6.������5(S�4/q�6�9o3صU���w6l�O6�~���h6 �6sԙ�f8�������"��$5������5E]6�5�1�S�)7[�¶'%5��-�@�[��7)���f&\6�1����5�99��
��G���o�5� 6��ƳK-?6��8�5����5~ʀ��������#�E���d/��&Es�J����5�f5^�p���G6��5����r#5�▴�?�5��0���5�
�/�R���~5������3�F60:�3���5Ȱ<6L{���06�����>�5��s6T�-6F�����5M5��"���9�N�6����:�
6���3�W<5���5�鶵76�ņ���D�PG�6���
@_6��ȋK�tތ6�6BQ6~n���f6pu�5�uD6�oE��%#�ę�䯌� (5(R�5]�F6��y6iѵ~06���T�?X_6MD�$zk�&_��\pl���66�=Ƕ0��6���tXy50%$��w%5���5X����7�j�6��)u5xƔ66��x�5��e6tk�4ξX�����dڴj�(|{��?�6�Hd6ظ5�=�#6ࠒ�R�#��E��Z�t5`�����6b6�B�S6�Y�5��ܵ�/���W5�:J556w�6��&5 E(�v8ݵ�6�}b5�}��@f85 �6 ��<.��%� }��T�5 Ť�(�%����[��������"�n�l�6��q6D�ȵ��H5�����Uܴ��06}�õX�g5���64l
6��µH:P�L�%5fb5h��4T��5�Ҵ�Cs6�Ե^h�5�d�5�<�5��"��{�5p挳B26�,�5�XL6o1�6�V��Y�6��)��n���P�6������6�^���P�5��6(��6P��1�5�+�<�M6 U�D-
6'�m6��p6����Ħ�5�g6�X�6�/�5����	64i��d�&;6�JW��&�4�M�6<��5���64�
6�e;��/�4[����SS���u6�'�M�6�6�5�8�,6 SX5 x�:�6K\̵�"60���H4>0�\#�6۪�����5v;�5�e���v��V"��A�5����~7�0�D4���6M;B68Fk5���Pp�B����u�pn7�m�4h���0ϋ��d7HJԵ��b5P�V��\��| ��a06�ċ��c^5 v���_��9�60��Q�6�f���7����E��)>6�'	6����\! 6M��vG;6 �¶c��0�50�I5�Tk3U��5���BH�:	�5��8�g�6�4�B����p� 6�O�5�͵��δ�B����j���i�E݌5�46Ќ$6����"�&6g��1��P54�紴�6�C����6~�6�g-���5=�5�ҧ���J6�}Ƶh����;5ޠ��E�6��5J���I;6���5����d�6hU(5$��P:7�V�5Vy´Q�˶�s�6W^5�B4�i�N��6 6|z��M��I�6��Ͷ@EH�r�=�3��5��+�<W6����r�ɶ�<N6��%����
p7@��$a�6xH6��Y�}y/�p��5 Y׵=��x�5�����,��}��WM5	Z�5?�54����c6:�a6Uߴ6�M��\Ñ6��6`[�3 �
�5����B	6�;�7C����5��5�`��
�����6�D�6�������6Dº��rj7�M�6�3���~7S�3��2ӵ�h�5-Nx�u�F��n7|�o�vrv5�`�6j�b��W����F6X�⵩H���$6�_�5�Ն5�0��$6leг���5 \v�A��5�I(�o�ٶ�c�5|7
7�<g6������� 7��j�6騶�N6p�3� 6�gO�c��wl�H��!��6�c��6vj`��%��L!��ߔ�6���68v�5!�36��>��2�J��5����Hq�6�6���5���4���x��6#�;6���w
���+�6��ⵔ�5��nA��l���7��P��+6�lص7����� 6w����%�����G 7�ֳ6<���~��X�56�"7;���`��096���6�D��x~6D� 75�5���k���H7��b���0����6t��6+ͯ5�����$��4|v7��6�1��G��6\��6Y�m�0?65�69��0��5#u�6u54 V6�t�6�.r����4���4���(�G��f6�`]�[5�6f�˵l����䵖�6���4�t��6�E5 �^�`���p�U5��ճ@�u��S5������d���`��5�:ʹ,|���%(�0���yǳ6��X6���6�*��$6Lg7Z��.���>�7�G6�z�5;�5=�
�3%7��6�C5X0���6S�a6���J䀶h2�T�n�^��jf��.��6Ԫ�5���Aw����6�-�6� z6�6�M��5�i6�������6o1϶BT�6��Z7��5D�'6��V^)6&��F=t4E6{ �����=$�6�74��R6Z[���(�(d�6n��6䕲�W���aE:5�7vcK�2�x�NK����6@0�4�$6~�97�E� -���⓵��@���ȶ���5J���i#7�j*6��4��2��r�Lȹ6��U6�Y7�Ϋ���*9��K��h^15�X~5|>�6��F7���6"藶�+s6�6E��{7Qg8�#�ֵ�����|N6�k 7�w6�'7UW"��������6�(�6�0��*7�Y��;�ٵWz7��E6���54H67��,Ӷu5�ȅ�������"`�Dm��7���^��6�MH�
H�5?�T6���6�.����r�"����e�6�L6f��6���6V�6Ô)6�|�6��;�~S(�h��	C5�R7����r����������6	6�\���_6�i�Fӣ5� �6�6�5\�5ލo6f�6<��x�5�qǶ���$�3�r��6��дH|���5��^�l|�5�w7eZ������oTC���봎y6k	6�_&5�oĶ�o1���	7�/߶|�6��ֵ�ߖ6z)���;7X]K7 %�Θ�6�w�6�̅5��13�"7��6����� ���7S��Y7�6�������5���Y�6��|6�����,�{?������6Ӓ�ʷ�4��6���6�+�6o������۫g6(���p�R�pN+5 }��{#07�%��춲�6W���^�6
���`�n5B����5~Q�6��6�_ 7cF6>\��;��6��7�|��7���;5ۺ�>W6^�ʶo*W6_�86| �6'�7p6�~27x��4Z�R�l�66�o,7xb��@��㍶�Ь�F�27���S��xS 7�ݍ6hs_��hǴԵ3�j?�6_��M���N-�xn����6
!��,@�6p��6��j�ƚ�5�D�6��6ש�T_6�#¶�,k�V)�5'�4�VʵN��69�z���4.Ɣ���5�D7�� ���5�}C��S����6VH06`s6�=�8��6��ŵ]�6���V�6�6��_;���6�
V��%��Jp5�_�⿭52��6�N�5��Y�Mk�5��63N5@�5B�ʖ�6���6��;�>b>����6I��5.�R� D�1X��DI��8K��+ �܎�5�S�6��7�"�6�1�6���4�3R��̮5EF�w�]�J�g5�+6 D6��)6��7��Q�p〶*X6Ҍ�V��� 6���4�����=��Aۡ���4���6�]����]5�Kf��t�6�5$M�n�6��@���Ƶ�� ��6T��6�̒5S���H��(��6Xn�6o�q�g6ܷ��]�16��6c�6���=jO���6�و��6��5���:�6P��6�H�⚪6:[:6M��6�	)�h�Ѷ�U�6�m]6�{�F�ܶ�5�e36�q*�Q
�4q��@�_58���Ϭ6�"�`	�4���>~�4��	7�[�4�ص��6��)�\y04Nz+5�b���96��7TiM�J�P6�/�5�p�����5.k��5ګ5�A����6�ӄ�*�6t�6���6 ���!���c��e6xԶ��5��w�����6ב�56i6�]����6Z��6��:6�6�#6�B�׼Q��� ��PF�U���6"~յ8�X5�Ԟ�z疵���68���-R������\6�x"��c������T�M�8)
7�N�6:��4���#�6�b��fl�6��5�����6V�6O�����5�O	h6u+D��/ӵ\c���6d�5@�2l�z�,��6]��6��5n��4~�60k��vr��Ͷ��4<��5�������5�#�6�?�6�˘��@.6u�����8��5�
7̅[��e|�x�z�{$���6�p�=2���g6|�5� 9��Y�6X����35\_��X�6� ����+���.7��P6`%x6��T5��� b��x2/5���5N/�5�B]�Az?7\��5�(�5lc�ll7(L�4���5���4��*M6޿6PF6�l�6o�g���5WÒ6Pn/7ڂ������ ϩ4l
��U��(���b�I8D6�w��g�5L�6� 5��(�)�~���6V9��>u�5~!�6f��<4%���6K�����6���O}����5��|���ֶ����)�q6��5�����\���с����4#�5m�96䵗4��,5�ڹ5�s�6�[��T�5�L�������o%�5�6�!S��ɉ6�0�6��6��1�0�#�L�|�|_�4�3j5���6V�6 H�0��H4Uhx6���4��~�v�h:�rs\6Ao���Xg�J6+*U6�ua5�*�Kt^6b!{5��H6푉6�`J6��`��Ù��
�6�E�5źh6�J��"B���C��
�>��6_~6�l�|�Ow�5x��`�z��� ��Vv�52�77�����'�5F�ȵ�+r���06��6A<�5�=C54�6�ps�6�"��N����a6���dB16H��6�S����=���7 ~�T�(7��2���3qHX7���3����bڵ��6X�Z�����rF�$�����|��b}6@�Ӄ������44 ��
к6�`�5X�+�"E�|���7l�h׵���5DJK�XT,�I626�}�6L�$����6˰��p������؅ȵ��t6.(^5�hb��}65X�6��}�5�v+�De6��6(�ĵ�6���'��*�5Jí��
�6�d{��߿5kB�6��x5�S�o"5� �x��6�+4�9�5[�Q�	'�6\i7'Sʶ�k66��۶@ԍ�8ڄ6��5���6���8�6�u6��#6�Q�5%�5�?�4-�6T��|���h�6�{����E7Iο6�l���Ե��t����6Pɶ@�{���74�H6`3�4�/���R��fw7Vdm69�������056���2��6ŏ�8M�7J� 6p��4�����7y��'6x��6mZ϶͚%7v��6પ4x펶[a}�20��Yo:7Fu�6��.��<�7g��5�_���� �i5l���=��6l�ɶ9U��ӓ�N�<�0�I��ޅ7.G��` ����g�F�7 �'2r�7���68
^�?��6���I���ΰ�6�*�6"m)60�6�{��� �+���׶�7ڰ��Q>�]�W6ஊ6�[��ͅ�6�5��5�SM7�)��Ѷ�� �-5.7�Z���5�⦵�m���'���L���s��+���6t7?���a��S4��Z��`���1H��:�6>_��n.ζPy�4��c�&s�5b{7↶ ��6L��6���|��5�}���W��.��6�357^*�m����Mp7�2^6"�ȶ�.ض�p5�Gζ)67V�6|Q�T���'�Ś��C��9���Y�6��B7�	6�C6B��6�M���Ū6����T)����6��ֶ��.7���C;V6��6�.d7�+6�Pg6�ty����6�@s�8��7.�5���=��a47�Wb�-쭶��64�¶�9�6`��i���qXJ��Ǖ��7S	6w���$�6j�6
|6�E�6�R6�^���u�6<K8�����ڬ��E�5���� Q�I=��A�[6w��W7<(��{v��s@!�K�1���7�wD7^㍶�##7�w���V�P�5��4�5#��Ny6ɧ[��8�6z�7�3��:���(}����=�V�䶔ܽ5�s���!7�O5�(����6� ���g���5ӵ������W7�����B��5�۽5�k�4p94W�%6u�5|d�Q�� 0�10�~4@n�z�5�S6\$��
�5l�u�^x��<T66������H�ڴ�_�5�N+�����6�q��S� _5?�5n.V6 �ɳ05�}#��d���a��5�0gb� 8h3 ���b��y��`X����Ț���I;�|�,5������5�2�]޵r[I�p��Jg4�5(,J�AX~6{�ᵸ }� Ȇ�ۯ�6�~�3�������6'�Zi �f�S6}6$����̲+6�'�4R��7{�5]��P�j5�`�H�6�S4z�ݵ��3�T�4�s@�,�|�-��K1�5p2�4����8л4�}��&*6���4�IY�r46�� 5Sd��D��� �1��:��0zE4<6ֵ���6 oǳ~:6�∴-���-���u]�p6X>�5 e�G�����5�X���3��5l���Wm�T�6�'�6�%$��^�5�<=���&5�����	%�5̛6 �����4�A76|�е� ?6:2�5#����
�@6t�\&m5�⺵���f\6�=��J#�� ��#Ρ��~E��+�^����uw6��4���5�(#6`��4@˥4BÈ5~�}5vt(5I���ƴz��5it��|S�5�R��6P���h��4"�46�_�=06`@�� ,�y^���ǩ5��Ƶ2o6 �94.Y�5d�g6�r6�͵c��5 �޵����.�5�Æ�����D��h[�@b�3�]x38�$5���4��>5�4ƗI��.�4������>]5.�ݳ��5�A�����)��5(��5 � 4,����6�X���_5)4U'����D��6�5R<u� K��\$6nX�5���K��5�ⶵx-85�"�k_� �4�ȭ��\���&4��5��6�]�5�S�4�7[���5���4X�(�p�4���zK6�d8��.6�ɵ(׾5(�R�2� �dji5�zJ�eõܝ�5?�f5$�س�IԵ�$ 6c�f�����!�"6��4�D6(ځ��)��_#6Pס5'�e�i�6d&6Ԁ����[6N䀶I#���[�6�]Z6�a���6�@�6� �4�![6c]�6�o4���(���$���"6 d����6?�5�_r4��_6ZrR6^�rj�5�6JTA6}Ɨ6���5i)�{��h��4F�n��o�6Ϳ5/��6n:�b�u��6�6&o�5;� �f5A.�px�5�O�5���6#�䵕G�=6V�<�b`g��C��xJ���J5r<��W����h�9x�6{��5fn	�c]6*F'64m6�(�7�6�\����������YK��H�5բ�6\�
6�P5�I5�,����L�'6�ՠ�0@�4��-6��06�6�+46~Q߶P �����5��6��1������ۆ5�$6���6:D�6X		6�:ٶ^K�4c��6,�I���5�Ϭ6��]6�/�4�h6�����p6���5Fy��}�5s7[~��fZ/4�f&6�+�%�����Q���455�}�l�65}ed�=o�5U�6���6w갶�k�5e�a�D z��^6��G6\�ô��6��6���� ̶��|�5���4��6@�6.�O��ȶ�j�5]� 5�w�� v�<b&�ު6�L���C6S�z���7�5%C5��Z6a�6�V�6�|���P�6��[5�a6�9���>6��5�p������N6�C(���7���>|Z4���j�w5�v�5��7ϗ}5��3��U�*���� ��h״;�+7�u"6��6��R6wR5(À6W�5���6TV)6hS´���6�$5�/Z61LL6�[�6�?���r���6��K���06��j6�n6O+F62p5�3�6��6���51텵	�P���7Aע5��X�8Me5˸�۱t6q ���~ɵ�ǳ2����D����6��5��5�ȶ���2�4����U_6b�6nތ���6 S�3I��57��5���56�4�ә6K�|6�ޝ�����iJ6��O6.DP��06�cz6|��5 �������&1G6֘9�T})�.\g����41ʀ5/_M�r��6��
5�,�6�Gj�n��5
P���c�6mN����5�H6�)q6Y)6;�H�6hHN����5,�4�ʞ�Q��6��56u5ˏ�5�m6߫\�m6 k3fKy5]���6?��6�T�-�\�5�5x�4�4��[5��6���2����5�eE5���4z�ݶ���5`'�� <�6����˅�5�)���?06I6^ɑ5R��x+�6j:K��T�y���@涻T|6���4�8�6���Ei��5���5��A��'6������� ����n<5dV�6  
3��v��f'����M긵KO�5|���~G{5_ɐ�*$x�VM6��5��[5�L$�h��j�$��*�������7����@�ܴ�(G���z��xc�)n5@w4������d૵|�58��3X��K���F6�4��B���6�\cx5����(}�4D�5��?5�y�y�Ԫ4�D�4�?5��Ƶ�����,5h ��J15#����JL5 b4���5�%ԵE:صR��5]�6 ����57v�	��5DI�5F2���3P5��5��=�`̣2Rm6_��2�5?�5���'P�^+6��m��K�5�.y3z�5!۵F�ĵ��6ݖ�5�L�6�;6e�5�t<4���$�$���|��4D�� u-6�6t_4�f�4RB�5d�k6���J���c�4�TX6���5%�'6��5�Q<4��S3��6 �ݲ$��5�H5�����%��0��6`�����5jZܵ��5ηԵ�m嵀�0��yx�����Iu��j}6 ��1����wn�59�U��,U6ٺc6z��5��T6�u-�0&v�9.ѵvor��%=��ra�Šb�=����o�0� 6���e6 Cܴ�b���6�Pe5amO�|��u��`/���@�5Jfe5@�5����<�:��~���h���A�5��Q���5�16f��� 6�{@5��W5���I��D��eS6�s��2YĵD��68�7HA)6���6 �g4��&6X���8�6�� 7�ض����T$���Ui4+��6>�6Sļ�pOڴD�5"u6 .��ԫ6�5��7�5g�6�Y�TE����E6���5:li6b�_6���� ��3���<�6�����w�4`v�7��5IO� ߣ�QJ6k*�5 R�J����N��%��{c�*�<6�A@4��#���6h�쵦+���ф6�%����3$�J���l5nB��3,�rT�6Nh����6Mߑ6�uW�r�ٵ8��4�F6^5f6���5V�"��������YHr�0H!��t�5���5�%״|{�����.��5fSs��16�̓�-~����Z�l$6�56���5r��5{���5�C�5�%
��5���6(����	�`�6̓��G�5ɱ6��g6жw5'��5�Y{���A�J�26̨d5��/�6��6��60��MS5 p64=�����5���k�6��6�ؘ��=26ڜ��@���v��fO�~��6*����U��56���5�UB4��>6Q��6���5H�1�V������51F�VbZ6��W6z[6R:ᵪ�0��u� 뱲�����J�v8�6lDr4���)�6F<�5�4�6��6��(���6�� 2���36���k�6�1���5�و5`T��/C6V	5P,4*=�5h�Z�0I�4�O5�΍5Ȍo�BiV6?�u6��5x�6���6��ߵ�ѵ6N)�'@6��Y6
��5���5�m6�n�6(�PO޳���6_�ݵ|@�6��;�8B�5�:95\3 ����Ã�5�Գ3�:X�譇���P6WJg6��O5J�+�w'ض ��5�6J�_���&5��5
�5r�5W��\�85�>��#H5�0P�t7��9�Q5,;�5 �����������v����5��ҵ��5���6��ִ�5n^6��5�!
��^R��M���4嵤�6���`D��T;4�ᵮ֞�J�$��S6��4�17��񾵴�,5''���(/ܵ��5�qJ6�0�6���!�d��<^�4�q��� ���o6��&6�V�(��4 B�5��'��~46�Z�6���4P�6�6�h�5�B��� ���5�u^6h����6��׵���ό�B��6'��l@�6ZIY���U�p�.��Y�1��F6fn�68p�43�]���%� �������C6��6u�6����D�d�)4Y�}5h�{�yԞ6zc��>�5��5����6`n��7�A6��#6M���?(�~ʚ6����wη5Pw��Zv7�w�/6uB�5�%u��0�A8s6`�V�K-�����"#�5�!���暵T�4��66ZP6��S5�]�5����(����6��j6�8)��ٰ2$�76%�6zQs��P����B6\
������D�n5�qg6�{��j����D6,86�$5<vQ4��<5!S&6��/5�w��[�6��ε�(���{]�Fy�����f�^��8;6ʀ�6��>4�Q�5n�X���� ��5̒�,##�JV^5d��}4޶�en��4�5��[�@A.�|�6�-׵�lx5�68�ȶ�%7��6pTj���5��絤q�6����Y6�,�����4�G���־����4���5���4�ܣ�`�T4 ��ܮ6�6�~B�hr�B����Q����6lS���[*6�K6.5@��}ᵷZ	6���6�x�4�Q5�Z����62���<ò5O��dN6�W��93H.96���5���HX���06vE(5�E6�tE5d+µ�kN�>p$6��)���6F��5x	A5��p6W�{6`o05�P6��6̒���ۻ���5nf�50��5�O�Q��$�4�a4T��6�J����5�d$6L�J�� 6��:)鵁�6�0"�t�V��F��癵�/���<�5�9`6`w4LF�5�j��CB�6Eo�6`b�� �6۪5\�6��𵆤X5��5����C����`�5@�04��>��5�����}6�mζ��5"�B6�7��]��2Q�5d�*5�_25`W�5��8���q6`Ճ3(�Ͷ�Wڶu��+�6j����4o�6��^�0ʺ���&52ە5#���fu�F�^����5�զ�2�46��P�M�C� �6l\6"�60W�5�V6�Nw��95[oe5zlB����*Ƕ5!ǵe*�6}P}6�͵$�*5�k�5I�(����6��|�����ۏ�� q�3'+�:���;�54X��8�g6�Ei4nHE��:L�/bi6db�����3�Ŷ�Z6�[6[�5FMX��e 6|�8�F�.6n�ô�J���lP52� �r:�- 6:%�5������6�;5���5#�4L�B��6����Mk��H�W6�,m�J&6�|0�w�4�[4O��4E9��z}��x ���х��L6�ґ�N����Ӵ��36&c�5B��5�}�������:V��6�����
�XĴݖ5@ݜ3���5�5F��`�5i�?��P�5S�5���E6�.Z��`�5~/b�>y6�\H6�aW6XQ�4�@�p՗60��eX�5y��3@Jo3-1*6-����t2��||�k~��C��5�/|��6��O��~T5-��6���`�;�r����n��6��{��-9��җ6
36Y�5�x1���(6�~C�� 	��* ����5Ƙ<5���6�T�G�Y6-��5fY�5�p3�A�5;ô@�5�U6@K�𢀶�\�� �೏��6��5�1��,�ܵ|3��m
��oW6�6�����Α6��ǶЅ94����T%o�H8�|+#5{=56���0�Z���*6�g9� ����2��@�5`%34��X�6E��
���m�4��v� 6�P��娵!5���5 ~'�|�%���5��5N�H6���(���$��5�%���ϵ������~8��߾5�G^����<6�e64��Q7�����5!7p�U�S�5�`d�hߵ�D����|6T�O���4��6NC6���6|	�6�Xε	��� ��,Ƶd�6�w��x�õ����H6�n�6�4�6�(�5#�6�\�5:��6W��6b钶��5�,�6[cI���c� �Y2ï�5 %7.��7AΊ�Va6*�6hO���PN5�h5P�5~6��z�6H+&5I06��5�g�� �5�h6�נ3zY�5	�b���ĵ��66�jX��Z���W�����6?���p�1�E�S��
�� G�9�6(�5�� �4	6�:���4�ʵ�.�6�5�6���6������2�
^^�&�����6�_�b[96�t��JK��û�f�6���6������n�*?Y��
���e�5�Z6��E5�5���,o~�����Nw5���Ͷ�8?6�(��0�}��m>5r�7 ļ�r����<���>��;�4�L5�µ�ͦ61��4H�5��ֵBe5��4���� 6��ȵVҴ��������V�5:aP5�}�5� �4����`k�3hTK5�Xg����4�ش�D�5�b6��~�V[Q�"�ε���xД5�T����6�
6��
5Q1�J,�
Uf6�f6����ާ��8��GP�.Tﶜ���ц�6�c��Nd6v�$���;��X6�[�556����	�5�Ƶ5[F���\6%Gd�i���!7���� 6��6ԑ�6�_���>6\S�6hY68_�6�k�5;y,6�~��|�P��6���<J�6$H��"�I6���3�b6��34C0v6���3 	E6�[;���#6썉��b���Yu��:���������5��6	��6�o5푏5��4_������#4��"�16�!���ǃ�6�������26�h�6��R��ʥ6��<�u5j�6���U?��z95��6Z^�54q�5�#6̻k�h�5z����m6��Y6��6����~!�6T����U7�m�5�φ6�;��6��6<r�G��g^�6į����6�`��5ў�6�C�������4, ��
�1��ڬ��Ы��9�6zݒ�����V�'�6�Գ4[���+����6QI�j��6���~�7����h �54O�6x6X77׽�@�4F6�5� 7��65�]��*7��P�cR�6d;7��i���e6��g5���68�6�E�2i���&����6/������ ��6�O�5���~���p]��P6H�Ҷ/������l�E6>��6��6��5S=�����	�\6�z<��s��1���5&��h�5z���ȵ�Pn5��7��K6�Mֵ~ �5�ҵ��8�4\D6��B5lQ 6 &t�L?���"��M\��w�6U6-6 ���P@ 44�7��6�N6l(���p��m�6�m�6P{�4਌�t]�5A`����
6`ǔ5ͭ���d56��]��8�6�F��_&��̶h�6���5��Y5�_���µ�t��PbE7x66x�6.Q�6���6���5iV6&6�6r�4�&6 �z�	+Ķ漳�����]?6.3F����6{%��+�6�!�6iɘ�n$��5ʎ�ǀ
�����TO���k�ʝ�r�Y�Nrr7���6͹��7�5�7����|`�r��5�%�6�;ζ8伵,�R����4��6���:Z4@ׇ5�����p�6a�6�6M���	�6.78��4�6>���}��@o���)7R��(;9�鉁���6�7*�J�� ~��������ڶv�6��6�W6I��@a)�Tֵ�D�6ʗM6^%G�te�6nˠ�v���A�1��+��,���q4@��� � �4�v��l�6tZ���Fg6>Hq�DE|6��6 �16Ђ84$\6~��������l'6�݌���G��'�6�5��Ƕ�~�6���6�a5W�P6L���J[6��5]��6��6��Y�k*�6��'6h�F��=���#4��5�J6L�0�5P�̵8ȵ�����79Y6e��4x�dfp6�78��Bٶp#<�w7���5H���6P��x.t44��6��6x�ֶ�]�H&��\T6p���>�4��� *4��6�x?��2�4/�Y6��6@��5 5�F$��^���۰5t��`J�4�ն�E6��R���� 26���6���6Į6�Zن����6�Uϵ�߯61�J6��-6D�N6>��@���l�ǵmZȶ�0ڶ${��lή54Xu6�8��
������Ʊ��W6�х�����|�A6�g6@��PG�5D m6�`Y6�d�lĶ���4�["�Ǹ�6��6�\�%3���K㶪EC���5�N�5@k�6��ɶ�o60\�6 kδ�6}7G6�5&5�86RIo��� ���c6���5Ls5���� 62ݞ����5�Vn6b�;6��=��A�5���4r�6:��4]��6V�4�dǵ�����v� J�4a0�P;�4)w�u0�#�:6L��6�,ҵ��2������䶽;K6�·��8�6�.6]���1�5��16�k_��Bg�׽�6��\1ٴ�2ҳ� $6��)3�L6a��6��5R�*���b�6.�	��x6�!e���Բ<w�5�=6�j��,��#���n�6U�5gz�5}g�5@��6���68�5�8�42������8�5ۍ���6L�j7?7�pϴo����@8��2�6H=��k8�A-��)�6�Պ���̲�3��$��6�m�5��&��0�64'ᵊb>6��8�k4o6�]�6�~��m6�dF5�I�@L�ٌ�6z޻�|N��B��4y���X+����̀��&�7%�}66�T�6��;pS�{a������@�,6.����S6!
5�� 5D�6x���.�51�I�_m6�~�5�����篴�9Z6poB����4⺋5/6�5⏚����SZ�8���(�H5�ګ5h( ��O �2׃6|5vc��t�6��F6NK6�_j��󑶌�56KA��0��6�+���6 '5�f����"�,�6����)�6lڶ��/���7�9A6�'46����ؽ�5��6�A��$+5�[�6�@�6���~�	7�/���6����A>�l��6;|>6�a�4���� �/��ߤ#6��e6�WM5�V�5���5�܂��R�����>�I��L"6�4�z�6��C��%}���6�O�5{+7��B��t��ƭ5�������'*J��������RB�6t�|�D<���y��G��C�����5�;�[=%�y�R6]�ܶ3���N��5�v�2k�X�9��6뚘���f6
�%6�^�5��`����o��&��;n6�V54 |�2X�=��ȶ}�,�aC��>*68��I�*5,�4�:�6�
7Л)�[>��K�7�j6���|9���Z���\6&�5���(׿5�n�4$���;�6��5�-W5�����մJd5|%��~�5)Ij3nI�6bܶ�������5L"�66-�6y7TW�@�a�q$@��Dp6@��5�.�6��6&�ж��6(z
�j~�5NQZ65a07���;�f��& 5d�5�|(5�ƅ��~	3���5n�_�7�i�R���p�5�|[�zC5���5)��6�$&5���.5c�6���3�|���/&�)�;6�6֧f���J�q�J�DA+��(��k��85�7?5�Ft6{�6\9��U�5��T4�+�|1q��9$6��6�}�Tێ�4|�3hrI6�6��.���"78��n�ߵ��j6��O4�/�5�$��R��$�o6���6�0�=vL�� ����K����k����Μ��X���ɜܶ���\n�4�팶906tGT6�T�6jiw�P�:��x]W�l���=F���5�%����4T6�е�^.6��4w)�5¶����5�m��8�y�`�4I��6V��:T����1�5d���鴺}��m�;4L-�5�,�0�d4�Oa��s9�(�46���5?�����5 p5�["��ҽ�D�5��(5�M���/3��!�9�Ƶfū3���5B�"��75u�6�E5,Z4�W�~�� �:5�j5���5J�6�SG���[X5y4�h�	6�et���M2)���M1� �a5�V
�4���T�4�2�5��4��/��S���16�ł4����5��5�5(���ѿ=5M��B�,�v5Lʼ5��4�5�>�4���4|'�5`����5W�M��Q5´���r2����G6��;��<����6��״ɘ���R5n5�Ԛ#6[3���_t48��6_�5��5��5*�6��52K����i���=4�r�5h��4�e^�ϋ50�?���O5H[�L4���:�����ԧ3H��M!���5����35�g�5�e2�lW�5ȁ�5�G���K���-�l5�(���3Y����5bT6���5;8x����X H4|���(���sϦ5�D?4W|M���Ĵ}y9����5U~6Ra�p�u��5�ڬ�zm��iC�ާ۵M(��]�6q�5�/L�ą���nݲ`k=5 ��4l잵�������4ǚ��z��������܊5P��3�5�v�ʹ1�~�52=t5ɾ̵��5�sR���E5��ݵ��Z���R���t5t����60H6L��4���@����Z�8�>�^x|�� �4�G�4Deo4s05+yG5�5d���}��15�71�����5  |��ﵝ]V�� �;�3�*60�%6�Ls6�hT�/?x����mϙ����롵虥5*���/qE��V^��5�4FB�40 �2�P�4�-�3)+@6F8���˵��6"�����4�+�@g��]���7Z��R�5>����L5j.6���52Rյ��5��5k��5���5P���U�5��7��o6UG�5$_�Z�_6	����5�6���yL������L���q5��4�7	6�_��Hw�H�6��5��ܶ&+�6rb�5�o6���iR��:��5O>���p�6�sZ������
�6��p���4�I�6N{Ķķ���&6��k4��E�sZ+��ǵ�86�Ή5�Q\6F=�5�Եt@��8��3�a85��6�I����5��Z�Uĸ���6k�5���6��J6�4�6���6�1ᵬH+4��86|$`7O���������8yX���"��"���w�&��5���6u���_�q`��|6���4�c��k�rl���7,���߳f�a7�%C6�Ƣ����Ȼ6��6��ٶ�
5V��3�F36�����-6�=������L������I�!5�w�4�.�]M��"��.�66(Y�5W�x6��V5t/7n��$�4B�J��u�D\�<��5���6xm6�n(�)^�4�M4e�36��@���65P�55����Kk6��5�86[�7�8���Ե��*6��z�"^9���H6��6F�ն��
�֣�6_$ 6�rf6 8�6�B�5���^50vŵ��5���6#7���0Z7M��6b���uB6LA�5\�5�ʵ��ӵ.5;�[l5�5E67J��L�74b��6����f�hv5�7��a5���5h4F5�4�6t��*_�BXi5뺶��5�!6ڢ�P�7�Y�=�6���6�a�4Ij���,} ��%�6��	�6�̴�:M+6l�����/6@`�3�4�T;�5PZ#����-��6��s�^t6X������4pL� v�6@H��~�r��I��`������×��_�6��`6�H�6�[j��ը5 �N���6�����a�6F7 \�<�6�|$7����%�)�M�*�06�e��(�6���6��6@=D3^0 6(i�4sUQ��-6�P뵝W�6�6ۅd6����.h5\h6 �w�K�*5ꎶ�aݵ
��5A���)	6��z4�ϵ>�7*�Y6p/�5T�c6 ��Zs602+5b�56�۳������6�收p���Un66|�1���U6�y5`{�4㉯��1B�+T�6�t������v 6���6�� �n5�x��Ǯ6J�5�xm6��6�5ܳZ�vz!�66�I75�}_6;t���D)��\6��A6�&ඬ�6�-6�GY6��5���5�5��P�u5F>o���D�P�I7=�ն�n6�@����D�5$ʀ�{�^��E4�T^6�	�ػ�6��5ˬ:5AJF�䀜4�B�6�qŵ�|"6Э,5�{6G�5.�0�\�6��[6]�i�u�2�o��6�m��
���6���.6<�=�l��6�6�.5�����4�~�6%}����6p�д�0�4P@�5�{XѶ�6�����P'����4&�l��T�6�|a�h�5��5t͐6j��h��W6|S��j�L6d�6ª�N��D�6��B��Q�P���͵�ym�J�}����5���5�S�6�c(6xJ�5��]5ʮ���;"6�]����>�0~5���cf��@uL����%��6>���<ݴH�s5�/�ü5qr 6d�ݶ���i�6k,!6􀿶@�3@�k5��O6�"o6�lC5�c�5�h�5��S6�Ҽ�\]�5p�4(�����5`X5Sͪ6��"����<��5TBv5��5����*��5�~8���^6�u-5P�O5���6a���5�����6Y��C���B6��s���6��4�sB6��"5��5H�嵔%�6�#Z�n6���h�y5��H�G�P�)5T�x65h5��6,&�6tIǵE�,���	�a85��q��]�6��O�(��4$0S6��=6������6@��6�KH6�6na86g�74��sl��d�J�6n�5�O7���?26Z������6�R�5ږZ61(�5O������PB�4�.5�@6o�B���i6
�6HH%5�I��X�E�T�56�R�����ߏ�t¨6M��L76dGQ��È���62ps�F-V��L�:��6#4NEX6��6�ݿ62B�6�~5Ėc6��6Lq�4���#62k+��!�5���5j�/� ��6{.�����6�6�6� [5;�]�����U)�S�7X�36_Y�5����T�o�6[��5��5�\66�6�
�6l@u7~�5����|�6�o�-���o�9�H56�A�)6/u���T6�D̶�&6��6ղx5ր��'���߫����-�6,[�5X��5��öh*8�9��6�Ŷ��c6L5ɡ�� !95�@�z}�"��w�)�a�6Ԅ���uT���f�
�� &m4 �Ux�5�,��ײ��(N6.K6�햴6��P{�"�G5��ɵ%k6F�2�D��5a��v ^�F��+���[��Bĳyy_6w���B��4��6�1�X�]��6�a�J�6��6��e��76�a���`4�k7����ֽ������@c��<굼��6��C��C$6�����۶=b���5��5���wW5uz,�2���\5�������6(�k��޵� ��h�5ܓy6m	7����%����6�;�6B7$���<�Z�a���jbF6�W�����v���G8��2�66��6a50�� v6�t�0�6<��5�oL���6.�Ӷ�@5�G�mN4����6��E����
����5�P5uʒ6dҵ���6r����4,|��v�6�Ӷ�+7wț��D�����@ʉ2 #y3j�7�d�5��Q���6⌃�)o��x?�5@l�����5i��6g���[�5?�6�6 U4��ڶg�⵻�s6�K 6л����O5��4���d�v5��6��6Jۇ�Co�6)L2�ڂ�5bö�`P��pе|ᙵ��� �޳�Ź5��M�d��6�%`4�c�5\X7ټ����뵯�ݵ�c����
���5^��� �ɴB�R�_��6��[5���5��`�b����8P5)U��sӵA�p6� ��*���@�r@�5_ƴ H!4̧���&�5Ю�5�ᵨщ�JQܵ�1k����$ӴF�6�I���u��S�5�\5�_5����x�����6�绵�QеQ�5��6��6F�5d�r5R�����..�5��4�_�5i!6`Ӈ�ʦ��[f��}�5k��46� �58�_�*iH5aA>6�8����^�T6���!�H6D{�aZ6���Pk�5ok�4p��6�r���ܵ�y�51{�t�!6�&��_g���*���O��!����5L��a�d@6/�굥q�5�#/6�󏶐�6��w��365�V`6���5��>6�@����-B6Ύ���ݼ��x�@];�L��5�lm���;4�4���i 57.R5D�5ٌ��@P%��@������V')��|�5w���0$�4b�86��6�mk�Ӯ��$��x��6$F�5Dr?6������P�t�R�*�#6�l�`-�]�5��K���5��H3z�`6���6�,�5݋����5_�86d����a76��5�L��,/5���N���5�
k5x4���έ5<uT�6|�5n�"�d����4qa6�����&�{6{�6�H�5�/�6-��Ɨ�,m���6'[�5�x���P�o����4�S���fO������C����@�6��4
Y�44�4�O��J6	7�m��<�˴u5!��lCt����5��Ե�ly6�%l�$!6�����n4͵;��6��4�
�jF$6�>6��5P6��e�vyS�,xy6x��*)������rLW68������	j6�ݰ5����U��_9W6 ��2Dr5��x6gE{�lǶ��86����
4��6@�3t�E6G5Y6X�c4��{��+�6�l0�A�4����5U��6HM��6�5�4���V6��47��5���5��4:����M���Ѵ0ը�I-6�mN5�x����=6TȽ4����DR��W5�P�4O��6�4:��N�fN�6�&�6�1����Q���p"7JT�V^��0�`q;71|&� 9}�%iƵ�ڙ�-�I6�l)�[����6�4A6ҷ�����5�I�6���5�K�e!?7�������6�6YEE���6�nh����6�S
6��3�>�F�D*7����^x6�_=6P�k��lu3�}�6&96t:$�(�6�Ƣ���13��"��6j�A�k4�5�/3��hd7���648�J��5%��6f�D�Xv�6�~?7>}�f�K7�V�4ݓ˶�t7����e��b{�L����������E%7�z���M�5�p^6�6ҝյ�	��et6F��6j�w� �&R���6�Y����^����4&�s��e$7��7<������6*��������Ӵ��Ȃ����a�f��68��6����
���P�[�;�ooW����6:����6�Ҝ6������嵰�A�ݬ�,մ�Q�6�����@6k7�d��
Ds�@����6���M7�{s3�z6��5���v%7�G�x���r۶\�7��7��㶳޶_G6m�Z6ڤ���y�Tj�����Q��6��6bB�6l�
�І6�X�6Vg�7s��5J^�5~)ʶ8��4�^���I6��*�����Wi����O7T��f?�@3��ޛ�6��5,�25x���!6���6
o���s&����6`�z5�2�X�ն 6��P7��k��6⭴5�aw�,���7���5�ݶN��,�5�$�6Ի�5(F(��YA70t<�TT� I5��5	�I��0\58�6�Z?�<�~50P���j7DE�d�����R����Ƕ��E6ɚ��������1��z9���,�|�6���S��6P���u�����5"��e�H��6��[5X�%7�u�X>�44d��^������R	z�ݵ��ו�
u�Q*+7l��6���6lN	7��H�}A�:��6 ���u������Ѷ Nѵ:"���J�� 6��E6{�۶��H�/���&���1�L\7䀸����5����б�5bSg���T��5;_6�����I[�9,�t�~7`Nó��y�ƺ]6��6�p�5���l7���'7�Y47fB�5.�:�6���6*�赞�F�/2�����a�j5<�6rO��Ux��;�5'!�4���5�-7�6N�� �A��Xp5,X�����6dX���w}6fk7]~C6:&�6�����6>J�^>7t��6��?����6��o��o7J�6�����W6-�6�P 7��6�n�7(�6e��5xѶݤ�%}�6F���|�7���6��"6�)3��\"�8�7��+7�m �E�\�����r6O&C��=Z�1�µP��5�&�6@T)�n�q6��(��X⴮�����8�^7v������6���:�٥��i�B7y7�6�<�6�ö�_�N0�5E����K��$�7f�6Ӧd��ȟ6w��6����pN�5��6DŶA>{��2\7��¶�77QBӵ
���k��$�׵0����5�/4n
��� 6_�s���6:k$7��N�<�)���H6�;�6
�ȶޥI6��6z�5ᅂ6��^7���7w86 �_�t)���r��2�7�*�6�Ww�tbd���i5��B�z�ö({M�U�ֳ���x�6t�%6p�J����6ȳ7�z��޺6t9�6�u���T���5b~��V47��w5�.�y�6E��6i��6��������ȇz6d�T�Zi����k6b�6��
7�D<�J����:7���62}36"�*6�_�%gs�_�b�! 6�N���6�h_���5�~6
,.��!��"���"79A���46j6�{�6���5�ʵ;�R6ik96�p���5�����W���i@6����T���6HӘ5P6l5iޙ�o�5�B��Q�y6H�ôwb��70��58��Bp�6B�6�1&���65��6�z�>�b��5��K��c�6L�5,v���?05��6����жV36�n�8O���6D�7��e�,����6H��@�`��z�6�!+��N5���6R'Ƕ���4��7¡���#���l[t6�I5�@1�5̔	�R�����W7qT޶��6���� �c7�b27J�����_6>#��p�6���6
V���6��6�����p�>�`6�2�9��6���6AkM��a+�x�@���&��c�5�׵�T�6{*Ѷ��6�/E7XA��^?�r]7��)��uj���Ƶ*2-6��%���i�8_�5��c5�+A6�gö�r�6nN�6�P�c�f����6��ڴ�[�h�����5���u��V&6e-�6��7͵X��J6�� �^�϶ Ph5:��5��F5��7�ϟ6���6J�.��Eж���6�jM7�9�6���p�"���W6��?6��?6z�6Pk6l:�6��ضH6@�e�ޝ17�2"�
�+6t7�U5��w5�����4���%��y�6��0�h3�5�F.6W-�D�ɵ�A�6P�n����4��5e���
*�J�=6�Z6��o6N����ݕ6���r��6���h�﵄��6�
*7Ja7��\6#��X�7 R���[(�児7^I�Q7������$���]7ܨ�6h��6ޜ^7�6'`�6���7��6�h"���+����5���5��6p;�m�7��Z���W7ps6K��, 85ƍǶ���5 K{32���6<������]5B�f6�?7�z���}�5�,�6�����䪒5�:�5���5��77�J��=�6�8�7�`�6��6M4Z6�����W7�#86B�6A6XI�7d�O6���>(��"y����6��7Rd���c�5N �6�df����5���6as��4��6���6f��6��U7 �x��\6*�Z�<�/��X�6C��r�7u�ǵ���5pJn40,2���%7�|��J��6}���#��5������6��46����{�6���6P��5xN7h�76��5�<õ�VD�"fc6�-66γ-6b�5jD86���6E�5��w�59�`��5����_D���L�6 b2A,�5��Z5"Ğ6��6��Pp�IUk6 ��5�����<�:$�5֭5��ǳ"��`�1����6�6xĶb	���l�6��5�C
���964�5J7�6|ث5p,u5���5*�?�����6�S�6ݵ9�s��QG�ȹ�����6R_�,Y��J5p���v�4.76F��5=r��1�/�7����E�6(qG5K��60@6�@�H���i�5d�%��A6p0��W#��'��~SZ�2p5BE�����5�����3�Y>5奝6����=��A�ݶEr6��H5��@���	�����e6@7�5�����@G��1��@GE�P�6({�:��6�,�����6(#$6��o�V|�5�56���5�3޳5̶Y#� Ĝ6.��5$j��xb��]��>����X6��b6��u6�i4�ĵ����	7$��3 �7E��L����5��(�^�o��a�5.�4�d�5̈́#�2Z+6C�6.���עH6>-%�Y����6�q�X��5'�y��	����6�Ge�Nr6.?R����6��@5%�V6���� )3z)�4�v����6]����{:�$�x�P')6�EN����5�796��O���4H7��Ъ�.�4��t6W����y�4��|�WQL�p[�6>;�R�6 �6/V��)���3S��7�����E5�!��l�7�.\�����6��?��o�5O����6�j�6�s�����Uh�6�7�5���5 2���&²�4�6���5jϏ6n�6d�5]޵(�5�X6�Md5�͞6Jxض�:f����Lɕ�Pb:��3�4`���%�6k��6�Xƶ��6̣ ��W�5@T�6��S�̕�5H}z����.�Ǵ���6�.~�0\����
��oL6$�/6�\�5zj�5N�Z�l����6������6s��6=G��*7*K��Xq5�U�!�5�� W�5L`�5J�޵n#�4�d$�f��X�f��SQ�"��3 |�4�������4��9��$#��֎55|�6g�5M� �5Cƨ5/�6��ɵ ��5p�4`�޵���5 =��Hw��฼4T��5�󵴂����r3(�õn��5�n-6��D���i�-k�5s+6�4��t��4�*V�16����L뵀�>4�3;�N�	6���񀵌��5���5P�24�(	�(Q��`��2���ܵ�x���5�046T����5 �o3��嵂��	�4@@1�75��6I*�$��ZCG6�+�5 �a������B2���d�ސ����[4�ֵ ��`�س�y��U5�
}58�B4��´����8��j:6`qG3��K�@y5�j&6Jbm����5��A6�6Tz�L�9���д�K�4[]赐'���r�5�1�3j�R5��K�f\�5H��4ld\�Qљ�$�������w�z����6PQ?5�G���y'�>�9�i�5>IO5d b5��5��3 ��3�4�ŵ��n40]��$h�� �-1�]�4��6� �O��5TM,5F�64@^6��506��7�d�5���5�0_60u�0��#`6�a6�Y��D�5(��4�p5����Kt4浢�	3��5�;�@C�5F�6��5�`E�>Z�5�5P	X4aȵ�[R5l�L5	�<6�ѵ�Ӵ�<5���5�T��йF5�ۜ����P��5���3RM�5����A6�4�4h���
�5����V5��35 < 2PQ���_�3���4�[5`т�ࢠ5f�260Z+�B7ӵ������hI�8��4(��pM��,�350�5 �^6`�&�����)�5._a��� �Z�ʵ��#5���5$�⵴lh4,߄�@� ��85�k�g�6������
6����l��5d�S�9�P���5и�� #4&Ȟ5�1�r6��z�5��ε�$�4�z�5��X6�a4���5�p�_�����7���I5��s���-{�U�v�L{B�^+� b44� 6��V6�ƶ<E�5��Ķ�cs6u�2�탆�i��5�6���5�17�hx[6��6�kŵЮ6���5��/Ե��ϴՊ_����	K�	���H�����6��3��ҵZA5��� ���4HF5�A��P�6"������69t�!𣶸��6�	4�6�V6,6ܕ���6�� ����6)���e���G�5@����26O[�5���JO�(E8��b�63�#6n-���;�6����[ �}p�6��J��A�5`;ʳ5�66U�7�r%����̶h��5�F6�d��T�2�m�Hg���5L=6S$T6��5Ķ4}�6ހ5x��Y*��y	6��ٳ�ꍶ<�06p����m�5�i5����|�d��3B�	6��n6�m��T5�E�5�2�6�����i6N6�^V�ܞ�5��նЁ��[�6��$��EU��v�5����)z�?G	6¼���2��ڴDQ��h'��aD�ߒ5�_6Tm��gB�FH�4�e�5�R^���$���P4첓6�^�6��5�(�`@�3 `q2ӓk�6�-7�:-�Pca�<6�����(�5xل�8��6!C�6w<�������3�f�6�`�W����g�5��6b'�6��5;�6m�Y��4d6!���u��B*&6���� �W�p+�5�����Ơ6�K��{?:6��6C�6w�5��紶�ķ6 �Q��Z6@,׵�a�4˳p5��v6$���5.�j;U5�5�.(�{�6�SS�.C5�C4n���0�4��P�~=t6�Y\��e���_�Hu ����5��6�Ov��/�5�.6?1�6��S6q�ĵH�4��.�FNi6��U����6���5�Ķ���5�ɵ:b5��S6��&6�(ų�l�6��ɵ�r"44뙶;�������8��V�6�&�5B���A�u6�F4 Y{5�I6��̵�q���5���4�J5�ځ5�25R��x���<5�_��x���LL�5�6.�76E�9�.#����������}���'@�X>ҵA!���5O6z5{V�e�	6�!Ķ ���E��2�5��j5������A���5H;�4�޵�{�
�0�9�3��∵��h����.5H�6���ȼ��H��4ZN����@I�3�j��Զ�˄�|౴�@��S�6���xK+6�!ֵhju�U�K6�7G6�{�5��`5~�<���ֶڧ�58:4�5D�6�+�,��hj�4�����c6��5b��6�2���j���L�b�6� 5��;�B6�Q6�%h�]J�5>ݘ���6Z�5��5(��6���5��u�NB�쵉6�ựx\�x�t��j���Ӟ5�W�8Cp�}s�5� 6κs5��8R_5٢��na�޹,6�M�5DQd������5�� 60#���̵�/�4��6�����H>4��[5L	�5b(�6=a�������5,X�N��4@Q8���n6B�#�`��4��4ԖG�.Gd6P*3��U�X�����3�1|�5��	4ӽ���,�!�5[6͡� ��0H���C�50l6�$b�l��u��dKf5��j5pl7��i�3mG<��ۣ����6�R�5�y(6�%�5�$�6\��� �16:Զ5��e��d6��4PB�����5ī6�A#��D�5�6_�'6!Cj5��S6"�?6�S�U��;�5�5�M5�	����D��%�5vc5�d�%,����Z6>�-6� ��k��d�96��6B<�|�մ ����6�6h�6����y�4�쵍���`�_3��6�㻶d�^4�uC6�_�4H��/"�6��C3w�67�6ְa��Ck5? 6n�5^��p�"�`��3&�5���4�n�5���8퉵����C����b��k>6�>��;6�^�5�j���6���53M��n�G�v�50�4����L�3�O)�C�µ>�g�_�86�na��j5j�6�U�6�\�6䕍���6���5�s�5&n�{�6���6�U�5��6��
5�%;��17˟�)O���w�6���6PH��k�r��17�)�BB��'{��n�6��u6��8�Ф� �$�:��6xP�6�Y���6p�>��5-ݶ��5l�6b�6@~w���6wM��X����6��y� �A5��5�ľ�H�h����3܈5W������%�5/H�6W�6@��
h��^�5j֟6�9���ؔ���������7N��������h77l76J�7�j7���!6@<峊Rȵ�U�6/p�����TR7���6'�7��a5��6������64�7�GͶ*�6n��6Y�蘔6&�&7wҶ�^7��f��{=7�坶�P6�˓��Ƕ��7�d춆�7o�f���"���<7 h�6)!�4�����4��~6�
�6�/6���K/�ʴp ���7�R���6𰲶V�6���6��6�U��<��T��6����N�6��5�%���a{��&��vo�{|�&[66!MK6��6�$�52׶�(�7�5�6J�����5�[Ķ��6���6[Dl�k�%X��v%5kj�}�6.뺶�G�����rT�6?(����7oV����6�@�6zơ6qD6R$6���6������6]Nx�2��6Q�%����x�z��7q�U���66�6-̶P��7��6o�37�pB�R5�����X��5��?��W�
�7�Q(6��7X{w6�,��}ow6�6&ڥ6���7%{�H�6���6  ~.�+�6��W�%�N�`6�9ɶ��f6z�/�ص6�� 6rv��i�6Ć���37�L�6����mڵؗ괈�ߵX�m��؃6@��h�4n8�68c����66f��Jc޵��K7H�Ķ ��4.t��P��<��5V�����6S,7�`���)e6���6��6'��6ʨI7��-6cAp6��5�:���6���.��5���L:���}J���붿��'�6�R7��5T&X6�~�6F���z�l�I��5�.�E�5�#նn���0�7&�5�,7*�ɶ�6ִ+7o�67-�����Ӷ"����$7&27l~1������T6t�.6x/w5P	d5�h	�Y�n6��>�ߒM�sn��mk���� ��5�3�E냵��{�lUB6���� �1���rB$��%d6N��5��Ƕ^r��n6�7<oT�b��5�6B�Q�����64�A�~���a������6�4k626t���7���6wA�覒��7��f5ڦ�5�BH�u �6�O̶��*5�U���9�6Ϲ�6�5���6�d}6,�"�ʶ�q�6
�B���'��S������3�I7�C��FU6R$b��=��GN{�u!޶�X{��<\4�hS�������6R)�UV�5�Pp5�o��H������q�6�;��ax+6��r6?4�6�[6�ބ7��6V��(8�6�:6�]�6�Vc�u26�1�0<�H���B��!�[�H6�\	�޿���.���凶'�㶼�/�_6 �G6Uo���?45������b�����6 o�����6����)B��2�6Z|��2��m�5���6�!6��6.O���c��wHe6��X^����{�tP��N�0��(ϴ1�79v"796�!3���%���7��0�ಮ�p)S7�')�kc)����6%97�+���Ǧ���7P����5�<v�����3�s(�e	����߶�0Q��P������>16l�b7��d��4b��]��wj¶cZ춓G����6n�\6g���?5|���6���mT�6��6�+�6�]u���:�q�6�Ȃ�^��H5��9����ʍ(6���ѥ-���4n�7J	�6`6���6�8�����۬!7"��50�SF��� �62PԶyW-�>'\6�_�j�F�-��HD@�dr�Щöp4�j����Z��ԏ�́���68Դ������ �>_%6�ޝ5pL����s����5Q�5,6�NqP6v�5Y6����&΋�	�6x	�64�6(�<7�An���5%\H��r�5o]�5��$�.�e6 ����	_4:L۵!������N�6�w�5�#p�$��6��R4�T��-6�����<��p��;�6���5F�15�x0��/7�7�12��4xS�4�n�5$�6"懶4�7�p��bp�]�7 3c4�x�q��6
�7�DOA������5t�i� Nu7v*�6�O���y�����糒��6��tN�5��J28���5��6�a�5����zҶ�8����N.�6@���y�5$+�5� F�������3�� ߄�͘�5��i6�Pr���5�^�5��˵�d�Θ��޸6d]�vZ"��|�6N͵�,��5*���/b4�[ն�k�x'ʶx ��Т6�@=��V��\�E7\�g6\�-6Ff�'�6����F�}���t6'�>�.W�5N
���g.�'�[6�C�6'Y�6�)���v�D#г.t�`�m�V5\�T��7\6�ű6� �5?�Ѷ�{�$,{5���6P��7��K�������@��N|����-����L����6�Q��Ї
725�lb�J�56���>�5x�6$|�!]�6�춌�7�-5�O76*�)�[�7"��>&�6A�6q�50M7���AT��J��5x�ε/�����	�['6�t�5�Ǫ��6�6��I���6�;C��϶d��6��6�<7V��68�`�xU7�&�6�m76�6���5iW����߶�"�!!�5f>7%��62��6Kt37�N�6��5�mA7��������������5���4ɪ&6�9�.���H7Ϡ�6��p��_��Wu6=�v�i�D6��6��7��x�=3��D�LѠ�~����B�6HT!����6��6X_�5�s0�36��36ъ6��εe0�5}�0�1�6��6O|V�Sx�57Y��T�6~"r���~6��=6�#06/� 60=���� �F��ż��FV4�e\��n����57y���Q4T�ìd��	^6�v���6N�ɶd�O�K�6?GH�(�6L�|5 G��c¶~l�6ޅ�mͅ������5&2|�G�5�ʿ�5��7��>7Y¶�"6����&ܴ��6A�t���+�6F66K��5�g�5��e6x.�6ܡ6�uT}74�6��e⬵ޒ51[6�e16ɽ�6�g���D��v.6�pY��2
��b�5�O5��	�H�l�Цo6�0�]�&ɔ�o�d��3�64[6�5ew�6��6w_����4x[Ķ6������3�6Dh����L4�Э6|<��ֹ�6*'����,7Rv䵋t7�s��ݞ���^6Ը/6��6� 6}KĶ#�=6�Q�6p�|���3��4��H�5V�5�c��3i6Ǜ�6O�6��|�{O6�iԶ��)6Dk��ԋ6nl36�:Ŵ�q6��ɶ`Ѳ3~w7~�.�ᙶ�@Ӷu���ބ6S��5��V����6 �M57�W�5!�c�=g�5�N�6��e6*q<���$�"N���6Hu�5��5}w�54�6�Y�6���,���7lp��8|6:Z���P"��?L6�s������$�6mGL���ٵ=5�5r�:�]G�6�,�6!�����t��S��60x6����ʵ��5�j�^�R61*A6��7ӗ6/�r6|,y6)k_��Ё��6�D��5|"�5��5A�a6D��6����X���ж��4%�!�V�Ѷ���`����4F��6��>�*T�6F�/6/�{�G2�tM����?���׵�&G7n����6��O7�7z���VBT6����dR��:6�϶��6����5��5�Ё����R�L]W7M�5��&6?�0�@�c6鮶���6�65���4����Z�l6@�[����,���(���O����\5��ƶ<#N��^
6!ܚ��|67�����6s�26p1!���6-��6�.��Di6��6�,�5QH#6Ţ�5�5��E�74�ǴT�36�`��p�涂��5e{��c㶿U5*y�5}g7p�6�Ǩ6��6 R�6ߢ�62��6�O��D/�6���5�EK����HV/4j^��\~��`�5<-�6�7�5��4�})��06���������\���4~��6�A�ܸY�.$˵)�36
ӭ6���5���e�&������S5�ԴA�۶�1��(��6jO��?궩h�5��6*m�6<��{Nm6���ʸ�*;6�16�Fi5�=�6�w�2`��Q��x6����R�5��6�d?6 Y;6���_�ٵ����W�5^���h�3��L�4�ƅ�����P���d;�5{�5�	6E�6���zɑ5@��3�?`�]�x6�J�6HR���>�_J
�.�6���69a�����s�5��5f߶��H���o6�œ����{
��{�_j���ݏ�6��Զ"�&5�=7�=�6}4�����7�_��̣��D6��6s�?��< ������ٵ�)��؏���5�t���Wܵ���3��)6���������L���e��6X36�u�5F#���"߶�WE6#s)�&�6��6T[R��ڼ5 Q0�k6�R�(G����54;5�ݬ6v����(���i�Z-���p6@Z�5hѥ4�	b6�q洼�J
�6�4�5���6$�V���ضL�鵤P���/
7����N{�}����<�6����3t
6�q�6�*��026)S�6�v��t�ݵX:O�����������W�7����Y�E6�6 ��>���m��67ЕR�lY/�7ڌ5Ǟ���M7_�[6��2�6�&6$��5@KH����	3���v5�0j��#�6���5q<H�~�̶C_�(�)��{��rP6j;6�
��c6B�նH��t%���� ~�j!����Q��/R5�d6���N�5^VV5�*[6�X7��v4	;|6��P5"�64k�45�"Ե�@�4�-U��|6�����6�7(6�	�6l�6g��5of5TM�@FX6��Y�rY�
$��X]�=��L��6��6B}A�?��6��6���5�z6s+�6��X�u=�6	ߌ6�"S��j4P�'�^^�j7`���ɠa6x`���5��5|�S���_�n3�T�6�[��V6Et56l76�Z�����ӊ68<��^fX6.����ե5��&��56\)����G��\��g66k�ѵ��<5��96P���O5,n5���5�4���5�5֊�6�������@�����u�>W����5�ص%��`l�5�;���du��O5���4�o.4�[�_��5Zp5��/�v[���U���5p��3sYt6��O��y��5�u���O���j�II�����#�\��z6������6������6�L6t:Ͷ񍂶�0�6�3ô�494�m5�ό�(U�4]{ٵ?�5>q�6z٘���5�2�+�[6��6���6x!�5�Hp���5s�5��f�4eҵXȴ��S�J�W6jec5" y�j� 5�KH3���6�V6a�p����5����f�6.�2�V%&�v��շ�5����h^��MM��z�6���4>�\�tR��5�A�6lBy��9��h�6��&��A@���4���"�x�O޺6^ͅ6��D�}⒵�b�5���~�?6�8�6�f�j-�6�-�3�Ķ�;6��&���6x�?6����4�)5�Un5x��6tEִ���6�G���y6��6Q��5>�(5T�f5������6�C 5x6��5=��6S��k���'��5卆���6�vN\4l�:�� ٶk�5)>��l��5�ĳ6�7�32&7
Vx��q+��J4�à�D�/����5�#5��-�;��6��6,�6!�6��� �D���H5�y"�\6�쏵��۶߾�6�[���5ۚ�5bJ6r���l~�\X�����6L���:56������@��t��U��6�J6Xz�����6�'��x��6�h���wѶӽ�6ر�>�q�5�5�J;6N����5E��6\N�}�6��!5�L���6�����퉶㷵�؁�����^)��#!��� �5�56��46᜵�{ݵ���h~H6�]�6�A3�A�H5 ֎3��o�A�V�݃ ��Y5DL�6���6^m��bw��%�6r鯵�c�6�H�6�&� @6ś���t��&,\7�:����@6 m�5\w[6N_6�F���]�6���5���5���w���6Y k�<j�6̴55�6MYN�r����ؾ6(�Ǵ�5V��x���W:��X�67��6�h4��w6Y�q��f�5��
5��6�=�P���ݶ@YG�ol�6�>�5F���q�ö�"����6���� �c4��6��5�Y3��Q����$6�&f��ʢ6�0�5k��|��6M66\�����'�5�����ж���6��O���NJ������>���0����V���Գ�5\�"���t��b5�rU��렶���4d�������
6�gP6�l�6hW(5���5.o5���6�6Wm-5Ԋ;��r�>C\�l����H�ᵚ�'�|J6��/6ψ�5z1���D�6�r�9�f���a8(���6!�ȶ���5W�6{�5��U�Pd�4��o��"�6��p58r�6�x�����5*��6�U#���ƶ���x�4{6 u4&���C�6U��5�85��k��d26����x�5%��6hk!�Ddp5"H̶O36"[¶̈ٴ�>h���g6Q�뵆8�5�7� �!���h����P�Ni�B��5r�$5��5���6�!M��t��NĪ�( �eO����5�е�[)��=ȵ�_�5-64�>�c�l����|����͵�tW���5��L�5@DI6�ɞ6�
 �PƐ4�������g�5�Z��dR�t�D���e�4>A�6:L��`�Bż��v6t܈4q�X6Ơö��5������508�5xgR�\�t�^�j6�<���)��j�!��6�5�B��3�:��_s6]��ЫW5hmb�U��H��6�$�5�35��Ƶ��Y�N{<6�d�E�6��<�6t�7%��fq�6�M���O�6h���@/� �d5�mĵu�(��^�6�~T��*$m�NA��7V�� ��n,Q�����r�5H� �4M¶����$}6Ҷ٫��3�5��6�����!���(+�6O��5�b������ �6��s�^�����R�)6�H��x�(��6\�c5�2�6h���}������H�6b؏���7���7�\ض�;���&�6t�7�\ڶԜ#������ 6 E3���5�e6�7�`@6v7�:�5:p����5;�}6	��Ţ���6���6"���F6<���l�ٶ8�6��7nk ��s5j3�@ݾ�Z6�64�����"7��A�d.��J�6r�����{6�џ�Y�ȵ�b_6������6��6t���:6������'��Q����>�6P���`��6��6L�6�P��J71���e�6 ����5>,`6E��T77�r�6XIj� ���v�6�A6(W`6�]���';��-G6�˶��_U��,�6zH�6$o�6�-�5Vyɶp.���U�5D�ȴH�4�C�6fN���ٵxKǴ���5%�6P/�&\� ;5D�@��a�6Y�|���Y�-�g���6%\
�	1��p�Ͷ�ߐ6��6N��5D\µx�D�0`44zO7Ҷ)5L��6�n�6�T5��9�e�ȵ*�	7<��6�[7i��	>�0a6�� �nc�5��"6@��4���6퐝6Z���(g)7o�E�ƞ^6ƿѴ����$�E���Q5�A�� ד4Η���%/5�?06���Bf���6\��P�S�'��6 �4��x�64�6(�.6�,5 ��2�?��Hr6�E6rc��R�i����5,�4�_T��u75��6�s��p�7���1��z=67�5�����6%Ђ5�۵�[5*k
����3�h�ȇ+��l6Iy�ἵJ��O0��1)���p4Ϯ�5xn���8�4nif���s�������#��D�D�ԫ�}�25��9�������5�~6�x2&�96���6<(����_����tŤ5��5��������E
6r�6�?6$�Ҵ}���m�ܥ�q�7�4�5�F������ě�5=m��c��5�*g6��*�@.436��h�9��4^46�%�5B����p߻��+�4�`+60�37����u5�յ8�p�16|	���D%6 �B4����:cg�~�1��96��58�����5�/6� 4Ħ��"B��c�6��;����5F��5t75M��4mݽ���,63�9��D��i��GA��@����5��5��6h-�"�����S4�m�=�!5�C�8�@6�/u6D��5TJ%��53�6lP�>&5��V6�:�C��vgr�<Q�5�� �ǞK6h��������}��M���*�6��5_�5.������0���dP	5X"�"���VQ˶�b#5NX`6���V���M�67W6�h�6��쳸�40>���Z6h<��6^���@u������e_�����O��/�4�VV5��5P�#5�#]����6��i5����݂6���ʷ���f'��[�<l6;$6YML�Y�5�eU4�.�5�6�%�����I4�Ct��J6��
���6�i	5:5h�@����6�9O�4�c�+`�Y��?�]��� ����d�6��/�66�6�&��F$;��/� �뵈9.��`76�i��`F����6p6�Cq���P69���0��5�W���e��pĄ�Ғ��$6��ֵx��5$�����N�Dõ��O5��35�浄we�j���aᆵ��4��$6����zrC6}�4ŋ��H~�4���3�5� ��6�J����K6�H?�֔d�[Os��T���S�O��m|���w������#�r�>�$�o5hD�5X �P� ���5��#�v�� �L�68�B�zn0�H����
�P��5�F6�ؤ5dik�R�I��g�5H�����j�}�۵,���������5D�3�NYյ�����3�I����6������V�.V�(�q4�m�5j�7�~lB�|���}?�5վ5���5��4��	�46��6��P6���$*�4�9s��~6Ά6��96gB���/�6�s�5�55�\��R��5���5-�	6X�u6�>2�J�ŵ\a��6��D5X�4��,�^�=5�� �(�P6ߛ축
D6���5�R56��B6�|52^^5�pL6�����w��J6�T7��26J�P��͟��y6T-z����4	�x�`ɜ4<�k�}�6��v5�p�5�,6�^��׵�x�5+m���}��k6��#����]�.�\P5r�3��B6+f������m�~%��(B�҉<�,��4��3�y5G��5�(���v6&�r�^(��H�:5ܵ�4�Y6]8�5������.����5�|6�7+6��6��6B뵀�}���Q��4�53 '�C�5���3,�26SZ16�G�5��]5 2�� �K1�Ze�D ���D� �,40�����4*\�6�u�5�C`4K�i6�IF5a?�5�{)5�\�5�^�tPz6 ��1[&G���6�3�3FE<6�b��&�4;�+6������|l��5>�^6��6SW�5�t(��uǶ��45j�6��b��Q��(G3�)�6���66�P�F���p��4�:0��5Z�M� �U;���wK��m�0�8i�4t566����e%�z�	����6�̗�k��5�|A�V���nN4�0�3��ȵ�^t��y�4�����9I5�,����5��M5�D7��6���5�o���>6P��5���4��4�8�4�ﯵt��d{���.�ad�� 54�ԝ���5hz۴�V7�wK4\�H��4�┵�[6�M۶⯄��7��V�������r(Ѷ�Q5����6X���vD6��6����<����=1h�h��5�,36��9��k���Y��n����?4W�x6Z�͵������w6�}�;4<�`�2���55	Q�>�K6�!����5h� 6�0µ��5����nA�5i��6�>6���5��F�����x-µ�~�5��56[����6L���� ���O�5���6��4P�7�s6d)��z50��"�յ(q����J�(��ܚ<6 ��3�ߦ6p�~6�o�6�ۚ6�}�����@o��uJ�57`E�������(�H.�5�3
7�m�~�6r�G����\�˶8�5񌒶��5!6�|k6TT�5Tg���+�5�${4���6��y5�᪶Dy5������?���^��6�Ƃ�����5)����:H6 )G�̙�|k;�7�w6ׯ9�hh�5�j�6��6H�6��嵠k���f6��16��M4�-�*N��CP�6��T6�~��D6�o⵿/�6�k��pQ���K���-����6`��5�߳�*�6�u��������5�@�����d�5�w���[7C�@rZ5�Ƕ�iV�BWR6���2�t�5�B!�p 06@[J6�D%5�]v��*z5�, 6@Y�5�9������B@�p"#�4���������4K�.6ڨn4m�K���u6O�L6pm,5l�J��i 6n�?�P��5�5(�B�!�W������x��Fİ�^r6��5�jŶ� �P�@5������6��'��}A6&�46�N��nϼ6<�C��[#6`�����w5���@��3���o*����5e�<����5.�������Z�Ƶ|<����D�6�4*<�5\�6�P�5=}6�g46�6lH��w96�o6�N68� 6���6z�N�6����K6d�j6�|a6�ZK�,?_5qg� ��6���j��5�O7Ť5���6
6�P4`F4�㭴��6.N1�����8�d6�I��lV�5H/��)�5����'9��\�s�6���4�5��s6�]�\G�����O�6CCX5tby�sԵv_��6寧�e�X5���4�e6��g6[��5Wɟ5v���[*����5ށ �Z�X ���4kܡ5zeֵ%疵�G-��Gn�L�&��]�{�;�\�160��5K\�5���2���5�6�\��>�v{�5�R~��v6��66��5Ȣ5G�C���O5P�v�i-�5�I��E���Tί4Z�?�ص�8 6b�p����5 �6RG6$�j4"C)���K�
0j5J�j��c����3�w5�Tٵ6��7�P6�;'5��|6�u�3x���G����0����Ⱥ���V6MU%6�p{5`��5;�C6#� 6d�h32"�4�z�(�4�gF�z{P6�)9��P�l�S6؁ � �����s���26ԟ��p�5g*o6������-6𝺵r��|
5�h�5�Պ�]����m4�_s5�X�4q�6���>�ɴz�_6�E�55*����y�3��5�K��S��+�6���5�ﾵ޼<�)y�5��	5x����HB�ڹa��0���l�p��3@��18D(� µpo�3�N�����`~���5�%�>��5�����ᨵ��?�z���hK��Ƹ�8p65;����<_Z�����ĵ�f8���r�B!�*�h�Hj6��\�c��5,�d���	�  �j7���X�4���6�w ���=5����)65�� ���5`�g�<a}56�W�)a���S46|M7Z54�ƵBK�5���5Rʦ5`�5�n5��޴����4�d6�iB6�����s5�\p�w�)�0��nMܴr��4�H�5��565��51%N5�_/61�k�w!��A�д,���5xe!656�Ѓ�$���$k6N�26̚ ��P6�I˴ ����v{5M��6(�A�$�q5œ6��5�@6�����(5嵧��/#�@��<^�hf56H���� �LEX� ����[6�6c,�5d"`5�6]�'��ֵ�{4@�ٵ�-�� 4���55v��5�ғ5p���������6@0�4@��4�B�5B����W��Y�QV6.��6�VJ�b~�5(#w6�7�6����Z���n6,������]6�6ؐ5`�	�C����s���6�	7@{��"��5��P5�n���I����\6�1ٲp��4�6��%��u궫�,� �T��F�6 0�� ��0-I����6D��@ �50�6��V6x�ߵ)��5`伴^��nFw6��S����6�8�5���6�d�������O�5@p6�f�5�85�S�5#y�c����֊4��6�^6�K6 �g� �Q����5'����� 55Ǧ����6$ж{4\����`�5��<����6@7e4�K�5�QH�;�5�-�'ǐ��DT5K�6��7�`�G��+���W����'� �O4"��@6��~�f�õ ��3
3O��@�Uʱ�}~�k&56Zx���7��������"5)�V�O6 Wᴬ��5��5�j�5�OJ5�x:6��(66��\�`��4�	ԶZ�6Rvu6��3&W���x�5�6�`��h5Za�6׃����'�|م�֙�w��{58�� N$5��s6,2�*ܣ5p�7�F�5�����P�5�n���M6�lQ�Ծɵ:������6!EB6����j�5�֒6�E��"b:6%�6�d1�b%�6{��5�060����G� !�@g�6������
V���P���O6��j�@�Ҵ(� �H5�-!�&�;6 r(4��)�h���n
}�`:6Ɛ�5$�$6��+��5Ӵ.������3Dq�3q�/�D	6
b6
9O��2ҵ�����5�2��U55��j6cG6Dh���6�G�"�%5����Sr��HƵi�%���5J�"5����w�6���Ci�`�6~N��K�e6���m	�5�6Z�5"0z������2�31�H�y��r���E�B;�2�[��@�6$a�,�G��q7��+µ"�p�����Ը���l�W�^6 e��rc��p��3��K�o�7��޶4����n�6 .6�`M6ڛ����#6E�����U�m�H�����յ�3�5�e{5����@�5S�6��b�](�@��Ѓ��^��6�6@�3�M����6;�ߵ*!6
�޵ �z�����|�����6�l�6��ݶPg_�?_o�FE6&ʜ�4D�5�_�1�7�-���7�4Yď5%Q6P��6Hg6���6P���mn%��%5�5�O6������_�	�Pץ5J�.6=$�E�x6���4�L���A"6H��-���4�5n�7��5����46�!4����H;��6F�P� C��d�l�5�W�Yf�6��t6���Z�Եɀ�37��40��60�5�U!66Xn����ƶ����@.��b5�s�5�D6t�϶���5�H6�}�5Q��5'�;6@k�3$;���%��Nf�$s��?��6���6���? �6ԛܵ��3����6���5����@�s4��@5Ȕ:6��6^�`� {�4��G�:�!6q'����06o67Tb6���4H`�50ݷ��g6��7�0��"N�4�641�
�68�5226?T�6��6���6��J5���ӯ�(��4�qZ6�T5���g6�����6v+5��K��~�6�B�5��)�C6��еxY6L0.��S(3��B6H1*���z5���YA6/��6����rF�5F^�1 �� �b6|�V��Ve6�$�6��k����i�g5�D�3��4ӗ�6`�����4H�
6jȩ5&ڵ���4R��[5�I��� 6bڶ�\�A6�7�@��4�p
6�v���,6	�j�P�i6�ֵ��'6=�e��"� ��4�Q6�2�6�ϵ>�ҵ0��=�A�`6�
�X\`��z�6�56�C�4�+�5&)4�;1�4��6�Ӂ6VJV5B��6-6��<���f5?e�5&%�58=�5Xk�5[�W�R��L�S��JL6�q	6A��F���7�r�58]�Ru�����6�r����ض(M�6��6�"��x�ֵo��\6�^f�.V����5��v6�3{62!^6PC�6���اu5P�4^m��?5�؝�����b�m\��a��P��4;}4p9�6%�5�xL6�v�5�c���J�|Kt6%� 6���5F6�/s�k	6�6�
������@6���5�]�1����4�p�Ј��j�4�Q��+$6��装�H���!�5-ģ�<`���66���fa�/����Ee����d6����$�S���6,�|�5��6:���!��j��4�݊����5&�m�x+u�"d�5���4��h�x�ö>d+��ա58B�6w�6{I��B�:�VN�6��ʴ��������w��XB��R6�Du��m��D��C6�	6H��S�27V;�����5��D5����Ln�m=E6����.O5,"N���5鈵6�Y�6���5�I��Ꭵ�Ν�� U�2{ �6��Ķ���+��6�ۊ5R�6H�A�jN=6^Я5|��6��2���s���47�n���ôD�%5[Tx6,w,�����yY��>�[�,�p�Я�4�����$�5�5D�60�ٴ2��5�0Ѷ󈡵ȍK6�搵\�����6մ���35��5�=j63��p'+��P�8	�4��"_6<}6��h5k�+��<54�@��씶X�6�45�z�5�V5D����ZN�ꍶ�86�Q6�(�6��� ;3�%.5�6�6i�36��6C�`�8�5��6�I��ӡ5`0��I���dJ��?�!�g�"̠5�5,�4��6"�^� (4Y���stF�0T��݅�Lu� �j6@Z����501%5d�6�0r6�Lr�����5����d�h��c޵�����͓���3�G)��&�4t 60މ��L�5͟4b�5 R 4بϵ�r����:���R5�Iu���.��3�5�����T7�� ��#�J�6�������TgQ5�5�ʅ6�k8��<6F�e��/�$/6n M�.�6�m�6r��6xP�"���6��	6��d5�������5D�m��qq���5�ﰳR�,�|F6��
�
A7X������6����Z6��6hP���:J��Pg��HM6_�	5Np����!6"��y�u6��6bt��N�v4�P_����4��6�{�>�i�p%�6N�5i#��Dȶ�
@5���5"4vA{��|жhG�4�.����R��g���f66�i6����{׵���5-a�6���4Xcx�SLK��������6ͨ�6���}�_�u��Pδ戟6�����76:<�7��6؃�6X��54~�6PH�,o�5o96`���Ͽ�֘�6�P�6�r6n��5:H3�h=��]~�6�.���4u Q6d�6�`|4t�@5��6P��/습Ų;�~�6�u6����"D��N#����5��P6T'�5�5�ǉ6��S5OC2�(�;6�/B�|�>5���5[��5F���]�C�61x)6dЅ��ׁ���5}3Y6	U�#��Vކ6Y���6Ig6,1-5f恶 t2��E6��A6v헶�?M6�(��u��6���nN�5a 6�]�6�EN��=f��&50���q����23ִҵ������5d$=6e����Ŋ5�_R�񺞶�TN6VN�� 3&����4�h��cd5�q�6� A5\p�5j�6�4�H�3�?6.w�5�e´�[�O97��h5�|7Z�J6�qc6�d���|5���6�N�6���6�a��ƌ4`������Z?�6�y�`+��p�7�>�6���5�`7 ���!u����9��~;�4�v���x5�5������A6�δ�]��4���|�ŵ2p�����36�6��
��!�6�T�<h6,'6�R۴�F1�`]F��>$6���5���5�.�5 U���մ^�5~���`���6�I5�>-4P�+4�Ŋ��'�5���3��34xˠ4�$�4�����!�4��γ��_5e����6�=�h�5` �
W5�(�5��S����5�I��%�5�](5�J ��Q/���S�����L5Ъ5�� ��b�5�5 �"�6���O��o��n'ص�m�5"�M�%�5f:u�� :�y`��Pƣ3xC��N6���3�Y�`̼�p�	�N�6�"6��ʵ��õ0��P=����O5�  6!E�������4zX;�m�5��H��b6��5��.4ھv5�r?��826u��5y�5�r ���4�Դɞ�4;߫�T�w6�?�5lb6;+���j�5xpF5�)��L���u����5���5�ʵ�N��04����<I���?`6!�6J�5z��4N��44$h4?6_y�5P^%�*�5���4����k5�e�5M�K6� 85���4xT�44J^4���5�?%�+���^�5��5�~#��#5P>�5�LL�h>Z5@�n�|��5"7��HT6�(6�bc5�6F,-�d��5ƶ6
�N�2�,5�^^�Sߵ��洯�#�S@�;�4����-��L�R�5�*b5<�%������6P}��!��W��v 06�d{��g�5F��5`���v6<-�4�$�5�B�0��3LPʵ�z�5X�5��36x�5�H36d��H�/���5?����,6�ل��~ߵ�C56��P������Ե@U3�lC�B���:��:N���!U��]2���&�W�̳��6|qܴ�S6.�ʹ�Q�5�@ڴ��͵�^�545���a=62��5��95j}<�*���5>�t��4O�66鳟�8�-�l���_�5�=��UB��2���q?6`�4y�
�3z!�5@��2�+;����54�65��ϵ��
{̴i�/6�(�5ȸ�3�*5���@5,1b���|�8���@*е��)�H��4���� �O3��5+��2�I6I|� �5���I�o6�A7�~����U�B���$6�͑5j����Y�6�><�
�Q��w�5VU�6�� 6��ѵlG�5�$�6�N��D��6T/6�^Ĵ��~6��!4���w^�����6�������w;6���5�]��)��wm6:G���7Wӵ)d16=��5qЄ�mꖶ�ǁ6 l�4�6�8���-6f��6���4��������j4����|�5�?6Nf̵�P�<��sD6��k�1��6�T2�RsJ6�&ĵ�6@6�5�A����v�峅5x8�6���4vY������5%55`"6�u��f��4nEɵ��6��5nNٵ��%�Z�j�`o�3�����;5@n23�}�0A�� �����L�6X��뼝�n��6 �x�����!-6g9l���Ͷ�����O��T��
�f߶����#Ķ�\�O��x���s��_� ���24A�̵L��4~ɶa�&6h:e6��R���6��5��_����LN��T��5��3.4r�HA�5�o�5�>س���Rl���7�9�52�X5�pW�@^�2?&����(���U�-c�5q=y�r6�/T5�n���F�� �1e�6 �6���5Jڜ6.W����5a�6�M���#���=4hI��6fzR�]V�5v�?�v��4pR���UC6��!6t������������a6-&��ʛ6��޵S�H6K��5���5���v�k#6��3��{6�6����}��H�u�,⮶�_6��ζ<�O�0�$��n��i8��ш]6a4�5��&4.v}��K��/�V6(�Z�|�63*�t�K���ض�[�5 ���Y2�5|�4Tװ�<և����5`����6d�8�����������ضlE������ǡ���\�6 �6>�6�4ȶK��56�����5<	68u0��(�K�Q���a6��5�X� /��s$�FFǵ>cG�Uwa��Q������u5%���х�F4�|�p��2�y���&���"=6 RC3 sE����5$��6D�(�Ί��v86�?A�0,��2_�5$���7�5���s02�U����5�2���#o�VL7E���`�3M����6���6�=� 卑�:궿�;7:7�E���@,���77��T5�jp5 8��K�ѵ�i�5�~��K^d6���5��69島��s6��^�qZ5��)7S4i��x#6c��6����`�-5Ѹ^� I4�[s�37�B���G�$7εEǍ6�6��衝����5��7>���5��R7��6P��4䵲�(����_6���#�g6^�5�d?6F�6�H	�|
�c�A6���5��6Ә�>%%6�r7x���l���
Iy�1 |��2�6l�7 �6 ��60�L��'"69�� �0�A�r���^��a����I=6������v5�3�5��6Rඒ��0��=W��)6F!�6����E>54��5�:�� ǵ��N���*5���/ �ʻE6�S�3![����.6��5X�3����5O��m�6ӵ��󏒶�F5�	�J47�T�4`-�3�;�6蝙�û~�,��6�)v�16Z����`ئ6|���A5���{<-�r�Q60�4p��66%"���h��6V6������`���4a�6`��3��^������-6������6�I��|��r6��ж�W��bo6�����$6�f����
7��R� �&3�w6ȥ�5�c6y?L6���6d����	X6��6g`6j�?�]k��7g�6�}�z՛�ޛ�����5�o�6�抶����=6NӀ�뤓�*F76bj��KI"6xd¶aU6l�3�3_7�,6),5ھ�6��6T\�D�6�䁶����~���润���e-6`6���ЊU4��n��v6���5j*6̅�5nP6tzZ6=�����h4�7N�K^�D�5E��י6���6hK�4�V7�ȇ6�8�6��6=&6�C6`�/�J��5^Rq6�	�4���ޝ5�76Z��� ��(�ݴ�{I���(6 a�q�{5t������F �$��X�A�3��ƶH<d6d	��L)`6p}��J6��[6��^6Em����4�/Z6h�d� Ӿ3`A4+{����h�pʳ�%�)������b�b��5H��� �������7�6�Σ��oz�2Ia5ڋ5����z�j5���p:�#��6��ܳ��_5ʤ��(�5/�_�d�����7�n05J掴�6��tj689�4��5�iV6\g���z5>��)��gf5��76�����B��qʆ�#е��r����4f_�(�6����P0�5��|�n��6���6_L�5k,6���T�5�ǝ�����*G6>6���R����5�����6�dF��
7[`L6�c6�Q۵�̔�Z�,5J���7NR6��G�̓[�p�3zs�6�6������A$���Cf�������e�5��6d����c�5� ��j�$6Q�5rO�6����`����6�;���w�5C'7�,赬rҶ��.�8��5��!����5o9P6�86(�;�&�61@ŵH�Ѷ��4��6Iˌ��p޵U���d�0��5&66��5��5�!6ʁ̵���50��Nd����6D*R�^k�5T��^ꔵrz���浽�3��Qw��5@3����(�|U<�8	6$-�6�,���6�Ե$�ȝK5��/��t 6�}�ܕ��k�4��6�+�6�l�@f�4�6�, �邑5M��5�����'����rq���C5������g���4��>5Ȑ��󉚶�?��}����p��l���6`?�4�#6���6�D0�4�^��Ƞ��t�q�����+�x��6\_.6�;����R�804�6���)ⵯ��p�R3Kx�B�6���5L5�6�g�3�[�4~�Y�W��i27@$Y3�4]�������Y6f��W6-N36�.'��D�5��I6����䴈�$5��O5X"�1�ݶE�5�6�M�5V� 6�(��H�6ȐC�1،597~��uu5�ڃ6��.�.���s6R���ĵb����j�6 �6�$�P����Z�4��F5�w��L�5��5�4�6�v6���M"��G6s�5ĕ���1� H6 :��C�5��ö�8ʴh��4�k���A5dy6�Q�c�k������5$Ϊ�Ё�5� #�XY6 W)5�H�{r%6��h���^��!�5� 6�#6�KQ��*n�&�'���5뢶��̵n>�5H��6��6
�$62P���Cy5 hϴ"h_5徂6B�����5<ߙ5��.6��/6xk6ޫ��h״�n�5�5�x�6�X�x�U6`14�?��M�)6���G� �5(i�5���6X�0��s���E3�#��16\~ ��&�#-6�鸴��48
B��0l��6��16 �o4L�q��m�5Rc�6��4�6��4�Ҏ�d���4�>,5�#6d���Ӎ&�����"�6�c6���4�5pS5
I\5��@6��;56汵e޻�`�<�Tg���M��u�6�k6��<���86C]D�x��4��5�:���4�6~L����$6�)_��߉����M&�6`Hl4�p۵�|)4^I�9*�5dP����ٴ�-���K�5DTA5ss����5p
*5���6[��5�����6�U��Y�%��5�ؑ5�ꦵ~!��Ѝ+�@O�@��z�6�6W�4���<��5M�6|�5��6(鴴:��6�Lz��&6.Ú5 �:4��6Rb6rܖ�@Nr�:<���҄5\87l傶��64 Tm�d��%m��:6��24�@F6@�������H4�j��5��&5U�5��#6�qT6h#�52*6���4 e��mr6� 5�q�\�#�qA�x�b6ʻҵLZ'5�>`6�j���KP���i6|^ԴěX5~��&����3���4#pR6���57���e-6v���{6 �0��4�֒��6�+����i�6�
!�}�1�7��6������6Xޓ�����8A�4�	6�ִ�Sw64��56��6�
����b���4� &�6�	7�ӽ����6FG�6"}�4췲6��5��7b唴�4�=���1��.���6�Ι6�=�6C���6��4�9w6�!T��Mʵ���5n|��uö�t�6���5�}&������Q6��8��	�ȴ�6�R�3�l6������+�Ď��&����(�6��S5eb�5�Z$�)֛��␶b��|]�4p&5h;���06w0b6����푤6�B��W�5�6�M64���F׵���7L�|�K6��e6 ^�6�9�z4
6j�6��m6"�5�ȯ��.5��5�_6��36��o�j;5*0$6��,6�2=�j�36����\Z�6��*��l8���i�fi��c��A�jگ61X��`�����L6������"6:e�5N�¶�'�5��t��B��Ԅ6^g`��Xa�?V�6R�5n4������7T�"3E�����RK��U?��f!��t-�n��5n��cx6����|R���Ҷ�(�k#���=�ր6K��6d�5c6���5`G
���|6�h���[77��Ys5"-��ܛO4k��5+Gභh15�޶>x"��� 5��D6��նx7��4��!5�;�6��w6�?l6�]6���6~*յ*ƴ6 8>�Iݎ6��<�� ��!?�6��� ��6'e6ai6V۴�A�!6j\I67SS7[0�5H��5w�+�`/{4T���Nj�6 1�6��4��7��6+k�ړx6��7�6>D$6�\��`2͵�!�@f65���]�6�訶�\ �́�6x�T5��c�k�W6���4�����`6�`7��6ɍ�5�C�s����[%6�{y��>ȶH���Ն��GE6�6� e�2v%�K޵$��
`�6��������j����[66��m�Ɂ�6�ש6^?����60O�	�[���,���O��ˢ�F`����6V霶�菵̔5"&��*�5��Q�"�ƶz�<5��ֳ��~��)�Y"��<��6����-%����6!�|5H�7®�����8<�66�7��6���5^�4j�l55Ɛ�D��4��2�f����6�%;5�e6?��ܣ�E]ж���6y�06�j50�I6�0�5��b6Xz���p��h��S,6�	����\*b���ζٵ�5-H6<��9.5T�63�-�t\����r���5jJ���A�e7���w5�&6���"����6܄*��_ܴx�|4K���n��6���6��O��9���A6� 6�6y{��D�6��Ĵ�G۵�?�5�J5��<�6*���&�6E�ǵ���5����>5�Cڵ��r���a6ķ���� ���R�6�u���5~�6n֮5X뺵'�E�y����c5��.ؖ��_}6l>׶R'����4���5��:6���+(����5�Pg6�ܢ��G7í36VG�5����H�6�i�C7	6&�U6E5��)6��^��C�5La��b�"6 Î����R(��<85��I6{˶Zʜ���R5�Y�6�W-��'�5-`&66��6��i���E��K�6g��z�6�D6ʭE6<a��W/5���񦲵?`��Z�6�=����5p�W6�:�3��6nD�5F�6���A�5��1�|
H��@��J�6h�k��o�6�W�<E>4�T�6@B�6��I6�J���L6�%�Kof6�h6�Lp654�J�E6�A�gV6��5�I������h�6Z
4�)r�A+�6�K 6s/�6r�����5�I[5�Ѹ4�����Rބ��[��|(�nc����g4f�����67R/6S�J6�x6�(�4�ѵq�ϵ[3���n��F���n��\�6�m59 6H̘5*ţ���5�i�[��5�6����	�5�cz54\���P� ��4�Z����4\����N6O����5��23�5�5�*�5B؛5���5L��а��D'6&�㵐�;5`m��N�H6۱W6��\5-:9�Q�p6��6 �=� ��q���n��+�6X��5x�,�L�4����C��d�v6�5P�7�R5�x�����5� ��{���ص'�)6��6�ء�I~�6�#�5%a5bJ��>T���A6�	56�	�
"G6Jэ6�V*6�J����P�Q6Hb|���5l9�N(j6j]:6�T6�F�o���d+M6�6�'?6o�26����������s�]��5�W��K��V 5ոJ6�1k6���:ߵז6$L�6�"]��堵]��%�6յL��56��0� 5v�3tכ�똃6V#�6��6�$����+����	�@���=�ސ�6�>�6���6����!�5? ���6����V�I5�U�@o���O6ͽ��2$^6��48���6�h͵Gg���8 6���� 8�1���5��5p��a��6d��4��~~62��5S�Ķ5�b?6tk�j}K6�ֈ�����M���Ƭ���=6�S"�4Ⴕ�w���"��+\�.^����6Ku>�4�����6�A 6�锳��y6�V6D����z+6��s6o��6f�o��[������&)����5
�6
~�P�r4S�j6��D6�pݴ�^����%6��I�4i]6
#�4�3���ރ�����/E� #�6����&6MW6�7Ѳo�l���Q6�Q�x��6�'63��5P��<����#3xDF6��6��6�~��П�44?���p6�b��]q^6j�7��5�����5S_���94�N�[6�J3t��p�y��*���}2�_�6&���;��ې�p�=6x�]5��k5���55��5�)�5�)�6�ד69�N�������)484���Ƕ%0x��G��r'���p�
�d�".�6�++�<�~��5�6�]w��͙�d����4ɷ15
)�h��6�Rd5��6r\�6t�P��?�����6�j޶Ʌ!6�6-���㙵�D6jC.601�4� r6 �8�Nl��o��1�x��5"�64퉵������5�J6�D��R�5��5E�e6~�h6Г,4ُ�4(�85a6�`�5��R7�6�f4�ٵ�h0���4�?G��2�4�n6J���I5�t6���ȁ�6 [��h���J��6Js4��6P�ݴ߾9�ְ�6�@���T6w�5��6�>z50v�5��>6�跴pH5��ϵp�����H6��u��ɶ��"�6���l��6Z��6��y6812���5 6$�Q6�AE�:�>��@o4DXQ����X��5V?�5r�"��6:���B5��\6{Oh5֛T5������𵒉�6��%�@�k6��76�6bD'��ӵЄ�5�9��t�A�>� 62N5��6����6�8��F�4q6x�=�����5��*/5xS%5
�6��Ҷ�(�4�R�6�-���-���_���
�7.96ʑP� T�5�J�5���5W+�\D�5���5�ڏ5q�@�NQZ6 ,�3d�c��D3��.�7 5���6([����@��d6����6�e6��~5S5�%6^�,�[p68~}5D_����5յ ]��P>P�pmG6���m5.W9���5��5W��g��6�S(�$���s�е�v�� 5k����4�p5���|p\5|�"6���5}��5�8����6���5���D6����*?�Ze�5 ���0�6��6���tϿ�`"�5p��4���5977���5� �\�[66m;6H_����е�-M6�<;6����60�Z��h�l�5 xݳɠ6����߶��4nG�5�מ��[4�:��N6nq�6r �6�O,�t�B����443~����5��6~9�u�QcK��ɸ��时�g����6hy���6�.��K�|���+��i6|5�$T���&�5�P���^���6��k�|*�6�ͦ4�x�6^�S���x��� �ࡄ3���5��h����y���L-��/y��w�5�ǆ�� 56lB�6d�75+X6R��6�����P�6p��4�Z6Q������_5`K��T��ɻ5�|6=(�6�a}6�:�6 ��6o�6d��Ų����6����
� �D�0��������٘6� ��E�5��>6$n�5{6��5�9��^�I6�+�6�v���F���=6�"̵v7p�T���6�X���U����6 �D5�D �ߍҵ`�4����`�6b��6��6N6v�e��.��5䇹���l6�145��6��ɵtՂ4�G��W�Fp�5?6����P��sϞ�����)�h	7�[��pv�5��k6�x~�*�6�,6��o6�h�����6��e�ʎʶ�8=5��Z�_����6���6���n�õ�㶍8�Z��(�36�ߵ�H�L���U6�W���6z(�6�̄�딹����4.]"��p?6��p4Ԭ3�pB�X�5\�E��6�R�3Zz6�p04
�p�|!���i��	ؤ���{�<�E���{���5��N���_�0��4`m�F���ޞj6l�6��w�N[h6X�5U�ᶨٲ5#�b6أW��[6C�6�~��"O 6p6Ȇy�B��5�p��^?6��[�LN����3�o�Ψ,6��9�i�z5_�4ȞB6���*=�5r��C�G6��76����T�6
�/��d�6��q�)�66�Ʃ6Åu6y9$5@v�4d�45įK��H��3�7��Y�٦l6)#6��4��L6��7c�p�԰�6,)6������7��}��OW6*u��A��6��5����'�6	\��\86�7\��~�5>�6�e��]6E踵�)�bQ�.Zʵ�:�ih���\e6d�5^,�H5K�$��7�ۖ6(mP3�v�5��6#hx�������d6�ޭ�������6��6��5��%�N5~��������5tRе컃4t��5Xq{�a�G6F��>O��Ͽ�̫	5H��5�~��;�Q�Dʷ��������kz��bl�Z
7%�5d~�5&؏6��66�^7vⵧх6tګ�	)6��74Tv�5TQ��ϥ4"�6��6+І6p
�[.�6�2�6�@���c,��f����52;��1Ѕ���p�}��w�i�xO�6��z60H��>�6�I60�4j{'7m�Z6�x�d�!5���6K����n5QQ����j�7�����t6|l8�K5�C�6�7¶@�6䇴.EA��]T��i16X�s�q+d6nR���3�y�6p�'��Ň6(�~�TV�����x;�5�6�Ķx67��6�Ђ��ӟ�@�A�8�6��5�)t��E�5��5��A��϶m��6X]5�b>�ڪ˶-�6(sa�h��4W�@� ef��v�6pA@��W��b
K����6���6����vה4|ϟ5�I��lݶh��5�dh5�x5�Z5#ݶ���4�ܶ]B�6�@6VS6X���'����5BѪ�/��6$�F�6`�ڵW��	������6�_T6ښ�#�6r�5`�5�d6bz6��6�~3�<��� ��y�6^`�6=g�6�`6�[�-u�6 D,4L����>^"�֘)��Y�3�)��������家Kb�6,��6�Ҿ�_I�5a �@1�60�?�.�����6,�I�]�ն<޾��5���N#3�?i6؃��|���2��-58Q�5����t<]6�Ƕ����t�vA�KĶ���6ĤԶ���5(�� W�EJ�5\�@5/۷5��ڶ\�64
w���5\�c5�}-�^��5SZ���Z��ِ�$O������n6������I�`s��gN7N���&�62�6��+�3J6ᮗ6|d �p!�4�ج6?���ZP�QV���Ԋ�(�̶����E&�ދȵ�`�6��߂S6B�6[5&��6�{����366&ٴ(;R5�
6��6�Ķ�-6���5�l�6̫q6�ǯ46�M6��6O3��56ᶦ��6�t$6Ɓ	��77�����5���U@���5)DP6�g�T��Y�8�;޳6�|4��6A��nO=6�:��=��q���B��H�5{2�0�r��5,�5�o���3r�(6�a�5�F��6@����\6J`_�\ �4��s6 H��Q��
��@�
4r��Or��F"���f�5�3�5�"�~�����������60c�4Ζ[5��E�5��[4���ϝ�5��T�[5�55�5�5�ͳ�˖6.60����"J�rOյ4�p5��2�B6<Q76b76 f�f.c�X�X5�û5��ܶ(��36K�&Y5�9ӵ�?�5�5�4�9�4���A�pt���X4%{5��|���´�$�(6*���������^�Z�56�6��[�e����ӵ-���rC�6��7��7@u�4�%5Ȧ�5��y�^K
6\0Z��H6�# 6��4�56�y6����ó���5�I�� ��4 ��2�PK�N��6&˛5�w�5 <)4�ڰ��I2�غ=6��a�u��5}�u5?��=D����6�A6�AH6s����%"���76P�6|�|6.�¯5��M��M��/KG6q{Z����Re�6l 6�ǳ��NT��y���d6��6�oҳ�sk�|06�g�6]�5��v5
uF6�dgC6��k����h���ʟ�� y�#6��5�H^5�N�6�4�5@!6�c8�� �3՗6���5�,��~��_ôc�M���5�ʍ56����.�@y�4pb�4�Dܵ���5��@5�F&6X{1��։���)��Hm���;5�P��G66J�5�퀶������*5j6*46Գ<6E7s5�hi���	7�^�5`�{5Jo6$&�5T��53T6J�l6�Y��lC�J�%�0��3e۾�-���D�⤓6�[�6]2��@O4��68Jf����4�5�i�6T��6���L�J6n� =f6��5�@t�n��5��v��u��@��)n�6�E�5�jµ�-6@�մ�'�5�Փ5X�5��96���4�U�6�6ʨ�4��C��k.�Fd6�!�6��q�l��4��4 �b� ��3�7��\��5��+3&a�4(�@l/�N뚶�8����2: �� `	6�J���V5x�5���p8��r�w���6���6I����|�7�5C�񠑶|�
5>�6�"� 6i5!�(5�v�c��|��6�o�36nؒ�0˔���	��5���4���5�z�5�D��$�*�����66��6`�5�e�G���X:���4� |6�؂�`{�3���𼛴?�S�@M��ă ��.6�5�-��s�5�+,�����l`'6`�H%�5�v��~��5��5x�5Q �5�ϵ��~6��d5RZ)��w�q�&��5���nK5�}̴T�!�ط�6����bU�5@�k�z�9�5U���"]6��ߵ�
	�(�4@u�6zm*���'��r��'n�`<P�zT@6M6�)6 X�L_���{r6P�5��5���6H��4쒯��l�4��45<�6 �T3X�6��;b�к�5�4�.5������5P�����4�|e�h���b(l��Ԅ5�.��*��>�� ���;+��'*6��pw�\��@���z���#w�5���5ޓ�5�R�5���4�lP6$����� E,��6�ч�JC���i�8�l5���6�f64�_6֊���]��<�6.6g�8C5[�|6ro��L �5{�5©
6�P5f&���L���.��%��W0�������KB��	^赴ĵ�M���窵���3<j6\�赼��� X#��O�j�y���l�0
76 d�2|��5%�>�׶Ą�5�3��o��r6���6���䈵��4�����J�u�H�+���ǵ���5)GI���5����rPe6j`�4��еh!5�,��O���:6�26gV6�q��@!&5N��|j���6��D�5x�5̷p6��`|c�n�~����(26���6�?��0�L5��6T�5��6�9�<�6X*6������Y���ݴ%�_��2��,���16 [�6�Ъ��<��T&�� �6��!6�&.6��@5�������4��21�z������n5s��6��6�$��%2\6#��6�"�6D�ö��5A�������Hȵ���4J�P������6<z[6��r�_&�6�B�5{��)6"��� R�4���4T
�6��p6�(:�)�5���5�7{����6�f�6�v��<��z8��,쌴�D*5 @��S��X����L �2��('68-��9?60g�6~K6������ �2D��6�J�69�:5��
��Ӆ��c�5)���7@ݶLW@���5�@�� L�3v�Q�o��5�� �v��Ԣ6�5��V�������d�e6䩛��=6Q3�56P�5!桶H���@��3��6 	��k�S4���e�M����$35F}{����5�m6���6%Yn��I�5��7z]6��F�^�#��'�5`=�hjk6�u�5��6J�%6� A6��6�����N6x��g@��۴T�c5hH/�ὦ6���������52�5�1��*�T��6�6�P�6ɶ���3�؀5�⃶Qi���4�Z��6���6ʄ����ҵ l'1���5�ӊ� �@�+r�6�G6H+ֵ�0W6�[�5�ɉ�6��s�927���PQ��!�ޓ��7�6(ܣ4ׄ3��ڜ6'�6T2���#R6�!�V_���ĶP[�6�_�Pϵ�p#���Yi5�,I5��6�.c�D�6�_��z�ZQ|6���ҵ�y���*���Z��P땶��������!k4X>�60��1'�5`���d5P��|�4�ٴ6n��5H	
���6�uI�%HO��.a��j�6�vc�f@6�~�4�L�6��78Q���a|5 ����W$�>��5�����@��2S��Yŵ@|K�W�6�>�6��6�ȥ6� 7�x�K��5�]�R10���T��f��6�j2��%�5��6�㉵���4XU~��ȵ���5��=6���63I��Ʌ��V>3������E}��t8b5U�}67h/��!D5AJе0�I5�6���5,��z&A��m�5��j�565 ⃱�ܵ����袵�ɔ5�.n6�t��׌u�*�5�6��e���sY6�K�TX�4�)u�F������|4hv�5��d3�E�5ɹǵpa4�H�4�v�4Y~"��Ǔ6(��4sR+���e�46`6�o"�5@�<3\2?�X�����U�V^���X5�6}��1*6nԯ5�5��#5Ƙݵ� w�Ǹ�5��1�P��4�,��4bD5��{6$C5���5ʎe�ҿ76896h�ݵƊ�Z�T66@쵎]�b���Q:�5(�b��5a\�5��y6&V�\`{���o5J`鵥?�5fҴ�@����z�%U6n��U�]]�6F)3��=��0�
�۵]����66�u�n�v5NKɶ��Q��]i6H�-hZ6Їb57����� "S��e�6���48�����X��5lW��O��j�5�B}4X_�mj�5@��3��ߴ����Qv6�A6t�x4�4L�+���-p��[��U6�o�5L#6NʵO-�Hk����O5VR6�ڊ6�|����q�B���b�D�2�ƵI6�50��ظ�4����	�4�
�5c�4�ȼ5��9�����!�5���4y��\ v����dڵm56�6��4��6�P6R�~%2�@*g4�b�R/26TcA5�� �I6nO5��� {��N��P{�40�涐X���� �:Q0�G�5���6����T�4��3�����3`�յ��i�r{5� �4E���uw5 ��5�cT��U-6xڄ���4"�����h5p⺵}TK�\N6?��fǒ5���5�����R(��<`7 ��5ԕ��V4!�'6�fM�r��6� /�l��k59�R�6��\���մ��:��í4��6WQ85�QL������v��D.z6FV⶘ʺ5Xd�4C6�6x,m�WX��J6B�q�B̞�yHJ�L�W4g�Y5cE�6iJ5H��5��&6]�\7׵D�����9�ŵ5c65��*ƈ6k_:6����������6!�6�k ��6,�5D�5I�5�ݟ��Ì4|š6($R5��*��.���d�5x�6D���Ǣ50�j���&����슮6 �� ���;U5[a>��	6�J6:�X@:�,�S�����C5���2P���y�6z�5��5�4�A�5l�6�%�5�T^���{����5S55�25[�5��x��4�'����0���x�R�M5�em6�r�5DL%�}lu5`��3��дpV�6�\n5-�2�����!5����B3�@�����=��� 6x�(����5�&5@���X��,D	�8*85����\жP��3x��5HH����4��X6��3j���8�56��6a��6 c�����5p�m��BT����5[T�5 pM64��vE��=6�'�6(ն5�36`��5:tx���5�g� t�4y�5 �6��Ƌ5�w�A �����5�� 6�m>4�5A�4�;�|��b��K4�6����b���Aa4�6�V=�X26���0�4�t5Ę�5�wq��sI6`6��4�[����V6t^59�4���<DS4�_�^�&6�Й5�4�;c�l*�5�y�5�E�6~�!6�i�4�Ie6��ǵ0�5��D3�C�4Ȍ�6���5�=6���5 *8�0Ub5ƦT��H45B�o���6 WL� �h�ֵh}R���U5�Zn��Q=6x��4���4�..�wl 6(�"�;h͵��5�J5�6��5������ѳ�b���S5�n6�[?4Y4.6|���ާ2��+�X�ֵ�T�x�N�p6��Oa�:���փ6��5�n�5P�_4�TF�ᘶof?��H�����xO5Zcs��S�jĠ��6]4�Hյ7��6��25�Y�V����� 1q������5k��yJ�� �{��S>��7�5�l����ٵ�\���F|�h6��L�/B�2r��o8�w�6�� ���8��5����>ݟ5P�y4L-����5�;7��5ɊӶY��@��3�l�5���{6�?�5��%��dյ�7t���066�6G�5���5�CR��]5��6�"o��6�zJ�.L���a�4��=�~ �bQW��q6��N6i9���u��#�t�p��6ۮ��O�6�m+6�n5�F��Z�?�n5'46K���Bn&7�c����6��>�vR�{�79Mҵth.�߁&�6R�5��46��47i�6�Ӵ����@/���Ƶ���5kk�6�ܱ6R�5H[/�Vۊ���ߵCÛ��!��2���E6�E��/
16Zǂ����56��p��6ŎT5��ȶ�B�5"�6|����5Z�Z5�}�5b;�50�x�0=6��6�<_��7Ҷ�6��6L�p�b^5Q�����5fI5�"k5N	5��+�cc`5к���EW������5�͘6���5P�5���4�f4������`6d1�6�A�4BQ�
���R��F$�5^5H��CV�5�h�5��6�[��A;]�6�e53�5�j6���5��Y5)7�5@��XR�~޴���(�q�[��6��5��7�+�Ϝ6i�2K��a�6�.Ե�j7::Z�᠁��!6������H6ҥE6��̵9�P6�	67?A�Nlk���6�6�y��WXy�&R��?>���!���!6�1�� 5�6�0�4y�a6�x7|�����Ĳ��8�5D�7�DV6V�D6�1r6̪��
��h6�W�6�"	����5ı6�A���Ƶ��@�n.�5Px����P6U�"6Ge36�7�p�3��j5��T�66�tg6����S�ܱ�������6���6R	�5+z6��6h9�6r�&5�1��5J��6�6�6z�5�W���I6����_�h�C�vz�5�0U6ؚ�5pT��N�$E6B̥5X��5��5��(�
�e6��w�����k��?�6��2�ʶ%;�5c�5�e]�HF&5BВ����4�6�Q�Q��؈�l6�4{D���eK6V&���6ra�4l΂�|5r��5�:���%�hʀ6��f�t��җ}5������6&����d5����߷�5�I�5P����(�-�\6�,���� �P��4��5�ʚ6ת�6�˥��*��6ʊ��s�6�����(��g������M��nd^�<\�/0��<H5�b������#�5X6,5�
�5}]���-c���z4;r�6�g65��W�cN6�n[�'��5)
36 *崞�}��݁��V�P,W6X�ε�	�6�6<�6"6Te��L�5�=�:�'6���5})��05�t6T�2��Ȋ� ��t%����ʵ���5׈�5��@4~����A� T��r��5d�ڵ�Z+7�5��r�U�6��6�c[���7쳈,����6���Õ3�H�5J���:��6 �鵑����0f5W���"�_6�Y.���5bL�5@I�4�^�5ꈶ���6��f��(�6�j^��Z|�<��#�6��=60����޶��6X��䵺5��cĶ�M���n4X��5"]�""6&U�5AU6����N5,��5 >6.]����6t��&�v��T6Ə�6�C���ٵ�5�3�5S����$�5`���5�63&���ګ��Oz�����-K'�`����:5v�������=��6N����6�\���Q���C6�����T4&�W��N�6���5��5�6�⁵A����m��;q�l�a6ptd���^��m5P�.�L���p0�4l��4�傶�H�5L/�5v?P6bC�6 ��3��4���5!�� ��5b��5P@�5��1����V���Ձ5��6R6&!�5~�6?Q�����5�V�4����w3nbе���3��5��3�M녵�L�5䦽5أ�X�k��͈�"�v5��V�,L�5�>6�2�b4��_5]�5��6���F�M6�P�5b��5��\�P���+��6�hS5���5�څ���V54��5M"{5�p���S5�J�5zІ�����14�T�4�J����������Q6 :�3��5�0�5M��p����4z6&Ң��t��մR%��!�4P��A�i5�4�4r���t5�T)6�H���Y4��#��4
6����,m6��5�5�2��5*��w.��]�5��f��j�5Xi[�|05
/5�L}��;���)4`�S����5��
6j�5�S���`�3M�õ�?�5G�6�^����r���	G50��4Z�5��5_ޯ�$�����Q�6��ĵwJ����3AL޵/d5��2�X򴴵U�5*�5��4��~5@�=�kٶ5��Q��/6�ާ3�D�5���5�B�4�f26ڐ�5��J���5�s6�#���P��ې�,�ȕ�3���5d�>�P�$��Ay�H��5t��5��?�5�q�5f46I5�i�h�3l��5��6!]r�H���
�%�5�Mt3�l4�u�4=�5D�$5BoN5��5R15{k�44Y9440ɵFֿ4�x�5�.��U�5��3��*�67K5�Ø5@�>5Ԗ4�$<4�S5��������w/5��y5hr���K�����PT�V�x���4�{6�xd����5A�5>X��w�5��s��G���&�4�*�5to5����,�<a!�X@4�5G��,n�p�5��5l۵��>�Lk�4�.����5=��4���5��	�o���,-��~�5�
_���6��5��.5n�59�$�nJ�� �3�P6��3=�u�!�4�͵W�j5�ͱ��Lm��6X�ӳ����9	5T�5r�C6�7�4g��4�t��%���������5���50�c3��(6��4����5��6�y�h�`�:#�5@JT��;����PC�5 ���r\?6@�P���@�5�4� �xb4d�-6��"6�h6��\�P;A��d�5�S�4�*��}�5d|O�.�;�f���T�66�6���fI}���X��Ȥ6/XR����B^]�"�6��E6�϶��/�4�_����6�T� �3q/6w\�5��9�)o/6��6(��"7�;r�~]c5��86Ɗ����5��m�@��6N�R���O�h�;6d��4��"6�7�"*���l�@j��悶,ę5 eW��Y?6S#�6��/5"���V�64[y6��5�V|�r��6���+�6@u�4���6= [6���55���v<6
)�6(��6�������5��86*�8�0��5��Ƶ�A���72j&6���4��6`�[q�5'����e�5�ٶ�ޜ�h��5Z�5�6N5
xܶzڤ��a�6�6n^R�8��5Y�5��l6��%62v�6 �4DZ޴����(T5�#�6zK�Ѝڶ}p�2,�f	q6h35�W�5���6qM�5b�!���6٦|����5������˯��>c��H��6�,�6��(4b�6�۶�� 6��6�|C� �3�b��/ܬ5`�T4�B��-��8��,6&����#^5��ö^���B�66���6��%������v��V*�6h�5�-B�*5����P0C�5S�(~Q5�~C6He�64����ܺ��+����r6�}l�4�6l��5�^���d���m6:�;Y�6/\w�o�i6�w5��Y�����5>�Y6B�V��=���!6i�<���굸d@4���5��9��6e�t6T���iJ5�6����Y��/����5��Z�ϭ��↴�ϒ�܈56$�%5�Q��[3�5t����U���6����H6�, �f����/ϴ���5�j3�`'��76L�3��V�C�:H�B�36@7ݴ>���G������<�4��u5�N)6��6��c��3���ĵr�d����
����ݴp��5d�@���\ҹ�n�,6���6�84�GQ6H)�6��U3֏���5�6������6��6��/?�6�K	5'&$��=6^��5&��7<��zջ��ɴ�5��+5��49��5Xs�Vb�5���U�u�N*6����f�p��$���6?�6:����@����8?�4�0�5����f&�՜����+��F���j�@���0�6�|T6��$6:6��$6�7��Ky�6��6�rYٶƪ���׬6f1Q����6tܮ5��������7�5@d��w6j�P�@�;�zz�6���.E�t�#��5�"4���Y5��6�~��%y�5W�6ʍ��
둶/������5 Ǵ���+6�!���$7
(����6dYɶE��`д��Â����5�?6�
4��5��6��6�V��Uw{�E1?�(�5��
���!�̻�5H�5z��6��0@޴p��5Т䶷�ʶl\��ԓ/6�0h���߃����6@�4?��_76�6�`�4a�o�������7��6L����\	7 ö����5ۡ_�Rk��>�4���3�>��ʶ���B��NF�5����@�µ�Gm6P��4�n�`?t�Q��65��5�	ٶ�D����	���d��.����A���"ER�����x��4�O]���5h�������&;`6p=�@��3�55U!_�ɑ6��7�<Zb6. �6 �\4�.#��t��K��[��`XY��7J�&�D���Ң��o��6M@g6wo��l���sU�b�t6<��h�\��Kl6�(���0�2���6V�Q�P�4���6�D�PYB��$� ?�5=P�6�-6v�z��.i�5�����5��a6�W>��Z�6ܞA6�sζ�P���xIg�.��%���"4ʾ�6����5�/���F6�"ƶ�X<��2�5�#U����5��4.@6B��5P�+�$�ﵒ �5�����6��l��{��Ͷru��)5�c�5)ŵ��$�@�2��T5I���1�N6�^�3�����4���5��4��5O׏��f�؀\6U~εK����F5�]R6�a<5��̵�̤��P���6R:I�-!6@���u5��5��s5:텴XU5�6�"�::6�uS���ʵ`��4{5������N��d�����@j8�	���B �5���M���&I�x��I��5�w�U]�5�9A��Eҵ]ON6X6����=4�6��5>�K���x��:#6���� �6*��5�E��i�ܵ�b��]-���ʵM2�5� �6�B�P��5�����R��L6tt���S��]���O��,x5=�54)���D%4"�z��A5��`4��5..52u5;/���೴�%���"�"5@�36�[�6��5���5P�3���5Bߢ��E�n3ǵ՜6�[6��� �5�`�5.U6�v�5�k�B@?6h�6P�=�zt�5���2ە���LA4c�5(�ǵ~��5_�൙~�50��5dY�56�6+�5g�4��Դ`�;6��A�V流j�5�[�� �6+�5 5��=������ԋ������:µ^�<5�����6����Y�	�%5Q���:�3�d���5~!7��O��zQ�6�hK5����!P�l�4tyŴkϔ5�My�vr��
���4H ��R�-���m�6���5p6��zV�4����6��<�&6 pճ�ߵ�����e�}�������A5Z��5z�䓽5p���fJ�7��� Ӳ���4[�#5���4n��Ig6�.5�O(4��	����5ͷ+6�6J��K�5^�s��C�J�����'���L6��d�K4̴���؅E����5������jL��M�����0�D��䳶5\�67�25$��4��5K��V45��5	�6䥍��+]6�~'6�o��!�96��U5t��4��5̔<�%f5Y� 6d�=�Fw6���3�6P5���5T��5@��YL���t6�}����̴��J����68����5�6N��ӡ6f���0�˶!�6#���höza�5��:����6��5e27N?����@6�����CY�5�o�?6�I�6[	Ҷ_5��p<34�����5�pD6�_�4
A�5r8�|6��46	�a7n&���W�6Ę�j�j5�\�6�\��.�O6�B�6mM!7�[�����{]S7xc�5��5a�B� ����n6�{n6Բ���w,7͚T�бB6M|f6Y+ֵS�]�`�5E7�bN��̶��U�_�6���6���@Գ3�z5�~�gc�5Y�?���(6�!�!��5}��B��� `�6MS'��5���𢵤�	5�����C�5�4����6�;���k���K��c���3�17�M�{�
�>�.@X�`2�5呟��"6;>������ �w�6k��b����,���`+ֳl��6��o5/�� ß4�'3��c6�o6���A�k6J���ȓ�N��5���6_��5˧�L'ͶE� �F�6Xx6���5R����S�6��Z6��1���h��67�c	7|����5�#�6 ^4�lv.6p���� 5w�P����B]�6��>Џ�hD� ��6�K5�4�(����"6�����p=6[iֶYҤ6u����5�(������j�6dR�6�1�6�/�60�ĳ���P)�6�P˶��@64o�4$3d�tX'���[6|.��V�'�DOX�\X6�T6�r�����_Cz���66��ҵ�p�����3���:�u�J6ؓ�RF�z�Z��%�&�ض59�]d45z)�5���,q�.��F�6DHĵ��T6��6�X׶g�6�E-4E�]���M��GA���.6�Z�����v`,6����	6��6׏D6�X�6F���d�U�������6(
,6\/$4�ø6I����`�� �2�����4ۚ��ʬ�� l��6�8�����
7�.f���6��)�H4�(_�6�۶:������CҵX z5����n6T.U��y����6�qζf�)5<ۉ5B�A5Ԛ����6%��,�µ` ����C6��*쨵·��b�����6Jtζ8��6a�5sd�.Q�50?��@�7��T�v�����5n��6"�5q6)D�@�6��5bS+6l�˴@6~�0$n6���6����D&��'R�5҄ �!n@609���7;5���6�����o���s6"J �Peq�0`X4�֟5��E���86��o���c��a,5�{b�#7t���H16_�5���5|�a5+�4���5�����Ԕ��EU6��6�77t��4�N6x�Y�+b�6<K¶��6XT����5`s�6�o6�S�5b�3�}f5���6B~
7�d�%p��F �f�g6��O����5�S�?�L� ��4���6~��8�j�6��5���5:q6��?��´���6%�Q��:7���3��ҵ[����@E��}6\��4�Yd��M6^-d5�⧶��]6�U6<jʵ�q2�*��-��`����6�G%�v5��P�;6�ք��d�5P�6^ҶrS6�y�����H��S�,�:Jc����>6���6}9�6Z�D6��w6��5�V����66���5�����Q�6Pu����V5NY��FP6]{:���7Z*6�`f6�C��r��{��6��=5&���.�@W6��<���M�HT75J�7e(���U0�p��X4�"����;������4x�?6�5��6ُ�6_Қ5�c�6ZM���6�6k���}R�6�s�6��6@`յ��6��{���q���7XV�6�d�6a{g6J�56^D6�R�H���o� ��6 �2��a6d��6���5�Kp����� ���(�5�.���7�I6�ϕ6W�6������6��0�.�6���8�^5(_l5�x4��]�\�6`<X6�,7 ��3�u�6&��6b�x5���6 kf6O�-�IF�5(����씶ds���b�q΀5���|��4�ʮ5����wϵ��25�0�Q�K6��s����,�4�c��$b��T�3�^]6��6�h�_�X�.N�6�y�5�k�6 �6rߵd�b6V_U5;娶$�S��0��s{��5ƛ�4�_�ň�6�4@p�M���ʭ6�+�4��@�3�u��5 ��� ;��Q9�D�'7�|�� v���{>�$ָ5{pᶃAy5���6S�5�5����i���k>6���6�56�:5��5أ`�]45�]
6����*H�6�r�5��6xt��然�iϵL�������,6���4�RR6Z��� &�3���B�p6|�<6 ��0�KM6u܃5�ï�`��1��6�2���6 �5/��4�ki�s�6~�6�Y�6`��BI�d�f5�X��xv�5
�4H4@62a5�#�3�f��<�5ք�6D����t/���5^u�4�瑶���5�U�p��5�bm�-5�����58�6$񒶉$6�R6hij�κ��V�6�բ�k�C�����o��Ȣ���6_8�5m��6�Ac�j���_ ��L;���6����bM6�8(��ܨ��k�ާ7��|g6B/�5�7�4{�5\?�Ɉ�5Mo5mi7������7����04�?���糶��'��r6����g�5qj�5h�ܵa�U6�˵�V&��:��D~�6��5u��!Γ6!7�5�	�6EI��$���@�E6����nමX[���6�C�6έ{6R�5�l��6L���R�4%p�5�+?��Y޶'���1�`g�6��+�1z�5hB�6y�6<�e�e営�6�[���e6��?�#�����6P6�J�527�6�<>�%��5F��6WFh6�r�j���PC�6���Li�3G6�i��65��3Y\*��� 5u�6Ҡ&�§�4@n��k/&6��5�Ut6�Vx�_�
ٳ���5D�����6r�56�O�Tܒ6�e����5%���f�5c�74�7����������o�6��r5�剶���5�r�6�Xr�Hz��6Z��~|���y6A�������@|�5�U�����5�_%7@���5&�6W95�tG6?T	6�&g����� Y3����0�����ZF5��5���<e��>둵��H66쌡5���6��	�>V���TQ7�].�B
���l6�R5�=��Daʶ�{�6��7���6Z����6�7'�6��6�T�6pA��|�j7fO��><����7e�6J<54L��ε6S���(᫶�%6��O����5�5�I56�ɭ���B4ǿ��ZJ�y~���0;�kT"�f�>�ȑԵTE����76`s4�^̶�<�6���x�(5�O�6�s	���Q5�N�5:3���Z?6Pqz���k7y�6��6��]�������6�Ї:7�?6�ʶ�J����4\22��99���66|뫶��ֶ�)	�0O�6̱a6�y5��ж~�	7��Z5*<���
7kR�6��P6@7F6r���x6�$;4'�E6"���i��04َ�6�YI����6��s�Ȯ���X�y�YQX6�#ڶX��5\��6Z�6�Y7��d�8�7Z�ٵ�g�6�Z��Uq#��B�6|�5�H����!6��]6��5Kj�6y�)�R���ovW�n�~�#ҵ�����P���6k�A6�e5�d�6 MA�����6��r6ď�4���6v��>_6�l�t8�6��34��y�$�ζ9�6LP��#7�g��t�6�5����5@�����춬/6��;5�t!6�9�8�q�ћQ�#���iY�?��6�yX6<�6N��5���5�is��h5�^6�յ�\���	��5�n�5��a��~r6��9�`n%4d��5�U2�p�5t޻�G&��N
��}.6b�36%D)���:6|y˴F�5A�ﶇs0���`6r�6�-7��P6q�S6(���4涶�86n�#�7��Ӷ9o!�E�5�U�� �e�FR5�ϼ5~�@�y��P6�����b6���Ĉ�|~��v'-�J�����6�Y�5�F�61C� j5&{a6��	�pT�3B.��,7�]N���� ��2��b��V�3D�l6��
6N5T�;�:�`�6W�6�4��a��5��5�tO5�	�5���5�&�FX6��t5�_5�k.4؄������r$K6J�D�p�'5�����n�;�6 �x���0����eܶ�f)5���5�x�5KqݶJq���6�������5��5|�5b'6����ضCI�H�n���6`�}��>e���P�0�5��&-����2"6�S���Q���#�5�6�h63����u��7���5ַ%�t���r�����6��Z4)j��W���x���7~H�5��5��6ش���
�6J;6��.�"�5��6[���C���g���. 5�p�6�/|6�C6�Q���S�۵|ٻ4t/6l(&����ƫ�v3���v���ƴ8��6>.˵>���f5��е��ᶣ쵸��6�"56$�*-Ӷ�lZ6s�ʕ`5��>���
�6�yq���X��J���䔵
@o6�#y6�C5�m��ñƶ�p�4�c0���S6?����
6�]����9�c+�5� g6�4�oe�6@g�4�5�4�����������B�5$�m��f��*A�5@�C�Tߵ�"����*��6g(�6o6�%36`�94��6����9���o�06N��UT�ޙj��5.l�6��ʶ��n����S94b15�L�����G�6-�w5t�5�S76j����M6���6n5�6�'�5��P����� �=:�6�eh����LM��hn��w��%/�5�صɏ<������6@@p5Z��
d�6�k�I��N�7^.$�5C"5~e̵��J�V�65�Ռ��=�� �5��T�V�7�x������  �����7&6m�5ޝ�]cI��Μ6⚤�=����@O��,�5?�$��;y��غ5F�ɵ '��$�b6w?�v��׿*6�{����+4���6��D6m�6�^�$�6�=���/5��H6�Zj��ȴ�\6.6Pv�5@����)����5�X�4����n�&�M5y	4��.���#6�����fu5����06��6� 4����5vy�����N��5��A:6�16��ڵ�Z(6h�/4H4o6���D���@?�4���6&�o6�y�@T'6���4ȓ-�\�ȵ�&P4�<�5��6Tǘ6i+����4��2��9R��};6��6\��5�(4�5�ec�œy6lq5007��6�5L�{�5��m5�ԵIX 6�٢5���4f�.6A�p��B�݈ߴy\6p����J6>�lO��"�q��%6��6��4�5��56a$46���I�+���,�26�����~�5��z�H�Z6���5�g5�FH6F�i�5,L6`�)60�3�a6�L��K6yy��Q���6~�6B=26�f�57	��Խ5��ԵL�	6��56��5'�#��0�5�o�5��l6�q6
` ���4\Gf��`|5el6$�ζt��5oH�
�5��4L����R͵X�e5�56�i�4�5ڵ��4�+C����5}�6�195Nt_�qӲ�;p6,�15Q�o���5�,�5Gs5��6�n�5@��\U� �2�i4"�6��"�()C6�v�5����&�������352���VP6do/��@z6=Vn5��⵨��5��96�' 6~�D�pHX��L�1b{��6�6t��5����7��5fa��U��Լ���%6��60��5�6#����50�*4�]S6@6JP�5l����L6��U��W�5��D����6�3�5V��6��M5{o�"%������6��N��O>5��5���8!�r�6���k6HzĴ�E]�z�P6{[6ֲ<6��(�QXq�p� ����[-�6��W3_���%w6�f���_5ț��L2ƶ�*6��5T�5$��5��ն8>����4� 6S�*a����C��\6� 趈���4�6.�5`L�� _b3��-��ۗ4R m�������5D +����.�����n6H\�6�/���*36�h?6_A6h��6
��5����U��H$�6pb5$v��)\�6x����m��p��3�C�5�� �/�f6On���5�j�5)��o|O6.
����(6۶c�"���*����?6�l͵�r�x���Cĵ��6��C6�96Zݬ�k��8y�5��r�@8���o�6�t�4��4�[�6�&$6��5ʇv���:60�
��6}��6 9�4�B�5./6VS��U6<-L6����RD]� p76Ĭ�5-Ƶ��\6�Aϵ���5�6O�6�tb5�n66rq6�H(�rb�5����6�����l��>5��3�
4�Q)�\z�������^��6�Y�40�����5���b(�6��d68j��nڬ64�p�N�6���v����O7���5p�A����5X"t���۵g��`Jd3n��4+}�5�������5~0^��R�6���o��z�1	5��56>ε�/� )�6�5�A6��5$(G5��6�'���9�5����'���q�-��5̎��dH6���V{�ָ�4��+6���5Z㘶��6 �\17F�Z�s5�t6���6�_�rv56^MA6�6������5�S�3M(t��}��X�δ�b���6&E�5yQ46�3���6��a�!z�5��6����V6 z�5fj�K6�Ć6dR��0[M4�u�b'���%�j��7�ۆ4�k_��=���w����5Nl8�x��6�&k���ε��6Z�3��u��2��6��A��%�3��6�Ƣ6�f�6k��T�568h����?6]����;���h�5����5 �3Щ	����5�ď��!�5[��5v�6-�=6]��&����p�5!�v��i�5	b�6x9D�<�6���5�\��ִ8"@4�E���6f8�^7���F�4���T�6�6�
6בn7������6�Z5�s��D�޵��6�6�}+�0��6�5���e66�~�6K�7n2G6�Ժ6��!�b͔50pU6��p51#��½��P��<6̶�y�6�K6��r5i�6U�6�&���6bF`6rO 6�v6B�6xeO���>�N�h�����@&7b�5�X�6�|m�=�;�~�"7m�66�6�����z_6���V�<�
7h45'�=�;� �y��4�<�l|�6�x��l��&��O�5�J��7|����5�7���5 Q�-���,@�Y�6xΈ6\���5��
�����Bg�6+ +�ٙ;6x9���6:��S���9�6��V�M�ʶ�6�]Ѷ��T��Z�5�8��:ѐ6�@8;647���zٵ�).���ɵ|��5<x�3�q 6���v�rm5���5�z����5������ٶ��{6��y���5Um�U��68yϴ(���p붰e�6"��5�!ж��5^y�6�t��ek�(L 6v-7��������C�\,�6)��6}z�6����X���6?��6�����za���g6΍d�к�4�g2��Yx5<�7�]�l�6އյ�n5�c���;����6O�$��pu����F�6X��Jе�����f˵j�l6vw
5��j��vM6Peq���6>�-��pŵ �u����5^c�5����d�Jچ���,6�1���萶z�6 X��|��n�7Q׵�c�#7P蚶��6��!68�+5%�06�Yy5��/61��4����
Ő4�W 5�����i=�����"7�5�ߝ�Vp�5�X#5��Ƶh��6�~��^��"O�6H.�5.��&x6���\��|�6�x"6�!/�t�~�ȴ��-�v����6X z6 g�2��6
\D��6\%��}�5��6	�T��~��GF�i��*�B��)\5���6<%�<���;T��;�����6��@���[7���F�ݵ���5�Y�٢B5���.�4��60%�3헌�ږ�5�p6=�5��{浉]6�b��C6�zc����5=��5R1��A���!�[��RX5ڊ����9�O~�5D��3#e26�6L)"6��$���޴x�6tz[5AW�c�5�"�5�6����4/������ �s��F�J��4d"6v,Ҷ��R:�5�k�579�4W�a4�i6��5�D��y����	6"��3�;��l޵qt�5�a�����5��8�
*�Ɔ5T�/��L]��y����5)9%6 �x0�l�5l.���9�5U�06.:t6�c65�)�4����Zy5�
��i�,6���?�4�G���5�z���I6��5ԅ���6���5'?�գ|���u��n ���6�����5���Pm��o�26�S�3�i�5LN���Ι5�愶��d6��!6 �3�]j2��6�yǵ��Դ�|h5#Gp�PX�4�����x��F�J5ƌ�5j`6d���5I3]6>��P�W��� 6M_ �.�q5Ȝ	5�x�,�V5��5�?����6P����84�56 �y���6-��5 㴧L:��浍�ʵ 	��M�B���6d���V��5n�5�4 5Ҁ
6�x�>���x.�5xR��p��5k�%�q�04F"ȵ��l4o*ȵk�Z��<�4���(9?6#j��iU�ظ����5�u�e��6E9��84���0m��J-6�vZ��G$5�5�3յ�6䴇 �5�2r�E"��c5X�?���5�U�5,�.��d�
�¶^>g5U!����5�����5��H���\6蛴5 ���Y�#�TI 4��u��861�6P49��#?6��46�y'6�g�5Y�6���y�G6��r���i�S!��?� ����6��_�P�b4��5ntѵ0Ŵ����b.�4��44���5.؋���C6%l5>�5�'����z>�����JE86Ȓ�5<���'�862��z�5��y5��ŵ4�-�B���}5�z�4Pޙ��5p�W6���tؠ6��7�ح�
��5�	յ~M6d�5��͵�E�6z󔶾��5Bh-5�I�6R��3Ћ.5�/~�U�6S�n�2�7��[�ƶ ӑ�(�!��Ĺ����ت6���6�':3�:Z��45g�6VQ6U��6���)97]�4��-� )D��f�5JCr���d7��7�ʹ6� ���p5���6O�l7z����4�#���G5���P�$6�ـ�������նqF��C��iE7Ƃ6�3� u��岭6ue��A�ж�:�5��7�v@��F��`j��)��m6B�]6�Y5Դ~�KF�5��
��6�X��ٵ6�����6?����8���w�4j@���ݵ��5X�����'�������@t�60ܱ��o3���{��8���	����f�5�N\5���6Z^�n�ж�Y;3�/T�켷�0!���'�4�c4�!'�+O��6�"���6��O6)��5�#���V6 �ֲH��4�獵��<�,5��5�� ����\��5�a;6Ŧ96i�=�`�D3�Cf6\}+���6ͳ�6�\S�lٵ�ܛ3�#�5$�j5R���EG��������dݒ6*{�5��α-�5�ő��@�5j�hO��"ڃ���p6��µ���+A$��5#6��ε*�j�Y����5`��>��D�z?\5~�5p�ث��U4!�5S�51ː6J.O�j�66á(6@N��o��5 4�톶��6�����^h���@7��5 �x�u|E�,�?6�@��VCZ��ez��aζY:�pK�:ܵ{k�66�9��K���B�>���+0��0R���X��ư���
62�6,_ɵ���8q}����k�E5�C�6TĊ6�U57�]���/6aI*�ԝ�4�u�4��_5�m6�\h6D�?���B6U47Rl����5���|������4ݬ�X-]��V��0~�4)�z56��6�a6ppH1�K+6I7�Ь5+S����V�5d^r��� E%6�6k��!$6���4h���&�����������25�b5���5Q�h5���6��������
�7� �?�*��5��6�76�[����h���5|!3601N5�d�4�˴0 6򭅵����5t�6 "������ҵ�jQ6�H����5��\��'�@�Ά�5������5���6|\��$���6���^�5���J����4��{޴(��x�5�ؽ�`����;b6Aεh���9勴���4||鵀 3��A95�0�5Y0]6��=�}|4m���ġ6�4tx.�l��5\�PO6�I6I̸�@����o��36|��6"Q@6�z����q�{ߕ6�������wJ6z�5��ݵ�2Q6�k�ț�qѵ��5
��5���6�4(I�P8�5�[��D�6'/�5�Щ�����X�4�t6��U5���5�����#6B�6�6bi�5Qڃ60�J����
 5i�K�x=*5��ĵ�����l6ƥ6���h��0ZT4Cv&��Q�6vrٵ(���6�)�����6��B���Y6���Fv�������Zε�b^�v!q5��6(��4)M�P�B�`u<��_�5TxY�E���ضs����I6.VE6�5�WJ���K6J�6P�Ŵ��n���jض��_�jd*�Zڵ	j��$�	6d��d ��ы6r=6��6��6 V94����
 $6̎��n�ض�	����m�6(�ܴSwk���6��6��ƵE�����6�B��u�c�ؙ*��פ5ѹ6g����wQ6�w�����5 �'�@��5@�_4��\��s� �L3��Ե���L�VH���t6�9�����5>���IW6&�_6�ƫ6>���N�x%Y6\=ݵ�w�6%�G6�����a6|��5�^���5
���6@]�6a�6@�G3$9�5_�961� �kfc5��\6���6��6<�y6���j6���3�홶��J���7�L�5N�� �^4ί�5�f�6={��Z1�f&g6x�@5�Bݵv�6���5��6����������6�R6���Ҷ�@�n����b(�����=�6�yζJ���=��r�/6�6�N����5P� ���6�`�5�/E�Ԙ�R`o6j�Ƶ�^����5�l���16���6��}��**��bC� ���6��5���6`�K����6ެ/�����5�76�	u6��0L����6��V6�݄5 Y5M�N�D6t�O�p�K04�L�5<�2�b�
��!�5�������6Ψ4��6��L��< �5��6�j��� v�~�6f7�.���Lɵ�Ԓ�a�6Zҍ����Lc�6�6��4�庵�f�6`X`�6�׶��6�Ӽ5wc96�����o 4jzF6���2�/6h- ��[�5-𢶔Z��c�3FR�]N7�35��/��J�6���5�x��Q?55`��C��^o���O6@�z6 �p6��3����5���Ѝ���W�Za���ώ��n5�;6@7���z��6�G@5v�d6�ӵ^L�5�8�4�G��}���D�5��6���6v��`y'��'���3��@7�'���/��66��
�T�6Ѷ3��|�ΰ6Q.���P�6ģ"��2v6��5�	6F�_�?�@6��>6��u6`��5�5<-�6ѣ�?}6�;5���6�%��Zgҵt��6p#A4�b16�_0�>�6���52��6`ދ���h�H%�6���ۥ�m����������#*@6M�>���[6n[����L6TJ3�Iu�6���4'&��BZ6���`:6 I9�D㿵�X49r�,�l��oϵ��"6$����ԍ5����p��Y6�3�P�����ĶP��4hꉴ� ������X���\�;<6�)��5���54xG���V��$�6 ��3��6�,��U��%6��!��$�6�����M5 �n3 I2��H5:�H6�)6E6�5�[�6������ҍ�6���  ���I��^�pz´Vd����<�5��P6@<�4��4$Ƣ6kqW66�����Y6Dql��L�5 d̶�g3�
��6ek:6,�R5�5P���lE6^ݴ@R��BTY5�����6vn���;�&p6̕����f��6���^%R����5�����5���0�5�K��:8c6�C�@\3��ݿ�JCg��-�5��G��	v6LԲ����5lR74Q��Z������r�5z�6]�v66�L6_!��`�5l�m��Nϵ�'��"��5��ض��,�@u6*��>���lh-�am�5����ݲ6� i�.�4�6"��6,����>�����5�Lh6�M?��M���b۵�4^6���5�Զ�.������X��4�57��x5�R��*�����5h�P���4��c6�:�sd6f��B;��޺5�S|6?EV5��"�v�\5@�γ��)6_t��/��x�g�h�M6 �����6��6>�L5 #e����6����s�,��u�����(4�Vѵ�zZ6�d�5V+�����6��Y⇵l���	o5X�=5�u�5�~,�6�(���6��E5�ԅ��Z4zr���ö���a��z�q6uw�4"?+6fNc6��6��6 83 ���>���Yw���͵�l6(�$��L6�/1��?	6���5&�ᶴ��5GY���"��f�6 �Z�R�5�t5X�A�@�5�Z�5\} 6��J��Ww6<(����6~׌6�'���Ϯ�sB6�j���w672�� �	6ҭ5��|R;�<\�����̟6���5�7l���G�5�� �
��ض����_h5�j.4�
���b��pvγ�Bε;6<�+5X�������0�O��05̲6B޸�j�B�(����52�5�9������56�`�5�h4���6JQ6[�6at���d�5(�� !�5�v���?�� 6���B!�H��4��[�|a6P��4�=p5^�.6}��o�׵��R4��U6�� ��w��ͱn6�#�+�N��wT6
���r=6�ζ�Iɶ��&�(�u��07�h���0XN6[^���N��5*�6�~�\6�	55�ӥ6 +��;q���Ъ���6�P�6���N�7�� ���tC�5/�l6�&G4i5�q�6�P�t��5���6~���4ʵw_.6b�3�K��6(�-��҄7���P�J�	X6%�|6b���������4�`�3e\k�@���6�\W7J���Ԝ�������6$A�t����Ӷ�A�6U!k7�;�����t�����6�]�6<��7�:��n���D��Hb�d{6���v�%��f6
�޶�9�6�O�L`&4�6]5B����O6���L�6�ڄ6��/4�7j�����lQ���[O6��5���6h��6̨K64���P7�^6��5�H
��r͵ÞZ6,ҟ��>�6������6���6mc3�r��y݁6��<���6�����N���+Q�26��h���	7���6�5�T��訶��6�U#�m��6�Uc�����t�5�
�6sg�6N^��@����e4�ώ���@5&)�5&����6x�6476M͵��.�v�'�/9�s����� 69i�6�U�5�?��5�w�66�I62o��o�6�ߴ��A���6�n6�ꕶ\p7,���,�'��6���k�6 w{�1j5^ݑ6E��6��J6�pֳ��ﶞ@�Tr����6.R��Qkg6�q	��I&��j6P�����48�}� ��5�ˬ����D��6d��5��W����6j)�6tz����6`��5��=6�6�艵&T6.5�6���64v����<6�)�6%�@�6ī� ��5����:)6�*7�"p6��7��05,0��P�6�=�����6��<6�s�[����sY5���5���6�f�6Pw4���1�~�w6B(�6�{X4|��5U��6+����޸�!� �����E�b6�6���@�3��m5��!6,~<5TA�����5<�69Aj��2����W��骴>�b66��5�{�5���� ���:XֵOJ�5��J6
�:!�hs�5���j��5e-6�_5��.6n5B��z�ߵ$�05�C˵B@�4,�5l�|��z��,��0&ŵ�iA��H&64���7H6 �i2�G�k�3��6�5�Xa�4n7h���5���?B��>'85N��5���5R���P�6���69�5��@�����c5�6~�	6٣��d��6�?i5P0 3�|(6/�l����-G���_6v*U6?v�w��t�5��j4��6Fі5e}��{�5�{o6�L��5�5��5��6�b�5�.��"	6��ܳ!���6�����KZ5��4&�����
6��3�Yj5���6���5����4�˿ʵ��N���@6˧���5�y�5��k5�嗶80S��45�V�5˼e5��P��4�����5����A^�L�'6�YE��66@qb�F��u�S6QϢ��#)�L^$��]4�f4aw6>�Z�,��4�]�4��V���ۘ6�t���I�s�5v䈶,nv���6�96$<޵�~5�h�L|�5�]<6ٷ�5��75�0���<w6�!�4��T6�^p�7���E	�6v 6�3���\5Y��5���6:Ӧ��Q5�۴4$�^)�5�<�5�We6�-��j��6r���<h7�i�5��76 ��l����4K����3��ҒE6F��5���60.��dZ�����b5�Ķj����ѵ��`��](5�<�:��� f6�pѵ0���%6(�W���Yb14����t�:�����-P� ���.���]V5;����5.ĵ�����96|4��r�_6|cg�x)r��Z45��߶�8��;z>�x���+��h�4:	�.@6�}��+���(5 ���[C�5��w�֚�5狈5 D]��E?5�C�5�����,d6�u95 ��4�K!�ȝG���>���4�'��L�a��X޵�����4U��5uյh�ǳ�W�4B���8�}X6�5�50��5i��5v�F6+��$5 ����+���x ��5�4Tm�5f4�5H]���+N6�P!6 �13�5�^��V򀵶���le5�G �[<���l��4���p$��(��B6,��=x6��	���g�6���X"6^Xw�9�K��M}5θ\���p��ˋ5�F��X�5đ�4�>�I����5=�6%�Y�`0���a��+M��?��<6����5��<��5���T47�0��d� �/�]�k�6�����~��6����4�p��xe5�.�Q�5�����6\�66���3(�&�y����D�������|��6���8�(�w��6L��xI�`� �ǧ:6��C����5+ڵrc6�_6p��3@����m6����끴�������4�fA6p]E6�`�5�ˠ6�.�5N),5�	�5��36^r!5_B5	͖�8)-��i����4/N��7�5�V+5#"����5�˯5ؐ���5��C4$���3�5 ��5��q���;6�2�5J��4T�4x_��,.4����j�5�㢵��5�o�������5@�ŵ��5�-5�l6���$��Z��6����з����Z����5�Q]5S\�5J�%5�/�����9o�5���6Xi�1���6*3����g�6��a�`�,4�c�p��� �5�*�������66��51cH6��/5���6���5�3�l�4诗4`�5h�D5 ��� a�3g�W6�Ƅ�s<�5�K�4��k��z�@�6��5֤06^�E6�+6��t4q�o5���5�!\�d`F5�/Y��5�|)���z5 Qh�yɃ6�,�ذ5f*-�d��4�/��)��JL��.���T��4d@�5�*��P6�ys�0�5Z�5"䠴�̯��ք�4%~5�ƃ����4�s�3��%6H>60m`�|`5h�s5��\�6�S�t��54n�5~Ǒ��0���ڵ�S嵚t�5k
�6愦��dx6�k��j����j
��X׵�_�6�@�� T�tE�6k)�5��6��(D��7�26J�I6��6���5��$6H6~���N5N������3D`6�@��;�6��;612��8�5s��7��46��5�+}6�St��pr6`���渶��5|��5|�4�*7��)�ye6z�6��d��45�E����6�oi6Pw����5�kI��s�ii6�{
���4��L6�O 6���j��56�#7����g��;hp�"�6�N�����6W,��u�6[8�6>M�6y˔�65Un��I�5i�6�V'�n$]6h�4� �GM66��\4pyʶln6�ٶ\���
���!��(s65.�6��&6ǌ���2`5��h6�5�>ߵ��B��
�TR/5���4u�a�k�׵@ζM3�6G�-	4�=���P�4rH5�Y
��p�����6g��61��6��t�嵪Fc6&%�5�s����5�*4p�b���a�M�N6=]�6'A6��P�����E6`ص,5�@�3x*�5 ��2NEF5�5f6^��+y�r�6u�|�*��V���a�s�6���5H
[6$T6��ൄ|Q�[l�5�rB�ҁG��6��k���5`ɳ���5A�0��ĵ��6�i;6*0ȵTO��
�붑�W����6 �3��7:���<6n�ݵb�"6L�5�j�4�A���R5��;6��6T05�鹶h�ڴm���6�y��(4���6���4lL	��s�6fa46S3=��J#5�ɶ����0ζ�[&��1��?$϶�&��J��X��4�m�5	��f�6hX�4
=���M5�+:�`�ԶL�5�u�`u@�8���"j� e
6��6>\��e�3�FeL�n�6�z��ȗ&6�.6I�5t�	�&���PM6����ƫ�&��736�S#��C˴l:6%Q��p�	����5G�yf��l5�q����6�����i6ج�5jb���Fp5rn�6�εF��@!2���59�N���f��)$6�"��Ğ�����!��T7��5Lk��w�4 C�6n����'5���6OK��7a�Ȅ�#���ܗ�8�5�5s�66��,��~W���3 6�:6,#��|6�u5ya 6�X+6 ��4`�BnR��~�+����2 ��.��H�P<5,�I5=�)6��������P�6�J��%��6��ɶ�H��<��0�K4���4�x�������)��k����y5�ۺ��7�"K��T���v޶J�����6�B���a�6�
7�����׶Yа�aۼ6 �6�K�҅���K�"/u6��I�ƣ���x 6��9��6��K6Ϋ#�d`����ɵ��5�ʬ��7�4��(5�6|#�5\:�����5�/���@��P7�(�4�O���6$�y6ݽ�7�6CJ5����L&�6V=��f�W�d��6��5�@� v����60W/���68�E�f�G�RJ%6	.��⑶��u���5xY5��4dLJ��e��k�ѵW��<�7 �����'6��&6ܴ��<�K64-�5��f��rK6�c�6%���d�v�q5/5-��Pq$6YF6��Q5V���S�5�gW5��ٵ�c6���5;;+6O�6YU6�=��F��N�R�p5Ԙ�@�5׻�6���6�:6���5�t��a�6�Ď��Ҵ &�"���mL?6�p�4��iaH6K9��r�6��ڵ�YV6��r�ֵ��7Mw3�����|�6`�8����5 v6ZZ6���4�O6�1��}�5�Hص@}�4�D�5��*�����y{6I��6�ZP�D?�6�6��Gө66�<���7�*֔�P;�5����4e��25�f|����5�b5��T%�Ԝ=6�4U5͌5V�D��uk�x�5r:>�"A��r��"l5��Ƕ�-6Oh鶂�ߵ�/6d6���6U�@��5qy�8?մ5��2@�H>-����yy��δ�t�5�ٵ�xD5�>S����2ȮY5���5����� �� �L6@�a�|�B5\�Z5�Q6�g 5�}����`��£��9�6
���4P4z}���6Փ6�M*5�ص����޴��x��$�5�6�F�45��56dY��}Z4���5�f�5���4w?[���(5�+���5��}5v�5�I��%e"���M6�/j�y6,� 5�.��g�5��6|��S�5�;4��5�u.�`.��珵�<5+!6���4Z15N4u� [{��(�5�����:���\5A����=�4��5�쬵t�_4 �#3 ��K�������5|��6h�5�&95��7���75�Y�4��4�r>5���5�"��i�ܮ+6�'�5���4E�5A�5S�5n����V�Ȫ�5��v��Vֵ�ƣ5�ﲵ"\S���4&��5��3Rē6G�=���������#��T+�NE���^�5�6\
��&� N�h��4H��=�5�ɕ��ؓ�ؘ���6���5%�ߵ�Q0�q�/6�3赯���f9��������3�5� J5��i�l��5���ڟ�5�;�5L��4r]6rY���V۵p�F6�n�4Xx���.�e�ʵ�5ps5�Q�Kc16LX����5!���k���ȴxn�3~���m�����'�6RMϵ��P4���d8�6�1�`a6 �k�İ����4�BC�\ӧ�D�����3�Xp8501ͳćT�p����64q��$��i�{�j��n���95�	���F3���1i�G��5@��*�LϷ5��5� B�F��1]�4���>��4`�5��R5dV�R��5B�w����5�I�5���&?U�vm]5r/84XӴ%�L5&��{>x�R��-���ԕ��zR\5X5x�<�-�,��m�5����V8����N[��P)5=
��?�@6���5��D�P�5�k�?�����N���5	5PK4�;� �  � PK                       checkpoint/data/17FB ZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�b�3�|h3���3�f3�`�3�I3[�Z3�-3��3[3�O�3T��3�F4�q3��3{t^3�s�3��t3�3�"3���3���3ل�2$3N�I3xa�3{3�q4Z�g3�pR3��3��3E�3�ۏ3ŗ�3�J31�3�4�J�3]P�3N>�3v��3��A3��r3WƵ3�Â3W�[3d��3'7�3FF�3�YM3�3P��3�t13J�|3:L3�E�3�}s3Z��3 �3�V93N�3.�(4���3�y3��2;t�32��3�3S3�43�+�3jr�38IU3a��3k,�3�_3j�23/�4<?h3&93D`�3�R�3~�S3�L�3�_�3{�.3�yV3���3P՛3��*3��3�_�3��3�|�3���3_9<3�Ǳ3`�p3�y�3�G?3 �u3n
3��3A��34��3PwT3�BI3K�c3?x�3&�3TI;3�Ќ3NQ�3b��3|��3}��2��3�SD3y�c3�5�3�!J3�3��3ۿ�3�#�39�H3)d3C�4�i3���3��s3Z�3�c�3V�C3�<3�R83t��3ͽ)4N��3Ɯ�3��03���3Y�i3�ѧ3��3��3�h�3���3LB�3�X}3�h<3�l3U��3VL�3c4���3�<�3��=3�i�3�k�33�3Ъ�3>/�3ۏ3|3��u3�k�3)m3��z3�T�3��\3��3|X83`��3e.N3�3�9Z3��3b�3�N�3�b�3Khc3��k3-��3ȓ�35C23���3>��3�p3�L"3m�q3���3��:3��3u��3���2Yf~3M4{3���3�R�3�K35E�3��"4�l�3�@d3�N3�x3=L3�]�3\�3�3��41R�3��3)[3�0O3�D�3o|�3��3���3ISa3we�3�
�35 �3Nc3�w+3��&3�	=4�S!3hud3K��3RV�3Zen3@<3cT�3��u3d�3Bd4t?�3y�}3�C3$�4`ވ3d�!3�
�3��B3�va3���3b��3/W{3n?3�3�6�3f��2��3os�2�3�˙2��3c�E3�b3 �2(�3�Y83�,3[+3���3�g&3��2��2� 3b�K332�2��4303n93���2	�}3A�3Z]:3��3�s!3��,3�3��%3X�2���2M�$3F~93��B30�2r�>3ٌ%3�]3ُ�2Ĉ3��3g��2��3�+3^�E3"�<3�S 4+Y83�=3�D3��,3�O3eY�2�34�&3�G3�4�3�r�3_q33Zg20[t3˄A3~��2Z��26�Q3�p_3L��2{"3��3�3�R�2�J�3���2C3n#3J>T3��3�;.3u��2���2!��2΀+3�(m3t6�2s(q2h�
3�oR3B��2�`3�9�2��3@�3=\3��3=�3�23[�w3h3�3��2�o3��3}��2C�3�&�2?�3�x3]
3H	D3w��2��3��3&�2�u"3 ��2��3��:3��3�fB3�3�3-|�3�o3+/3�d�2L�N3�2#Ze3��'3�7�2PE*3��3��3?)>3Z�3��*3��<3Y��2E� 3���2o� 3�b�2x�e3��3sE3IR�2�R�3��2�3r��2Gö2�3��330m3�ف2�k3���3c��3ķ	3��2��3ٴ3U{3*�83w�2�S83]�3f�K3�3�]H3�]+3M�3JV�2�P3�39�3�3��3+3Ɩ3�3xZ�3~��3
�2ӏ3�<32��2�D3w�L3���2�d3�y3:[�3�1�2X#3�m3�=�3�0o3�qa3;�834�43��3[E3��=3Gk�2�n3F�g38�3�T3V#�2�"3��	3�63!k3d�2i�F3|��2°\3�63?� 3s�2y1�3�l�2�a3G�Z3h2<3R3�	3
X3�2�M�2�u3>��3��U3쏮2�`:3q	3���2ʄz3;:�2�}i3-�83� 3AJL3��I3��l3w�3\n3 ϐ3�c3��3�63$�3�u�3֘�3[d/3�}�3��3�x�3@�+3?cu3I�53�C!34a�3{�X3x�^3���3ܿK3иr3��@3��c3M�4˨63-�w3О]3��3�B�3�V�3�3
%G3J�3�3�39�3&�3��3�3@�3I�#3�$�37�|3#?�3��q3%��31u�3)`3L�3�=4�(@3F�3��3h�35�3])�3��3�3�͡3���3�-�3Z[�3��3X�>3�Y�3w�3akF3k]3�ؖ3��,3EF�3�x�3l�f3b3��74��A3>�R3�$�34Â3��3��~3��3��3���3�@�3���3���3��&3=ag3.��3*�w3��Y3�e]3꩷3�/3V]�3�33��Z3U@)3!�.4�e-3�!3v�a3(:3-ca3	}3F��3�d3#r3]��3e"�3jS3I�?3TT�3Y�+3��73 N�3��2�M3�c3�٫3?�K3&2�3�u�3kn�33��3��G3��53Yv3���3E�v3	H3���2���3P�4j�3���3�d3,�3%�l3B�3���3~3��i3nEF3�tY3��v3\�3��3�C4��33��3��&3�bk3|4S3؏3�3_�j3�CH3��4F1�3�D3a�3��3B͓3��h3��3&�2-��3�Z3<�3u�3�#�2�@.3�Q4�]U3�r3�z�3��3�p3��G3S��3xrM3r�>3�Jq3��4-,3�[3ڊ�3�VG3�Ke3�23�83�IZ3�\13f��3��&3)��3�3p3��4�~)3�5�3�/r3�a3���2�Ra3��3Q3���3���3+W�3�s�3B�*3u��3��3/%y3z�j3�3��3C(T3�x37�r3��/37�>3�*4��j3L#�3k"�3�=3��Q3��W3Sn�3�H�2�3�"4
��3��3'b23[j3l��3C�W3G�3�<]3_�3�;h3�-4O.)3�^�3h��3 �48�3Q��3�3+��3B�3��N33� 3Zb34җ3AG3���3��3sb�3>m3�13��!3�G.34
�3��2�F�3�e3�o�32�:3)��3��3d1�3!�P3K��3B913C�3���3�d3AͿ3B��3��3�#3�34��3X�3{A%3�=G3y4]3|lQ3�L3�>�3�Fs3I��30�3	^4ժ03��\3��3�H�3�V3���3��3�t�3�q�3��3���3�I13׌3�ć3O�3�VH3!Lt3_f3/�3Xl3��3Vg�3$4��P3�4#��3}�3���3�6M3��3�~�31�3Ǚ;3��3�64�`�3��N3��3�>�3��C3�J3ᮬ3�13FV�3a|03��3�CN3��G3>��3�@�3<,�3��3A�3��^3�Ȏ3 �3g��3��3�r�3�3%��3��3�?3]�3�Ψ3?ds3���3-�>3ɜ3�"3:&f3N��3M�i3�3�94�YK3, i3 ˡ35��3ɐ-3�ʉ3�_3�*3G�b3߂�3l'�3���3�@)3v�4u��3a�3Ō�3�Q3�)�3��y35]�303
�x3��3+��3"=B3"dS3;>.3��H3��S3޵�3���3ڇ3$G�3�.�3q�3�]g3ne�3��33� 3�3C]O3'^R3|!c34{�!3o�q3O%�3>7�3@z>3b�D3��E3�ɑ3��3L|30��3��3���3�p�3��3N�Q3#$3�0�3+X�3\�R3�ӳ3z9 3�s�3^P}3��3�qE39T*3"7�3���3R�3�#�3C�3�ך3Q��3o�53��3Uq3�n3�04ᑾ3�Ԋ3B��2��;3�5�3�Og3CQn3�v�3HՐ3��63�4f�&31Y&3y�\3��4�/@3��3�37<�3D�3�a3<3�f3�@4���3@�3{#�3���20�3��l3�d3Z/33���2�=�3B��3��4�q�3M��3��3�Ӿ36�S3.�i3�:3�3M�c3�{3��|3��03λ3U��3D5�3��P3]�.3
��3^�h3GK$3��3��3�˿3��132)�3��m3Y�73�@�3��3`/3 
n3�N�3v�83I38�D3�WZ3hDF3�(�3c��3�қ3ߙj3�@3��{3?L3-4T3�^e3�+m3�r3oS3��3�n237�3��3��4�υ3%��3���3�q�36��3Pp�3�[3M�3��O3��24m�s392K3v�3H��3��C3�
)35��3.n�3qC3�� 3��3�Ox3�+3�S3>V�3!3�e3�^\3��s3k�3M�3��3��3d)�3u{�3�ux3M�}3� 32`�3{W4�Z3��F37>304�3��63 �3��/3�z3P3~}�3E|3�� 3 p@3%|3^�G3��3�9�3�B3��3�3��3��3�%�3	��3v�l34�i3�џ3�k3@�3���3�JB3��i3��^3jRJ3�4|8I3|�3�34}z3��e3�3�3f33�.3{�37#�3(�}3��A3���3᪆3�x3��t3�738�3ɩ3o�3dN3���3��	3	�3R3+Y�3Du3�GD3�� 3Ѫ13���3�-�2�?�33�3�|33��3T��2K�3:0*3n&?3'�3�_3�i�31:3x�3�ym3:�3Et13�H(4O�33|�73�S`3�:)3v�13%WZ3�c3��3��3�mk3.��3�{�3���2���3�u=3��3��3�w
3��43�d3��l3�b?3�q�3�^!3��3��t3pB3^�f3�(E3��s3��E3Ϧ�3#h3ED�3R��3��3��q3}3��3�
Z3�p�3��3E�@3���3�5(3,��3��:3�4�3��2��4�?3���3z��3b�3���2��}3
��3ת3� �3��3��H3Y4N3�!3o2�3b283��2���2k@ 3(`3�/3��4�4]3^w�3љ3���3(3�hn3MeJ3&�d3��43�q�3��3{B3��3��4��t3S;3K�3���3ք�3�2�s�2	 <3�Ӡ3�c3���3�O3�T~3�5�3'��3�h=3�C3��436�3ɼ<3/��3D��3и�230L3~��32�`3\�3�3a��3�z3��)3a�S3�9$3�P3
�t3&��3s�3X�/3��G3���3
N3`��20�c3i,E3-[�3cԎ3�@�3�j`3�g33�ݮ3��S3�R�2��3��3jX3��v3�3�^3��3!��3�s3��+3\�)3:�3�%33��3�?3�.F3��3�ڃ3(�V3e3O�=3�5�3�N�32�A3 w3pqy3��3�s43x�j3��93�f3�Y3M�23�b3���3�@3
�3g�3��L3aV;3�
3/�3z�~3���3C/Z3��3�ۤ3�:�3��L3��b3��3h��3�?93�ʒ3)ZU3�j]3��E3x��3w�3��23�Zv3�w4-�13c�3�Z3�^d3�q�2�ܑ3Bf43�3YUc3���3<�3��u3"#�2u�s3�3��3)�3ɶ 3Q�V3ۿ�3A��3�B3k�@3�*3Ū3�*3��\3�?:3�(+3�)=3�l�3�%�3��b3sv�3Q�3���3��K3��3o�(3�:3 cG3v9�3}YL3�[3�R]3�ˎ3�UT3֦3�3G� 4(�2��@3��(3��P3�G3S!3��3���2;P3��35I�3�W3u�2�B�31ψ3P��2���3�3�;3I�M3U��3��23v�H3$+3���3�p�3sΆ3��3��3&+x3t�43�1,3�E�2�O3�D�3�a�3T
�3(8�2��3l�r3�r�3�`3?T�2(#B3w�3��%3d3E3��2�4�3�3\!E3�h^3��3�/3(_�3 �3|��21�83B�3@*�3��3�Q	3��3�b�3�93��T3���2s8�3���2-3�C�3�M43R`4՟�3~��3V��3N�3�/3��39k�3$/3<��3r��3���3��^30�;3^�4�a}3%�33���3d�3(�3<73�3�3��v3�|X31:j3���3x�3e*r3T�d3��A3,��3�3���3���3��3Mʇ3��3��63z��3A~[3Z�q3�c3=�3
h�3�6|3���3Y��3{�3�'3�u�3<�	4&3Yh�3O�j3� p3�?�3=��3�ܰ3)~83݄i3v�4���3�6�3�u�2�uq3=_�3Q�>3lЮ3��@3��3ֽu3��3OU3��O37A3?74�J3��]3�Y�3�/�3�Qk3�Ͳ3���3\hW3#^�3qR4;�3�?~3��3��3%��3��3��>3�N3Z��3�" 3�H�3|N3D�U3��^3p4��3�-q3LӜ3��36 �3^>�3��e31�M3i��3BY�3Q�3u?3��53}��3}��3O�23���3:�)3��3x�13A��3�ܓ3{�3�<631I�3p�c3��r3�c3g�3�mF3}^�3���3��A3�0n3m��3��3K[�3�B;3��3�	R3�:3:(Q3�W3o3ʙh3��X3Dgz3(>3��=3��U4�[=3uw#3��3�532Z�3+"�3��3 4A3�h�3�=�3};�3O�3�.3�.�3�R3��3e`b3ËP3��3v�W3v�3ø�3�D3#�h3:u�3}�3q��3Ac3d�3|@q3�3�>�3�q3dZ�3cJ4u�4��93���2��3�]V3��>3�"�3J�.3]�3l�3�b�3Ӌ3^ i3�3x�X4��A3�13R'�3}��3�A�3^x3���3�	3�i�3�ٳ3AK�3�x63	�\3*Z�38�Y3�.(3�$a3��;3�Ú3�Y3�>�3\�>3RX�3��g3=�04��r3%د3.�3�`�3e[O3���3M��36e
3�+4 �4E�3i�3=�3�_t3^�R3-�O3[��3xk3�<�3��^3Q��3^��3B��3Г3^P�3���3��v3���3v��3��3%ѝ3d�3d�X3T�3�P�3���3$��3mh{3���3�6�3m@%3�]39�3P�`3�3Y��3��3Gp�3��_3�4"_[3��3�&3�	�3T��3O�j3hڷ3�9S3wW3v?�3}�Y3�ݏ3�i3qv�39�j3�!3�OQ3/^i3���3�b3n�	4at�3�x3a/�3�1�3*�3���33V]3p�3z)(3�3F3 �31I3%tb3�4��3րb3x�3��x3� 4�g3���3p[�3�E�3��3M|�3��B3��;3��F3��4{`3�k3~R3���31��3�3i3Q��3��2wA3���3'9�3�N�3u�3�F{3r@P3i��3�3ِj3���3�a�3E3Vmr3m}3lt�3�e�3�33cN�3Å;3ϗ3}�13�Bl3_�s3�3��W3w��3iC4n9R3ȆN32_4?Fw3崈3�3ߥ3�K�3dCP3�H�3��-3-�}3��'3�P4/ъ3]kZ3C.X3�V3.vK3=�A3Vf�3�A3^I�3���3O�39�3p 3��3Fª3g238�W3�3��X3l3ұ!4�P3iTq3J��3y�D4�os3��3[�T3�X�3"�(3���3��K32^3�u3!EI4�ߠ3��.3u�3�3et3��U3��w3
[�2��z3{gL3��3~30�3�h�3T4f@A3BV,3��K3��=3r�f3|n73�.�3�3��3���3��3yk]3�_�2n3�u[3I2S3���3p�3˳�3r)3��3}ن3�=3#(�3�!H4Oi@3�MH3�K`3a�p3i�C3��3XТ3�SQ3T{�3 r�3��g3BТ3��3ݫH3�s31F�3���32�2?��3���2Y6~3W?n3��73��2*��3�(,3�r=3�˦3#'3w�3�~3��3�D�2Ԑc3��3�s3�W3�&36��3��2۶�2n��3v�/3�E3�I3�3�3���31��3#Ws3��3��d3<��3D\�3��3$�3�z�3��3{�i3��f3v�3�T3;��3^u\3�r�3��3 &3��3Ec�3�%3�V3�r�3��3�Ձ3N��3� 4L�h3�-�3�э3�r�3QY3葎3�e3���3��g3f�4㭟3[Ӻ3�S:3T�Z3ʔ�3Q�53��3&�3���3��s3�W�3�.�3�+�3�?3~��3�P�3H��33P�39�30��3���3&]�3<�%3$�}3�Y4�_3��3�e�3���3��3=�\3�3���2˂3���3���3��3�g3C�3!=4'g�3�$3��3L��3I.3��3�;�3l-3[��3���3J�3���3�F3�r�3��3 d37� 4ҨS3��3j�3-��34�3P�e3	��3ҍ4�S�3�fD3�?f3C��3Ծ�3>�3ӟ�3` o3Ȗ3r��3�{�3�ŗ3��S3˫�3��3%k3��L3�`D3q3��j3���3&
}3�d3� �3S~G4/�a3q#�3�H�3�/�3��3�B�3Ұ�3O�"3��3!��3�B�3t��3�B3��4��3�N43��333��3�C�3pb�3|�$3��3�(3�4yA3�ɒ3&!V3�;3���3I��3�Ds3ے�3�<{3���3iġ3���3��!3���3�Ɇ3�>q33�3ƇJ3"Q�3�V�3��3Az3>��3��3-~4(�f3Qe3ߍ3P��3�3��35��3�u3ş�3�>4�3|�~3��I3+��3qv�3-��3�U�3��L3��3��a3G��3�P�3��-3F�3��*41��39�3KQ�3ƨ�3��3��v3�"�3��3�Ć3��3b��3���3v��2�=�3蒶3�n�3��3�u3�*�3:�H3ݺ3[2�3;�%3c93��G48�y3���3��s3�r�3ҟ*3��3D��3J�^3���3���3٤�3oz�3��3p~3
h3��53�z3�=3ے3�I13�� 4�-�3�[F3@	3&��3޸m3ڊA3�A�3)^3sA�2K433K�#3�3�uG3���3�;4u��3ޜ3��3T,3�q23��3���2TUI3_F3w~i3��43J�*3ה3�z�3��3E�3��*3��k3Z3!΃3�J53V�2��i3�f�3�0�3�-3ߦ3�S�3]�Q3`3:�`3��3��3k3�)z3<y93yK3p�3e��3��p3i803�39F3]��2I��2L2<32��2��3_�3�Rq3��3<�/3I�3�9�2 �38�63%��2K3Z�28�3�s3�3�΍3)��3��?3"/�3��x3�n>3}:W3U�3���3�1�2yv�3%��3�N~3��f3Z��2�m3tw�353��a3�,�2�փ3o�2�ئ36�3��63Ȭ?3U1�3��W3�"*3|Hr3�P3��>3�x3�3"�3�?3d��3���37%3�3�֔37�935
3*��3=�63��;3
�3�D�3���2 �3� �2q�3`A53v%�3K=�3:�<3'��2v3�2L�3l�13_\R3"7�3*C3�730
E3�B*3�Ex3��2QW/3^34L3�3z�3f��2w�37�2&m�3r��3Us:3��I3~3��2�k36IZ34W3�
�3y�3��.3�)S3��3�Ҫ3��3>�2�=w3T�=3��2n�#3h�3�=�3W3�f3|G�3gZ�2�e+31�93څ�2��W3P�)3,��3nO3>-[3ܸ3	�X3�*~3?ܮ2ټ+3D��3��2s��3�=�2�V�2]"h3�f3�'^3Ʒ�2�"�2��	46mZ3N�3���3ƇG3�4 38�3]>[3Ra�2�N13M.+3I�p37ߘ3H�3nC3sH�3�Yo3�sN3lx�2^<�3�-�3Z�:3?��3M��2X��2Һ3��2�w'3��3�0�2p3��3̆A3�"�2��.3rT�3���3���2���2��Q3��P36G�2�&3�-�2)�53�v!3�Y3�3�J�3"�3z4Zy3��3��V3���3�y�3@��3kIc3zE�3+�s3�v�3�J4���3- �3�3���363 ^3o�3�,�3��a3�4�҉3mE�3Hc�3ټ
4m��3�ݎ3� �35�4�a�3̐�3�I�3�g38o�3L��3TG4\@�34��3؛3��3���32�3�G�3ˏ�3-y�3�X4�q�3l�4��l3�D�3L�3�׏3v�3��q3,Xv3z�!4��3g�]3.��3؂49�3�k�3���3��3�!�3d3��3	a3��3�`3�[�3D\t3�3���3�6L4*#3�|�3[�3�{R3�e�3"ڤ3�3�3u��3�I�3��+4X�Z3�+4���2]�3ȋ�3"�=3љ3��3�۾3�0�3��H4�͈3�G�3L�3�Y�3�ϣ3.p�3UH}3v�Q3l�R3���3��3ee3o��3H4 x�3`z�3;�3�P�3��3'G3֋3�T3Z'�3Z�3!��3��3�3�3�o�3#`�3C�3xC�3Д�3 �~3�c�3k��3F�3��{3�'4Gi�3
�}3}�P3��4�G�3qT�3ho3"3M��3��3z��3.�3I�3�~�374���3{!46��3,��3Pa�3���3�J�3ӣ�3�@�3�o4k��3�s�3�i�3�J�3A�3��[3���3:[3��3f�2ʧ3��3O��3�M3�Z#4W4�3�K�3���3�1�3�l�33ʔ�3`�83�q�3[�4js'4�J�3bo3 ��3�z�3�m3�D�34B3ym�3Md�3��3܆3	ɖ3)�V3i14*)83b�e3٧�3Ny�3 �3�b;3���3�5�3s�4Nkb4�1�3j��3��2��3��3��n3���3�dS3���3Г�3f4�3��|3�I�3�A4]+w3 �3u��3"x3�\36�3�Y�33��3�C�3��4��3�b4v�<3��3��a3��3SN4��y3�W�3��3��3+��3�|4$�h3��3+co3<3�T�3�I�3g�h3�Xr3~r�3��V3n�f3�"4�}3��3�F�3Ø;3<��3�x3[�z3�
�3n�4&�93���3I��3�i�3��3���36A�3}]�3��3$��3.�3���3�׷3o�3�$4d� 4IB�3Ύ�3 O�3�=�3[�3c��3,�3��3�Q�3�^3��H4���37��3m3l��3��r3=R�3�s3ș3�.�3�H�3��3�l�3ّ�3r�3-��3T��3�?3%ِ3�_�3�	u3#�3��3���3kM3|�3��j3
�3���3��4�b{3��3�I�3}ҁ3=��3�H�3��
4!�?3�\49�3�J�3�֌3Fol3GV�3�W�3	χ3��i33r3|�'4e�Y3%o4B �3E3��=3N�4ϋ,3�%�3�Hb3���3�v3Da�3�3��*3[��3���3�2�3I��3S�3"�3�T�3KfV3t��3���3O�3� �3�=&43�i3Z�73��i3��%4�Ԯ3i��3�Է3���3���3gt�3���3o3Ï3>�!4���3�a3m��2���3�Ѷ3�p�3��]3(
V3�G�3^k3ˮ3��3��03o Q3�d84A�3�x�3��x3�Gg3���3�4�Ԋ3�c3��3cn�3��3�,�3<�^3" �3?73�3��3���36��3錖3�[�3���3�Hq3��M3���3$�63���3�|3u��38H�3�~�3��3�D�39l�3$z4�]4��3��v3M_�3�3\�3���3�3��3+��3��44g73�_3�{3�`,4돷3���3'�3���3���3�oA39Ѱ3W�]3>��3�^�3!4���3#�3�V3�O%4���3k��3�/3{��3͌G3���3�e�3�.~3�=�3��'4�ˣ3�P4��37�13{.m3ɀ�3��3^�*3���3��3N:�3�X�3K�39��3,��3Z�U3pb3�P.3{V�3B)�3G��3�ƍ3��g3CHN3���3	� 3��e3M�!34�3���2�3w8>3��a3�?3P޺3a�3 �:3�:W3$l4��43w��2h�[32r3K�"3!�+3ϕ�3�V�3ЂY3?��3�/�3�/3�93��_3((34e<3��*3�rQ3E	3U�2��`3�`�3��+3�(3�v�3"�u3d !3� �2��B3��^3��u3Y��3(Ձ3�!p3��3Q��3=1(3�S3��3��M3:�2b�73Ҭ�3�{3��3T��3,z3��53��3�!�3��37�3fi�3�c93���3�@3Ү3s_$3�!3\k@3�-4�O33\�3�Md3� 3��N3�Dd37J&3��3tۢ3�7�3#�]3�H�2(��3tt3t%3��^3g�3�\3R�2̻�3V!3�a3 3���3�<3m�+3�P
3���3�G#3���3X{33��3�r�3rN#3�3��)3{��3x"3�+*3�p30��2�R3��3�U3
3B��3o�3��3�3��P3/t�3k)43ǻ3�[j3�3��2��g3)��3��3ɏ3�b 3s�t3���3��2y�3%��2��S3�|.3l3�39�3K 3�l�3��3�F
3(�2�6*3G3#At3��23iv�2?�@3�g�3$��3�3ܖ3�3m�L3��3�ƃ3��2�pV3`�3�p3f��2�zC31�%3��4T;�3�+�2��3P��2�=3yE3���3o�)3��3�6�3���3-d23�l�2��3�3�L�2��3�N�25�\343���31}#3��H3'1�3�t�3; 3;�2�3�3�B�2�B>3�L3d6!3OxR3u�3��3��/3R]3h�%33glN3�a3���2�Ԕ3Xv
3�i�3��3��
3�k!3�&4��W3�yt3��"3�3��2ujb3j�g353�X}3=�3 �3|K 3tZ�2��b3�6!3=�31<@3���2;p3UU�2�Ұ38�3oCo3���2#IR3�_�28E3��3593�O�23.	3���2V(3K(3-�<3h&3Cv�3���2d83Ru�2�239��2��43���2E�3��%3d�2&o"3��3�83B�2g3��2�v3�]�2��3��.3�,3�Q3�_�2���20�2m�2L�3�]3�:�2 �2�� 3�ǲ2�	3`3�-3oF3��3B!�2� :3T�
3��
3|��2�"93>O:3��[3�k�2�T33<3��2{�3
�y3^EB3�23+3��F3�_ 3i�2Y3$z�2��63�>3 J�3�ԧ2֫3�r	3vh�2'�	3�)3XXd3���2���2�3;�=3k��2���2��3r�%3��3��3!&�2ה,3_��2�I3y��2dZ�2�
3><�3��2�Z�2;�3�!3_T�2В'3J�?3�L�2:c3��y3��3M�Y3ȕ�2��_3c$@3P��2,3�
�2��3�3��3��/3�>3�t�2�֖3�\83��83��2� 3D333�.,3��27A�2�T�3�X:3�i 3�}�2D��3�*3�#3}�%3}��25�a3&��2M�3U��2��3ki�2O#�3��3��3���2�o3�
3j3�q3M��2���2O��3R�n3C53��2��3���2w\�2+�{3��2�@.3�f�20SO3��3�;�2O��2�3��3ǡ3�	3�3��3��2�63s{�2�~>3��33P�q3WA#3���2�"3�38��2��3t|3��3p��2*He3o3��3s��2|��3��&3�D-3pv33k�"3�|3�3l73���2��!3o�I3c�-3��	3��2�:T3��"3"P�2{�3��3de.3���2P�E3J�3pH�2q+o2���3�l�2�s3#3�s3�J�2'm�2�M3t��2+�K3�`3�_3�V|3��2�63K��2��2���2���2	(3�F"3�?3��#3�K�3��j3��:4�U�3��3%Ԑ3���3p��3���3��3��d3Qov3[p�3��3#��3$]3痬3B\�3h]-3�p�3[�3�4}3��.3E`�3Iƽ3N	R3�a3��3���3\ S3vJ3�53,D3+��3d��3��`3W�q3�݌3E�3�ذ3;q3�}�3�E3��3�53��)3� u3�H3b��3!p3��,3e9�3g�3⢖3��63���3fe�3�_�3�R�3Ÿ�3w�_3�@3�Ni3�-�32�M3F/"33ƻ3��3f%$3L�3e�Z3ڭ�3��c3�Kx3$�H3���3� �3�h 4"[3�'\3mz�3�(r3��3J��3y��3.�3���3�!4Vع3`-3iH3�$E3\3�z�3��Z3y�w3ӝ}3E��3���3Q�3g�?3��R3AX4��B3ԞI3nM3��I3L�3�8P3�
�3j�53?��3��3{�[3�4�3�3l�d3b�03h�3b�Z3|_3�zN3�B3ν41{U3��b3H8�3�44!�93�A�3�S�38�u3m��3�]�3��3���2t�d3�-�3���3�l�3�t�3d�4fY�3�s3�T�3��3���3r�W3�{�3�T�3
�83��2�m�3aKi3K͐3j�.3r�l3��b3���3��B3���3�ն3J��3��35��3{593{��3��3��H3���3:$13��w3��x3b-�3��3կ�3�fT3ߕV4��J3 �3�?�3y�3�33Qg�3.\c3ڬr3�ތ3�t�3_Ҽ3f̀3�=3��3�:�3��=3㔞3>״3��3��)32ծ3SZ34��3�l33�v 4�g3��R3o��3*��3�L<3�ǅ3:p3i�]3aC3D��3I�3�*n3��43y2m3�o�3G^�3�x3F�f3D��3��3���3��_3�pX35D3]4��3f{3(��3��3�(73��N3d��3�q34��3=�.4" �3A�{3��2�~�3�83�3��3:��2ʊ}3��3.q�3�ug3,
3+�"3���3�7l3��3��3!��3��>3-j�3"sa32#3�S^33�3��3�T|3Ѕ-3�|3,s�2��3-�83RX3=5(3�3�M�3ݍ3�ݝ3MMi3�f�3�WP3,�q3D��3"�3��3��A3a&�3��L3�c�3���3���3w�N3`F3��_3 �n3��w3R3{X�3���3�pA3뱧3�D3�P3~t�3$�4<<�3�o�3#p,3R�K3ZnR3f�63��3��;3V̒3�3�3K4�3h./3V�,3v�3:39W3g33U��2��3�73���3^/R3c:�3� J3��3�,U3��'3	@3S/�3ޕ'3�H3C�W3<3v/N3o;�3L+/3�r3�'&3׎�3)]�3� 3|83;D�2 �3��,3���3:��2q'\3��2-��3��`3��3B"3�G3�r
3me33C�c3�3�'3RLf3�lh3��b3�O.3���3��31��2��q3��3�l3}t�2j��3�� 3���3�~43�|�3�r�2%9�3���3ک>3q4�3>�r3��@3��c3��73*��3�Ww3b�3���2�X|3���2��2ӕ�3���2?vI3�S03��]3�!$3�
D3��3S�3�}U3�҈3}��3�f3��
3�aY3�j03C33���3�&�30��3�G3\43���3H3Qs3R`3>��2j��3s��3V�31�D3�h43�03�@4H�i3��N3*`3��3ݏ53�s%3��B3�+3�y3�l3]��3�*3`�2��3�#3�3K��3n��2ᮎ3�1k3�i�3�J3>L>3�zG3��3�V3޶3�Q�3�3#3��*3"�T3���3>�3ي3��31	�3'I\3�>�2�Sz3��L3ч3;5V3s�&3�@3�z�2ܤ/3ZD]3KB�2�	3ҷ�3�%D3~�#3�G3N�N33��3ȼ3S$�2X�3[ґ3J��3�Z63��2a��3I(g3��3�>@3��2&�3ۧ�2���3��2q�4�^\3���3�yN3�n�3p�3L��3���2Zѭ3�f�3R��3��n3Bl�3���3�wa3Ii3�p�3)q�3��38l^3WӘ3c�3CQ3e"4� �3tn�3�!�3�Z>4@�3�<�3YK�3ɭ�3'�3˟�3d8"4�)O3�7�3:4!4��4�]�3j�3���3!��3}r�3���3283W��3@~m3� �3�om3Wb�3��3�S4�e-3�\.3��z3���3���3t�3��3���3�ި3�H$4
��3}�S3�3��3U�34j�3
�3��3a�35�U3��3�+�3,��3��3��A4�QT3x9|3)�3>}.34	U37��3��3�6!3]3X&\4Yڙ3*�*3؎I3�G�3rX�3W63ȼ�3�3���3`/]3��3��3?��3���3�4���3匱3�X�3R#�3V�3���3��3��3}��3��4�۪3{_�3��3��3��3�k�3!�3Hh�3���32-03���3���3�,�3Fp�31��3Y�A3��3+�3�D�33֓3�ñ3��3�ّ3�P|3��I4�p4�I�3��x3�K4�ŭ3�cZ3V`�3�Mz30��3�zG3sN�3��3�P�3�\3�R.4�tA3��R3�s�3�N�3�+j3h��3�Ӹ3(�c3zj�3��3Ÿ�3��3C�13N#�3⑘3,[�3��3�'/38=�3�po3��3��H3!��3��d3�ii4�Rr3�Ў3i��3D�~3���3�$�3��3�iY37y�3W� 4�u�32K�3�`r379�3d��3m|j3�3�sp3:�4ʾ�3�T4b��3!C�3D;�3��I4S7�3�K�3st�3�s�3(�3}T�33�3<�3���3�X	4T�3���3�i�3Bu�3B]�3�j3��3p��3x�3lߤ31m4���3y�:3��3�r+4��}3���3+4��3�3�C�3�G�3g�Z3Cq�36�3��4";"4�v3#3۫�3���3a��3f�3�\4��|3N��3��4���3':N3�?�3��)32��2��3tI3�3�$3nه3�3� 3�X3���3#͎3w>3�	73+E3H&�2��2���2�iG3@�3}�p3��S3�3�!T3���3tN3�&3f�`3@t3lA3'�
3Ӱ03�/�2lA63��3��3B@,3��3`Z[34�w3Ǥ836�3Ū�2���3VJ�2��3E3p�3�\�2��3�s\3'z3�&3���3[�3�?�2c,3y)�2``3u>�3p^3��?3� 3�A-3�Ck3�73ǭ)3R�3sy	3L��2+�Y3�dA3!��3i�U3���3��3��3��53x�a3�h�2��3Y�3��2dOK3���3���3�>�2��
3\`n3Mj3�3�+3�.3YqL3�Q<341~3��,3�3,�3-,�3�v3�PR3��J3�a3��2SVl3;�3,�3�3��3�|�3E3���2���3��e3�t3�S3I�23�QQ3��3�3%3J��2���2��3ε 3��r36VS3N��3�Q3E�)3�(>3��2�J3h�3&�3���2�21.3S��3��#3��3�}3��n3�P+35qD3�A3kE?3붜2���3�RE3��3<3�3�C33�b3�T3��43A�E3��3!V�3�3XG�2�5�3�m3$%3N�3�2�)�3��$34ʝ3�^03$�3��832�3,[3�(3�t3��3���2b�L3��3B�2��+3��3�&=3�X3�!'3,93xr�3� �2*�l3%�03;�s3�t3/BP3�	Y3��L3x%=3�64 
93��3�O3O�.38�3�k\3�Ն3U�3�Z3l43!.Y3��[3���2R;J3�Ѓ3�-W3vk3�3_W3���2<_�31�33z�2���2��3\�2)�(3A��2�3o��2T�63Z:�3��3023H'�3Ϗ�3�,31��2+�i3�3��2��93p�3���3�^�2d��3�K 3v|03�3�t�3��M3M73Z�13��g3ϐ�2��3�23\H3��(3f�3�m3
�3^3�Q�3<[3�. 3�H�3�ܔ3�lJ3��2��3�w3~)3a�e3_�3�3E�36�l3�E�3�C3J�@3�3x�H3��#3��a3�{�3�М3�Q3��B3/o 3�2#3��3�3c)3q�G3�W�3��~3��T3� #3k��3�13t�b3�83�ˍ3�3�W.3=Ds37U3��Q3�.�3E�33�.3�Ա2r��3��3�9�2�>M3�O33'�3��)3$6�3J��2C�z3�]�3��4=3MN3r�&3�c�2�?3[�q3�{3�L3j�3��3�^�3�#T3h�2Xެ3rp13�1�2U+3C�!3.��3
�#3ڀV3g�"3lE.3�13;*4��2��^3j=O3�y3�J30�z3�g3MA)3�#A3w�3��B3Z�3��3�Z�3E�3�2'��3�;3�=3A�3��t334A3.9&3�ո3=_�3��@3�~d32�37eI3�93��3*��2.p�3ޓy3 I�3���3�3���3�b�3��M3��3��j3�}�36�2\"3�.m3u#3�
�3�,4Pv�2���3Ʋ3;k3��3CI3��]3Z�3]�X3q%p3��3��O3��.3���3�Bq3ll*3�[j3�&3�Č3+`q3��3xtk3(�03ju�2��3-�/3�"@3��3�3�3��k3�3Q3��2FO3��l3�b�3��3�� 3�:�3�8Z3;�3w[n30�'3�rQ3�<3v��3~�g3��;31�:3@�3ᴕ3<�@3c3>�m3��/3A;$3-)g34�2�5D3���3�0�3�p3�=�2d�i3���34X38
F3���2Ų�3���25�3�/�3�y3N��2��4n�13�N3>�3'3�!3�,I3�`3�M3�Q�3��F3�	4��^3�2�~�3��G3*��2��?3�H3�e3��3�n3�n�2U��3(3���3���2��3�,(3V33�3�U3ڳ-3�,�2B�3;/_3�\3*s30�3�`�3��p3���2�}93և3b�Y3�>�2hn3�m3
|3nrH3��3��2;KK3q��2�q3*13�t3�<�3( 3t3I�33�.53��|3t9b3�q*3�(3>3�3-3_2;3s`Y3�$D3Y�G3���3�ˑ3�3�`m3%�
3�3"�3N
�3�35*3�3M��2W��3d�3�k53�) 3�2�2)�23zV3WѲ2j�O3̲F3�=36K�2�i�3��2��3_3
04d�3#43{]3�RE3�| 3Fq33�C3ˈ"3ƧO34�3s9<3��63��2��[3�:,3c~!3��]3�v3���3ɇ�2�37�=3�z28�3��3�V�2�,�2��M3G��2�%S36�?36s�3���2=3��c3�S@3C��2�s�26��3�=3]A�2�?3=l>3���2��2��3A�3�lj3z�:3���3t�Y3��]3#>�3U$3��3OЌ3Q3��P3�U3g��3Iݵ3��'3g4<3z��3�`D3I�38�X3?�,3 zn3e�<3�Í3i?U3�K3�ME3�2�3��#3��o3>Rs3��3�C
3�O3@t#3��O3-�3�4�?3K�3��2߄3�A{3Z53��t3�N
3�<3�|
3T�3--!3��u3�U&3�B�3Ř73���3��m3��63�>y3��_3�l93�I3j�\3�8{3�{~3yq83��3pck3��(3KA3?��3��3Y�o3�e3*�3]=&3=� 30p$3>4��S3�<E3��H3��O3��.3�3W�O3\$3��2{7c3��3�Qi3��	3z3+"h3
Jg3@A3�`�2��3O}#3bmm3��I3�3��2��3T�V3��V3)Y�3��3`�3v C3�_23��3��L3�Ȃ3���3ls3�L�2u�I3�l3�`3��z3���2/Ig3�� 3��x3�G3$�3�3��4�_�3���3t��3R׸3#�3�<�3�l�3q�e3���3/�H4��3]m�3�o�39��3�
�3�M3v�3���3g��3P�W3�.4t��3��u3�7]3:MF4{��3�	�3��3}ś3�!�3J@�3&Y�3N�3��3j�4[=4�Q�3W`�3	 �3d7�3}�3��3lR�3���3�(Z3��4��}3D��3��H33��3���3V�3
%X3��{3�3Ǚ�3�s�3�_�3|��3�ݎ4J�3KM�33oH3���3���3�C3���3�2�3���3��3q�45B�3�N�3��3G|`4Z&�3�I�3�n#4+�3���3]��3VY�3�£3��3�4;��3&�3��*3� 4��3�ڄ3��
4���3Lo�3ND�3���3KR�3M�3L�^3T��3�m38N�3ԟ�3�r3HH�3*H�3�@�3�9�3vO�3�>�3&R�3���3!_b3]
�3��3�ʖ3�P�3d�|3�.�3N�3RX4��4���3 M�3[=,4F�34q�3h��3xة3N�3�<�3c�3K�W3��3*��3=�3�i�3L�Y3���3���3��3�Z�3���3:�3hg�3:~�3b��3/�m3�Ψ3��4��4L�3>>�3�T�3욓3w.`3���3
�3�3l�4�44���3D C3�C�3Fp�3��y30X�3>3�i�3@�M3_��3��^3���32��3brj4���3���38��3��[3�\[3<.�3�K4��)3��3.�3�p�3��3�=�3�:�3;W�3lѢ3�$�3�\83D��3�9�3kI�3��3fR�3ؗ=3n�4��3H��3!�~3�r3?�w3fO�3���3��s3I74�94>?�39�3�M3I��3���3��3���3ahi3C�4�P�3+�4�/�3=�J3� J36x>4�D�3�v�3���3��3�ʣ3��u3"��3��A3�`�3]y�3574ݓ�3�T3z�3,��3��3���3��2/�4N>e3�*�3<��3o1�3�/H3�^�3�\�2*s�3��{3���3}և3˿r3��3�'�3KX_3�4U2�3W�p3�'I3�Ƞ3��i3��2�~_3Ð�2z�3�UT3�Ϲ3Mr33I~3K,G3e~4؆93�p�3��P3Pt3��v3���3���3/*�3S�3ua�3�6�3J��3��2X�3�\p3��3 ՚3f-�2�+b3^�E3�CR3�l3)r�3r>73�4\U3E�f3��%3Q�z3�M3��w37��3�6�2' g3�0�3�t�3��c3���2� g3ɮD3x��2Ǟ\3\@3�[�3�X3dz\3��_3_��3��]38�
4e+R3���3��Y39�2��P3�"f3AX3�.3y#23��4U��3i_3�<3/��3�EW3��3n�13�e�2(��3Ț�2*��3�3��w3��3��3�	3�{33܋3`S!3S�t3�m�3�{�3�A�3[I�3���31��3�53�3���3]̉3>+3���3��A3aIg3iX3���3(Fm3�}�3+3�)�3�3�gI3�u3��a3��3xak3[�3ds 3���3�3e�3d�3��=3�Ω3�1�3�3��93�]$3Y{3�v3�N�3��'3��[3a��2p�
4�_3��3u�!3�kl3�~,3�J3y�}3�"�2"�q3]�4d��3ͨ�3#�3l�3R�3�3S�3�*�2���3st�3��3�L34W-3pß3�4�U3��3�Q�3l]y3
D3�f3��s3��U3No3`\�3y�3$_�3�3Zi�3��3��3
�3�!3��3���3cS�3�.3@(63v��3l*4ܭ�3��i3���39L3���3�N�2PR�3��33p�3��#3/��3'�3�|3��O3y�3.B3Pf�2
s
3xlk3F�3�+�3PH�3�L3�a	3�614��"3G�m3�c,3�Ȉ3�4=3*�3��z3z� 3�߀3�?�3��3~�3�;�2�3{ڪ3�s3tV�32�F3<	f3��!32#�37҅3Bٙ3�J38��3r�3��/3���26X3R43E�m3kW3Դ3��l3M��3+1�32�3�3�ܥ3��3�3�25�M3+3�]W3��3��3�Kg3��b3�xF3
W3SV]3�K3Q�3���3�w�27H3<h3�1[3�C3O��3�ۼ3�G3R��2�I�3��U3�3�3ދ83�o;3��X3|h�3:i3u3fQ�3c��3���2WYQ3`[3��w3�$3�9U3�M�3���2y�e3J�3ʉ�3�C�23fC3�&&3`��2%E3�A3��63�lp3#JH3&I83�a3"�33k�3%+3Գ=3�Nb3��2K�M3�9�2Ͼf3Q�2�PK3@I�3�N�3�n3m��2"�^3�W3C�X3Vi�3�3���3�}+33zo3hpN3�}$3��.3��3�V3_<E3673[�3�f3��>3��3he3�Ch3h<`3|[3}j23�#3I��3�'3	�,3��3��2h�w31�3�׊3��?3G93��<3�,	4�S3�/�3�Nf3��:3�r�2��3J��3���2��[3jZ�3�Ȇ3we363�&�3Dby3�K3�u3l�#3r��3I�3P�i3�L3X�V3=ן3�4�3q�J3���2}e$3G�`36�A3�c�3��3�6�2��3���3Q�Q3�B 3��c3��3�gp3h3���2kͶ3�$3UT�3dB3�?3:<W3�3z��2#�%3�A3�:31�3�m3LiI3�2�2"HB3-�3�3P�3p�2�u33��@3� 3�}�3��28�3�J03�G�3�\3,��3`*c3��4��33��V3�gw3��3�$3��J3:Y34�73��3��3�Yn3Ǣ3�R307�3��3���3'@L3��h3��13��Q3�e�3U�-3�d<30N
3�D�3�B3�=3q��2��/3Q��2�3�[3�A/3:{3���3�o4��y3���28�K3X{3�@3+�|3RR�2֣3��)3!�3;d53/�L3�3��3�k�25�2�H�2�@�2��g2x�'3��3;b�2*��2��3���2��3<�3�*K3ݒ�2x��2�$�2��2F�2 �2���3F��2�� 3��2��_3�V�2LMD3��3"}�22��2*w�2��l3�3��3҂�3�L03�R$3��2��63�� 3H��2!נ2��2���2�<�2�{3s@3��b3��2���3+C�2<3��2�X�2���2
�2��3.��2G�3i|3a�3U�2�ZZ2��3���2�8�2qa�2�B�2��W3�B�2C�03X&Z3&�3�D38C�3���2���2��2-D�2�U32^��2"3݀3[n;3YHP3�`$3���2s��2��3���2�^�2nd�2.��2�3��3C�	3���2uZ�2�|�2@+3�n�2�,�2���2���2�ʁ2�3��2ck�2k�3.?�3�73 ��2�W�2�R3���2��22.�2���2;��2Q�2�	M3���2P��2'�3���3{��2��)3�3Gt3*��24�3�T3�3ּ�2���3~?�3>��2f��2��y3{E@3�f3+zB3��2ЄD3��*3oE-3%ڈ2^,�2JE�2AԮ3OU3��2 ��2���2��3M�@3BM3��2�63���3���2�2u��2ؤJ3�� 36u�2]�3j�2j�3ڻ�2�b3Y�3|2/3���2d��3��3%��2b/3A3���2:
3�M,3�Ѵ2�	�2�sT3nh3Z�+3q'�29*3&��2��2<P3�F�2��!3PP3�(3~��25.3���2u�c3O�2{�3B�\3CM 3e&�2+E�3H�83W�.3�0�2���3K3Fm�3ý�2��3��'3�>3M�"3ι�2h�3�{z2'�o36�3A��2`�2��N37U�2h23v$
3aQ	3� 33�8+3@�G3�2�3�*3��O3��2P'�2*�N3[�2R�3��3���2(z3]�3E�S3�k<3��3��%3�C�3�ٖ3"׆3a[3[K�3�?3�Ԃ3?g�3��&3	k3���3�,�3/�3�0�3x&�3I]�3�pC3�&3��3%q3�;�2h�3P8�3�e�3ĕ*3�O�3ɝ�3�@3I��3{6�3q3U@�3�ym3P� 3��n3��3R��3+�3&�2)�3WL3�Q3#�n3�>3=!�33�&�3�J3��\3,{A3�W�37�3���3TeB3J3q�3���36a3��3���3݁�3�`�3+�383�{�3�3�13V�3���3I�37��3�"V3N�Z3��3�{3�l4I�&3�a]3�Ǚ3t3Ɥ3֢3xy�3��3�G3���3B}�3F0i3L��2�c�3{�f3j�%3��?31�P3-=�3��)3��3�$�3��3��03�}4+oQ3H݂3��3�p3��J3��3�=�3��b3��3-
�3��3p�[3K+3k^i3�,3Ö3���3�s3*�3I��3�>�3읙3s�#3ea3C4��K3]$�3��3B��3�13g?�3���3�N
3�rm3X��3�X3-��3%�3�ƌ3���3%S�2��3�
S3���3B3A(D3��s3�r�3�H3��3��.3q��3N
3.�'3�ݍ3��3��3�y3���3C��3��f3�D3߬�3H��3�!H3�l3���3��w3�'�3�5K3w;�3V��3#�=3\ʃ3#�4���2��S3o}_3�(=3�)3r�k3��/3��3[�~3�w�3T÷3��_3?@�2%��3�3�r;38�3��3�+e3s'�3�t�3��3�C3���2h��3h�>3���3DU�3��@3�E[3��3�:u3y�B3Y�3�d�3�){3�ų3��3��93��3�n83a^3��E3��3=h3���3�	-3��2aI+3�@�38'3實3I�3_�Z3>�r3q�3^Q3+/3��3���3�A�3��3��3�Dg3�ӄ3��%3�T�3�[+3~P�3js�3 �H3�/�3�`3K�2`_3��2�38�3�3���2�:3�f{3٣�2v�2��3+�23�v3��L3xZ3��34��2e��2���2�;�3M��2F�:3J�G3��L3�>3�<�3w3���3M�a3~$3��X3x�w3���3U�K3��U391G3��t3��z3�-3�{�3*)3r�3��3�>3�c�3a��3�.3���3H8G3oh�2f��3��3t693�203,4+3�_�2K�;3BQ,3�Y�2��I3Y��3��k3��3@9�2L
�3�nd3��3�Z3S��2 3��2҃�3�%�2�	A3�4��3<�3�[�3>�3��2uِ3Q��3���3k�j3�G039�3-�3�F�2y�3�@�3��3�23�3V38e�3ܨa3�]3��<3�O23��[34�3�ڣ3��2�o3ܢ>3X�3�j3A�3��o31xh3��=30��35/t3��D3�93{04}J323�G3�3�/73\X3�?73Pu>3V��2�� 3$G�3��3��$3��N3�3��I3�nR3�;3�Z3[�`3��3q��3��3$:37�Q3E�e3O��2��m3�^3�3'c*3)��3Ձ3���3�
:3��4O 03+͟3��43�t3_��2��>3�H�3���2ʯ�3YOM3�ʴ3��`3�>�20r	3EJ3�Z83�a-3�:�2���3��3���3t�S3m+3�%3���3�m:38\�2I4�3:8�2��63��3�˛3�L�2�F�3]U�3X5^3��H3J�2;�U3�H3N��2g7x3�?�2��)3XwF3b{�3��-3� �2>�43��4�m3�Y3�539�35;3\�3W�&3`�3��H3	R3�S3?�73�`�2O�&3���3�=3��e3|�2(ѻ3�3�8v303�-30�2��32�3�)3�/93h3��3�o3��i3�#3��+3'�3&C3�;3f�2��%3\�3zs�2!��3Zg�2�3o�3���3���2�	�3˔Y3eEc4X��3�404W�&4��4��3W��3:�3H��3�.�3$kM4]�@4644�Or3L�4��54>g�3O��3O��3���3#�3�A%43��3�c�3�^�3��X4�A�3+n�3�7�3��3yw�3�L�3y,�3��3�ڳ3=$B49J4�&$4G!�3_�	4���3���3_�4�t�3)9$4�t�3kh4 �4�
�3�b�3_z�4T?�3?��3j��3V��3��3Q�3���3-�3_��3UeI4_�3�^�3�#3��3��3��3qe�3���3�4��3W��3���3��3"K�3f٭4T�3��\3l��3	4E$3���3N*4h`3~�4��3�3>�/4\\3�=�3�:94m�13�Q4��3,w4�u3u4�3�Mh3��l3^�P43�f�3 ��3���3a4s�B4X��3���3��3Q,4�L4��3-�X3�X!4���3��3/J4/~�3ޒ�3D�(45�64���3f�3�Ñ3�Wz4<��3�3�m4s9h4�s4�}4��3Ѻ�3g�3��I4�{4���3��3��4rh�3*��3�'"4j8�3~V�3�� 4ȿ>4�$�3�k�3 �r3S�4>R�3��3O�4!=�3�04�l�3T74�3M\4JT.4�$94@��3 �I3���3z'�3�ҿ3��3;�T3��4�h(4z�4/54���3�ے3��y4�h3�N3XfZ3J��3~�3�L4%�4�<3�6�3Q�94���3$�3,!�3���3�Y�3p��3cO]4#x[3*i4i��3��3���3Ϭ�3@��3e�q4�4M�a3ļ.4k��3�s�3N�3&^�3u[@3�4�_4�:4�4�Y�34�3b�4|ç3���3+�3.f42I�3E�+4��4�ߎ32��3���4~�3�N�3���3H5V3�7�39ry3c�3�3��3��
4�4$��3�LP3N��3���3��3뚱3�*3�/�3�@3�4/ҙ3� 4��3�o4�1�3u4��l3n�3U�+3+S3s�3��3쥯3��4m��3%��3�Ǣ3ԓH4�}�3S�3�ζ3x�3�]4C�A3aI'4��3/�3�f�3��"4�o�3���3�c3��3Z��3���3�*4�Q3�_�3Pm4>:�3��3'��3���3-<�3� �3]4o�_3�y�3B1�3�|�3�â3Ђ�3��3�4.��3 ��3���3�;�3��3z
�3�/�3D&�3dɗ3ox�3`֭3�n�3<�j3\��3�|�3�&�3�d4NF3ò4��3�^4�H�3DC�3��3�ˆ4-j�3�@�3+~�3�B�3o�e3%~3�^4s�p3%��3�04ai�3M��3���3�ʹ3���3P�t3T٨3Κ�3�m�3Yj3|?4��P3��/3���3��[4�z�3d��3b��3�>�3 i�3�3`��3�u)3cq�3�L�3H�44�4���3{�3��3�c�3�[�3�la3�y4�y�3���3���3B<�3Ү~3?�#4tϚ3d��3r��3M?�3�~3�?�3��3���3��j3��3ы4��3L,[3�&4���3�:r3{�3�D�30�4]H�3%q�3sü3���3Ff3��,4@ȁ3t��3Yː3Ԭ3��3G��3�'4��Y3Zu4Q4��04f�3�u3:�4N.�3$��3!�$4�;�3���3�8�3'4��3�p�3���3P�E4���3���3��3͇�3���3<��3�m�32�3Z�42F4 �
4���3�$G3�4�!�3�_�3��4Wz�3w�3��^3�6�3�9�3��]3��3- �4l�3F_�3*�3��3�3�i�3�π3��3��3ϒ�3�%:4r��3�33b�3��3o�3�ܦ3�+ 3�"�3W��3��	4��+3��
4B�3m�4؈{3���3�j�3�}3a�3*x�3 <4*�^3pk�3��3�94��3��@3�#[3���3o'3���3E��3$��3̑�3mҭ3��3���3R�3��4uH|36o�3�a�3f%�3�w[3T��3F�y3}o$3�3�4�3��3�߀3�t3 M�3�l�3J�<3�3e3�G3��3�3S�3I@�3$eN3+�%3v��3�P�3gas3^o�3���3�3iT3;r3a�!3o�Q3z6�3�y�3��3Q3�A�3���3\013�-|3�y�3Uh�3�j3��3es31[?3��W3 9�3CI�3�}�3IE&3h��3h��3%�93bK�3Ou43��93�r�3�f�3�W�3*�36��3���3�G83LG3i�3���3�j�3(�F36?3)#3fl
3s��3*�f3�,3��X3�Z83i��2�~q3�;�31�3�إ3��"4��3\353�u�2q1�3ڥ�3:i3�7/3H� 3��3< T3�п3��K3]��3d�(3�H42G3��3ԡ�3=m3$/t3�W�3�Ii3s.3��3Zַ3�ݚ3'j�3���2?�3��3}�3��3�73Yޟ3úB3"��3g�(3��U3��3���3�6S3~Z�3�d�3^�l30+�3縎34��3�AR3u�C3� �3B$�3p̩3�^3Vq�3��4�DL3�k3{��30��3�ï35y�3 �3+z&3*�<3��F4esB3�*`3��Q3���3(_(3a�3b`3�	�2�/W3Ĳ�3�=�37�V3�3�a93�&3d�U3�W�3���2��j3�#3�ׁ3���3B��3��3ȷ4f�v3+�o3�:�3�3�3�O3=��3�lC3�(r3oJ�3	��3�3�m-30}�3!b3�tp3Ĺ]3�N3�un3bVd3���3�<o3�Q3U6)3GR�3���3<��3{[�3V�2�YG3f;�3�d�3��x3tp�3h%4㯏3�Pu3�3-ܓ33~�3u��3��3c/3�h�3G13���3{C�37q(3��2��3��G3��n3ϐB3��3��24'�3��3p�C3x�u3��3�M�3O�T3P�3�,�3�03a	S3�g�3v�3��3|�3l8�3�v'3�$3��*3E#z3"3"{�2:�%3�I3<�d3��d3�xP3P��2�H3��3�H3��C3��3��|3:W3���2�m-3%<I33�R3��3��]37�2�L+3Uv3��3q��2�^3R+x3��3���2�53.�f3q��2�3�lv3�	�3�O53��2&,3�?>3�N3�{<3�3D093Y*
3���3�33m�3p]�2�ʵ3=\3�X3��3G3���2b�3��N3�3,S_3��3dV3MC3?�2U'83��H3_\�2�343�2?�@3h�3�3�x�2Zq3Wb3�i�3E�3�U3@m=3���2��3��53�t�3���2�d�2O��3��3��3�!�2v�b3�T3sE3 %.3��20 �3�Z3�*\3Z�Q3;'$36�73mN�39#H3J-3#r�2�03��3`=3��3z3�53p�3�<t3	0�2`3hV3�JK3��"3�3Y,�2�G3���2DƝ3$)3���2�3ĝy3N33�3�q�3�3)��2>�v3 |e3��3)6'3�͞3'r3��53�̒2i�,3��G3�j3�3�a�2���2?��2��G3�7E3�#3*;�2Ւ�3��93�0'3�93}�313�xT3��K3��R3gkI3��`3n�Q3��!3�>�2�n3P:3�(�2:7S35�3�83�[�2!wt3��"3|g�2^��2��3�m[3P�36�3XL�2���2A[3V�3sC�2�q3Š�3ȋ�3�3*��26-3V�h3��L3r�D3���2��`3R�3J�33?�2�h�2���2�n�3�+�3n�g3�4%34�p3��2L�q3� !3!��2'�@3��3x��3bS"33�291�2�yF3��2��O3���2��%3K�2�43i�2.�(3�)3.�4z�3;3 .3��3��2�r<3s33Q��2g�(3��3�ֆ3�w.3ɽ 3Q�%3<)93C�3�a3@��2��3`�2pYI3E�2i3��	3�TJ3��V3���3x|3�
d3�C3��13N�3��3�3@i`3�l�3�43��"3�N�3'�q3��/3D�<3!�3Zĕ3�k�2،3�ql3��k34At3�c�3��z3s!3A,b3�԰3�ݶ2
f3��K3iv3_&m3b�3��3�[v3=3V}3U53��2 ��2KN_3@4�31H3H�3q3:3��F3D�63B��3�x�2[093�d3=��3E�2D�3Lʜ3 Q�2��3��4؊3A�3`�2���3��13(2�2?wi3�r!3�@u36
#3�O3Hq3U�@3��(3�D4���2є
3+�e3GnL3��3�q3�X3�ʝ2"�Y3G��3�ދ3�$3��2�}P3�43|]3��3��"3���3�K�2:�z33EG43$*3OZ�3U�63�^13���2���2��!3�L3�-3<$�2�R3'V�3=�>3��"3&��2���3w�w3��3.�d3�� 3�z3�iF3��L34�=3�3Ywz3�y3IsE3�H+3��3b�V3�>3�%3&�g3�̷2��*3�?�31,�3\M3'��28l3��Z3x��2��B3�E$3�73{+3r��3��]3˨�3�53w�3��3��K3#� 3�o3x��34MY3�!3���2���3�K3o�?3��/3�xa3Ǵ;3�Ga3��63�03�30NO3���2 �3�<3��|3C��2��f3ƜG3��33�.�3��C3�z3sh+3vȱ3�}3��W3Fj3Ш�3i�*3z��2!��3�2��3#�u3�3�9a3��3�%=3��r3$�l3��2E
4�3�g�3L�W3y-3���2LQ3S�C3�_�2��3��3Zv�3�}�3�2�Gy3��j3��3@�3��33�t3���20��3T%"3P	�2|��2���3Ì3�53F͔3�O3�s#3�I3��O3���2��u3�@�3�Oe3�??3�i�2S�O3x�3�P389�3+�3�uZ3o( 3��3C&F3+��3.�3��3��_3�T�3-�F3;�3�Uo3^��31�m3-s83c�H3��3�S�3��3ߤg3�u�3��3�t&3S��3��3ɢ�3B�-3�V�3vYI3�VY3�kR3���3L3r�3�'4چ�3� �35Y�3Z�3h�3H֟3$��3���3�,�3PI3�g�3Mv	4. 3J�`3}�3���3���3�p�3b$R3�3�"3a��30�3�$\3b�3���3��D32��3r'�3�e3i�d3��4���3�'�3ZO3��W3/�3��j3��,3�ڰ3�&�3^W�3��3%V3�*�3�53 34�<�3y��3К�3�3��m3U&v3���3�Io3r��3\K'4�3y�%3�[3mY�3�a|3��:3il�3(#3�C�3]�+3:��3�y�3r�S34�k3���3�a�3JZ�3g~�3t+�3�6e3�g�3-ɩ3��*3(Ѷ3?4���3X�r3�9<3��4x 4xW^3�|�3,�]3�}�3G-J3$*�3 Q�3���3~��2�e�3�G�3�+|3k3�i�3��3D�3�}3���2a��3Q�4&-�3�b�3��3�?�39�3<%'33�3�gf3ދ�3ӑh3]a�3Q�Z3�w�3�"3�4�37��3߃�3��3S��3�W�3kF3_��3���3��%4���3QSE3��f3d��3sMd3��O3�p�3*�83g��3?�{3�$�3�ԑ3�vO3wVv3vU4c3�#@3Fp3�&�3;�j3�&�3�/�3�^I3��3�@�3<�3f�Y3`0E3>��3|��3��D3�ӣ3Q&30�f3['H3.�3��3䄍3��3s	B4�^�3|�3_��3��$3�6&3zX�3��3"f�3Ԋ�3���3#��3m�3ٕh3ku�3 ED3���3� �3�v>3���3e�3�b�3�UN3�l3���2�+�3ܤ
3�83�*�3�B]3|Df3���3���3�83ܦ�3�V�3j$�3Z
P3р'3�4�K3�hY3+��3�S<3���3�A3�Ӹ3s��3`31��3���3�[�3z``3�J3£�3��$3���37�3Ѹ34$�3���3BB�3��R3�>
3�w3���3fb�2?��2���3wB�3��3�u�3@s^3i�3�3��3�k3(;M3ڷ03��37�F3�93�~3�w&3u!\3).44�:3��3�2G��3��N3eI3Y�3�3r�3�]&3D��3��;3�3�A3a��3g�31�>3ZC�3_|t3��\3��.3���3%�3b�Z36:4U3R�J3W�2*�3��33x�[3I� 3�3�v3	�K3�,�3��{3Y�E3K>3B��3c�2��v3`qX38�W3�A�3�373M3�3�ӷ2Sp�3pE4�MB3K;F3+2
3re=3ĵT3��C3=��3	�3��3:�E3�3u�'3�jP3n�x34�;�2��}3H7{3�J3�ac3L��3�3F30)N3/�3D=�3�83��37�3J�3cv 3^HW3�Q�2�2�3�aa3	��3{<$3��<3��!3���3�N�3�zX3�fx3U�3І?3�3��3`~�2��-3B��3���3\{�3.W'3�^33%X3��3i�Q3Ĺ�2X߈3o�3j�h3�L43��d3]G33��31�:3ہX3 �w3��!3C~3��3�=W3�13��{3���3#=m3��@3v;3Cey3�Z 3�P~3�3�37,�2N�3x�Z3�8�3r�n3�Z3~C03�\�3dd3H38�23��_3�%I3�{3�3}3��\3�Ə3��4��3�σ3n�@3�&�3%9�3�G3�z�3|��3E�3;u�2�m4.�s3C�3Y3#�4zi_3��3��3h�3"[K3�Ck3��)3ft3���3d^3)��3^�3ڡ,3 �A3�]|3��03=Nf34�2&�t3̴e3R��3C�3��3�m23�t�3ik�2^�3^03�~N3��3�n3ٿp3 �2�	73�� 4��3wr�3��2��3�^�3A�3��=3�t230��3	��2��3p�3͗d39@3��3��&3�6�3�6�2&R3u@3�&�39�r3��3�o(3`�3�y3�%I3xJ,3��*3�"!3S��2��(3h7 3�a�3m�2�236�E3583�G3���3wR3^ǀ3V�2�$)3�)3�hj3Au3�Fg3h7p3�n3^�;3}�C3Qf�2FKA3NE03�~3r�K3~J3�_�3��2N]3��j3>_3J��2��3W35�(3�@F3�א3Y�2�L3�b�3���2�+!3��3��G3�װ2���2�M3��3�}�2��93c>3�>3hn�2�/83$��2��3�mF3�P�3313��T3N�3��3�`39�3��2JH�3�[�3KH�3�,3dݦ2L�3�q3G�3]��2T03��%3�#3c��3w�3Զ3T�3�W�34},3cH3;�3&J3�"3�_3K�3 83g�3oJT3�1�3t�;3��2h�G3��:3k��2A3��3إn3RZB3��3��f3��!3�]3)��3�`3��D3���2W�Z3&3��Y34�k3 ��2*3\Y�3׫d3�,3>�2��3��u3?�,3p��3I��2%k3���2�T[3��3:�Y3��3t��3�<H3��!3j�2�4�2Q�$30u83u@A3��3{�3(�3_�K3Y�31ߢ2��&3)�13_�,3�)3e|�2G�13�T3T�\3��3C�3Y��2	q�3��28�2U@63�3���2��J3�d3�~ 3{Da3�9�3l�o3�3̀�2!
X3�%3��27Op3��2��3�/3H�Q3�?E3(M3��3�]4�!3�3�!3c�3��2�`3>�m3993���2b�j3��+3y�3��2oT�3QK�3��3 3�h3�:3'p�2�93c,R3�%�2m��2�4�3
��2�43[��2��3M��2��E3qo=3��2�K3�؅3�Rv3�3KT�2;"u31H3�`�2��,32�2��G3�6�2,N�3��!3Թ@3�3� �3D�23��3���2oI�3�s2�>
3$�3c3���2�7u3f^%3�3��2�CL3�23r�2*3t�r3p�3��2���3�2@3"5�2�E=3�gN3�3�3�h"3V�3�J(3M�>3��X3�93=m3�ǐ3-ez3̩?3�e�2�[3�^�2��2~�;3�3��3Ȓ53k,W3ʪ'3PVc3��M3���3��o3��M3H�*3l�_3���2��R3:03�k3M\3��3��i3�)�2�Z�2��>3�iO3>��2�=3��X3��d3�3��3�u�2���2���2'L�3*��2�m3{3�2�83��2�h3"6\3���2���3�ױ3n��3�j23���2�D3y�|3W�2�HC3Et�2�9�2
�2!ǀ3��2��3�'G3� l3�b*3@3��@3��3�J3�<3�Ճ3�}�2�503T�3YI3�63k��29�O3�"3���2�3�33 �3���2�e3�B3IS3�+-3��3�3{�3	5�2l��2�%�2�	�2�3���2�03���39�3A�3ޞ@3CO3�BW3<R�2��3�R!3��3
:3p�3�� 3`2�23>�2���3M33Z43�NR3F_[33�2~ �3�׳3�*`2�3��x3��\3Xce3���2�(03��%3rx�2��k3,�2Ù�2�!�2���2�<@3HF3r[53�Ay3�2!��2�j3�	"3Ɣ�2���2]Z53f��2BNE3��3�t�3zW�3o�3��3c�%3{~�2�B3Sw�23�u3T>'3�+f3�i3��3e��2�:4���2�/3�qS35��2�k3dÈ2կS3�%3�JM3R��3/�33D߮2�3��l3U��3�pC3H�3_�3��24�3ls3�9�2�T�2*&�3�e�2��3�[�3��-3�G3��2&�30W�2��c3�93O�33�v3ݠ�2�t�3��N3�2K^W3�-�2,�&3O�2J��3c�43c 4��34�˄3��3� 4O�3{63���3���3Ij3v�3J4��"41a04��3�L�3Y��3+��3p"�3'4'�4��|3�4��;4D~�3}=�3_D_4 �3IL4��S3���3ڲ3�m�3g��3x=�3�ק3�4�e
4� &4���34��3��V38"�3V:�3�

4��3��
4�3ܩ�3�w3%)4"Y�3FΡ3���3���3
�N3L4*��3HG�3���3�4�4\�-4���3��B3$,4ٖ3�~3�X�3i0�3�4��3�|(4EƳ3���3γP4�+4i��3�ͧ3�X�3��4���3$�3櫏3B�I3$34$�4���3߷c3)^�2D��3Ǥ�3���3��3-��3BV�3k't3/�?4ѝ�3n��3���3�_54�p�3��3�v�3��3b�3�a�3З�3�r�3c�3�=4�7�3�e�3���3׬�3�(�3�-�3�?�3��s37'�3.T�3�e�3U�23�.Q3!�{3��&4>��3�3��F3�8�3��3���3��3}s;3��36I4���3ԉ�3(�d3܃�3�J4��<3��3�ؠ3�4��3��4���3�Uu3�D�3@[ 4E�:3w�3V�3��3�}�3=�#4�3�{�3د�3
�4�N�3�o4�f�3��4��3E��3��3{��3���3�6j3�`�3��4PFn3=�3��l4Z�3L��3!Q�3���3Z�4J|�3��3��]3i�3<�3��4��3��63�� 4��3��a3~[4m�m3�4�3C$�34<�3a�3(�3��3��.4qo�3:e�3��3�H�31�I3A�4���3j�3�
4�V4<a�3���3��38��3?-�3j|�3_�4G�3���3WY�3WH4�y�3B8E3��+38�E4�+3�.�3Uh�3舑3�{3��V3y��3��23r�3E��3}�34���3�Iq3(��3�ʘ3�`3��3|�733��3S�H3�74�Փ3R<|3.73&۰3�I%3NT�3#��3'��3o�3l[�3$�3�}�3��t3A"4r��3R!�3��3��3��>3�t,3�z�3�/|3N�3h�3Ϣ�3��3���3h�3��4��3c�~3T^�3T 4#ٌ3ɋ3.�3��L3�k3��3�X�3�!�3�33�x31Z�3��m3(�43?t3a��3�څ3_��30	�3䄗3_�g3���3�#3���3��f3�3�X�3e݄3_��3��A3�k�3e��3��3��d3�03���38d�3\QA3���3dJ�2�^3@�D3�m4�̠3���3"<�3�dX4���3U͖3^��3Z��3�:3T�3�Y�3�i�3�3�(4��3{!L3r3���3�3�u3��3�؁3��3�Q�3+�4�4�3��e3t]3��3�v3�_63�r@3��f3꽒3�_�32��3Oq3)�3( 4Vo�3���3�ON3Y�4P�A3߫*3��4�,3m�73�PR3���3~"�3�V?3��y3�4j��33���3��63�$s3D�3��3��33�t�3�#4��4Vܟ3��33��3� 4��K3S��3��3G��3@�*3�^�3pe�3�"3U��23V?4�0V3��3V�,3���3�n�3�S�3�/�3l�3�̦3�/4��3�`3�b_3.`�3��3>��3'�3mTf3��3$ȸ3���3bd�3�Jm3b�r3���3�)�3y�3���3�(4�~H3t�3VB�3XnJ3��v3Е3�V�3-.�3�O3(Z�3��k3�gR3�C�3�2<3�*�3_��3\ɷ3@7q3u�|3�93Y��3]$=3I�K3�;t3V�3`3]P�3�ƀ3�s3ո�3��4գ�3���3;
3a_n3м�3��$3U��3VQd3���3��X33P�3�?3U�F3��T3$$z4-�"3��3Pn=3�l3	��3�E�3N��3��3\�`3�7�3J��3�+?3��q3�#�3�o3{�Y3Sڏ3�^3L�3E�O3���3}?g3`��3��43�S�3DCe3���3&̒3V�3��2���3� �3�U3�,3�4��3��3��3���3%��3Z��2��W3�w�31�[3��3���3���3��3l��3��
46q3�؆3�>3h�j3�]3��M3��z3�u�3�I3?�3�V�3��|3��2l��3��{3U^3�P�3\3;�3�^]3���3���3�cP3��,3�	4��<3S{3�s3���3�l3J.33*��3�3���3:K�3U��3lA_3�-3��f3f��3��'3?:<3��3��3�Q~3m��3�H3��35�3{��3?�-3VR3��W3ta33�(3c��3��I353��=3�P�3�i�3"* 3K3Z��3�lf3���3�X�3��P3{J�3�j(3)f}3��38�'3�3�3b;�3�273Խ`3��33<b{3�H�3Cdg3͵`3��^3إ�3w|�3t��3���3��23D��3 ��3��W3���3ẉ3�Fh3)�;3��[3S�L3��3��3��4UB3�%�3d<�3�r3J�3��k3�3�3�=:3H�H3�)�3�f�3*l�3��3_`�3:
�3.��3	rN3`�y3��4c�!3��3:�j3�.73zc�2��4�yt3�M3�5u3&�Z3�A3"��3�[�3��3x^�3U��3U�3�]23�c.3v9�33kG3���3�	3u�x3>9L3:��3)�3�1�3��3I��3���3��3Α3z�p3���3pU3J��3l�F3T�3�)�3R^�3 ފ3�n�3�\�3Ȋ�3+��3�.�3�rL3�ä3��Z3	�4M�3!�3~#3��3ݴt3桕3�R3Kp3 �S3� ~3�&�3J�f3��3��4S�3hT�3U��2�3O��3�F�3~ X3j#3��k3��i3T��3�j3N;@3�%3���3T�:3��E3�=�3��3��;3��o3�	�3|�3��L3���3��3�̇3c��2뢼3�a3�*3,��3��3�3T�3��p3j��3��J3�*�3�x3*�3Mn�2��3c�Q3M��2~c�3�f�3�5�2�8)3��2�V
38�Z3y��2).3(�3E��2~��2��53	K*3��3��03%�g3��-3�_Z3ԋ3s�"3�H�2Ǻ3ke33|�35a,3L"3ޅ�2*?#39�3͝O3u	>3��2+9�3�V73o8 3ȳ(3 g3p�U3-3�yA3��2�-3g��2k)�3 �"3�I�2ݫ83yj3��2'3�(3q��2,sU3���3�;�2�#"3&�$2�0�3E3Kb�2��3iO3�r�2��{2��3���2a43�3�8�3�"�2=k	3͏�2Q��2�*3u� 3[P3�~2kC$3�]q3aQD3��3�2^_34m�2���2:G3�
3u�39" 3/3�P3�1�2�"K3�X3S�3*�
3h��2na�2:,3=�=3��S3�a3@�3L�M3���3��2i��2�iv3
`�2��2��3��B3��3�3!>3̍-3��3�R�2���3��3�s*3�0�2�y)3��3kg3`mg3�t�2�H=3d5�3W��3�j&3 ��2��2��;3���2�TH3��2Y-3��27f3��3?�3*;�2���3���2�3;�2��3���2D�83oB3e��26�G3ۜR3v�3G�32 1~3s��2�L�2B��2FR�2u&37��2��i3N�*3p:3�23��3�W�2��2���2A��2�5�2;U
3�xh3�W�2Nbu3��H3�O�3�S3ק�2T�"3�2���2��33���2t[
3j��2{�83��3�z3K3�221�3�3+�33c�A3L�K3��343��33�2��U3���3!r3��=3c��2L�I3HD>3��
33�+3A��2$�3l��2��'3�+�2�l�2-�2��W3�}�2`�3 38��2��2P�3��u3H3P�3H�g3��s3��*3+�2Gu3�H�2h��2Rd:3�2�$>3��3�;[3�36�k3Ѭ3,�e3)')3ܮ�3k�H3�hx3���3_�g3xD630�X3k�L3D{�3X�3߲�3Ĭ:3��3s�F3��03o�t3�F�3k"3w+`3�0�3��e3Oq<3uV�3�M4�
�223^73�{�3�_F3K��3a{�3�X{3u�3�Z3��\3`��3u�3#��3��3\Vq3d��3�73��2�,D3�3F6�3̜�3�@!3J��3�TW3J93o�`3v�v3(�,3��3�D�3x3�t3�4��3Xu_3��2�pq3��3!NE3vgl3M�83B��3�83�3�3�B�3즧3��%3-eI4��3��3�Uc3yb-3F�13+Mu3��3p�2o=3���3.r�3�3�*&3�D30�3��W3��`3�6�2Q�y3�3M�3�,Z3��2�v3�C�3/'3x�e3 X)3���3��2;�3�&�3���2��$3�k�3��{3�~u3�\�2e03�kV3f�3�<f3Zx�2��3~�2Uu�3��,3�8o3�K�3sw4A�s3��3^u�3���3�h.3�=}3��3���2�Y�3��3�(�3(D3'}35�u3��83�o3%��3]�03�=�3<{O3(�3��(3ѻ3ܴ�3�i
4��3�B32^s38K3�Ea3A�X3v�B3E�E3��r3&4OU@3���3%�	3�M�3j�38�<3�ci3���2�3�<V3�E�3�-S37-�3�}3u%�3?�3�s3�83x�j3E3\3��|3Ve3Յ3��?3,T�3]�3�yz3E�2�T3�lL3?*3�|�3p�
3D�3)��2�:4Y�3��3gm3Z�	4��E3'�3�^t3��23ʑS3�MK3�3r^;3��l3 $�3�'�3Ww�37�$3)�3�Ǔ3�P�2j��3-O3��3%�F3S�3��v3�>}3��83 � 4i63R�33�l�3@E3-�3��3�q�3(,3òo3�4�3���3'�3�0<3��3OnC3MfX3��3�3?�3�;3� �3�j3mP3� �3p�d3��'3���2��3�ɺ2��&3b�g3s�$3P3�^�3��i3v~�3<oH3�ړ3�Ƞ3�A/3L��2���3Kw�3��3�Ő3#ߢ3�a�3�J3�t3׏�3�o3��3_$3�3dSY3���35Jv3��%3���3�VK3�)3ե 3���3Svt3d�3H�G3�73��Z3@)L3���3��X3mA38;3�͇3���2��03I��2�lQ3*�3�:3N	A30.3��03�35�3ނ63q�2�/]3��V3s��2=�.3+�a3%�43%'J3��T3��[3�wW3q�N3�@4�=3<��3)��2x�3C?3f[s3���3�Q3ɜh38*�3�O�3��f3i�3Ic+3��3H�3�`�2�FJ3��p3e�2+�?3<�G3;XJ3�&�2ã4L�3�2��,3X�+3�{.3�L�3��\3 �2�23�c�3�4�3Z+V3���2w��3tH13>%$3,
U3l3q��3�3��u3-�h3��03FH3&��3�,�3ŝ�3��2��3#̓3H�_3��_3̦3e:3��{3E��3��3x��2��3�fm3s�3
�E3 &�2a�3g�3��3ἐ3c�3��L32��3�3��Y3�!3]DR3=�3��e3�03��$3���2GH�3��]3�B33�d�2��3�x3t-3[��3�H3��13�	3�F�3C�)3uƑ3�Q3`E�3��G3�>�3g��2�"3w>3�fM3�Y�3v��2	;3EC�3�-�3�lO3-G3:�v3㩐3��3E��3_��2893؇�2���3�38gF3�y3��3�V3~�[3���3��=3�d3tzO34833|:)3V�x3��3�63�k3Wi�2'�s3j��3@�O3�+39�3zEq3�o+3:��3PU3Y �2Q��2��4b�(3�73�=�2"�3T,�2,>�2<3$$3�ߕ3��3�*�3��N3h��2r�;3!+93�~=3��'3�{3 �E3%O�2 %�3L?3@��3G�F3�T3ᛄ3���3%T�3q��3&>43Ϝ3�Q�3!�F3�E�3�84~�X3��3o��3�e�3�d�3��M38d�3-?�3���3�`3Ӵ3�y�36�z3ŋb3�4�
i3�S�3UH�33Q��3o�3m��3F3C83���3��3P<�3��38W�3��39w3֙3(lE3�5�3�S�3p��3�3 Ҫ3�83�p�3��3���3�l�3��3/��3�"K3]��3�<>3�3�]�3b��3�673w��2^�3�pA3�Q3���3V"�3,�23r�]3"[
4(*3��b3���3���3Q�f3]>�3�ӛ3�P�3i��3���3��w3Z�-3[��3�D�3�׏3_�3TRl3��3R̶3J�A3O�Z3U�3G�[3nz3$��3�c03Mi�31�2���3\ד3���3��3��%3�L3�9�3G��3\��2�J?3�U 4ii�3�x}3�_D3ju�3\ɛ3��23� �3�N_3��3,�@3��24��N3/6k3�9�3�,4�ؐ3
�3��3p�3'E�3�Zi3�X>3�32;�3�O42Q�3��3��3E��3(��33�>3MRa3mg3=3�3��38��3�3v�3<o�2=wD4激3��]3�b�3�/�3��23䑥31T�3�_03	�3�4���35.3I�63�S�3��H3��3mЕ3u3��3�.3�*�3��23�A=3%�3�3�� 3#�83
�;3��g3:X?3�.�3�և3|�3�3ū�3�M�3�j3Xy�3);�3]sz3
al3��3�#t3��3��3�"4a�a3�}�3�w�3
I�3· 3��3�}4��W34s3���3�?�3ߣ3>��3fc*4 ��3aq�3�8h3�&�3�h�3�jS3���3E�F3zC�3b6I3� �3�w23�G=3R�%3�S4;�*3�93)5,3�mP3��Z3�a<3��3єP3N��3[˙3q�3I�)3��3+��32�3�6H3'kx3>��2��w3&(3�.�3���3�Վ3��.384�mU3�B�3>�a3���3x3��3a�3�~a3'�|3�3B?�3X�3��936)�3�4m3�Z�2:>3�4e3}��3��	3���3�yK3YOT3��3=D�3��;3l�=3�r�3��a3���2=�+3�k83Q�63�Kp3c��3x�3D�3}��2Mb�3�k43C 3��_3�f3�/A3
3�8a3�z�3;�Q38A�3е4!�3t�3��v3pڥ3�H 3��+3�|�3R53�/3Ws�3�B�3h�3�s3�;<3+u3h��2�͕3H3O,33��"3膄3-J3��x3��3�D40k3,�83l�3ha3�nF3I�3�g�3��3�6^3w�3v	�3�~�37�2|Db3ZM�3$c3G�73�	j3˔�3o"&3��3LY%3�#I3���2Y�3>	]3��732s3W�3�3�	�3#�J3k�b3uUV3cn�3睚3���2�^-3%�3w��3YKQ3l�Z3�3��j3<�>3��3�gc3��r3If3�#�3}�c3�@3_~�3��_3 53{3��3C^�34Kq35�4"��3P3���2Qe3vF 4�jS3=E3��!3J�o36�$3ڑ3�,~3VY�2*�b3u�4Ůc3�#�3Xwx3��u3��3Q�W3GRv3Pp 3���3vb4��b3-%3�#3*�3QqI3�43�@537�	3�)�3��T390�3
3Q]g3�g3F�~3#)�3F̂3\�3'�73I43��3D_3�3��b3�W�3��F3\��3.�3A	�32�3x=3�z3P.;36=H3e &3<��3)�o3^�3廁3�64�t�3/^�3	�	30�W3X#j3�B3f�r3�A=3�P>3���3�jv3�p+3�g:3W�83z$34a�3U�3�#3��I33�Z3��=3/�33��-3��3r�]3�U�3�n3M��3�!3>!#3�9b3I�3�{t3�M�3�!o39�P3C3�N�3���2�U3`N�3b��2��g3d�3��3h�3��3�3�3���3�3M36�J3�j�3��?3�Zn3��3#d3��_30r�3�}�3���3%q3�<q3��>3�8D3��3�ɧ3�3{&Y3	ɝ3���3�/3�Vp3,�4�x3��3�Sx3^}*3�FH3*or3}��3��Q3��<3�k�3o�N3��3A�3x6�3L�93U7�3�9�3�W53�ѓ3=Q3&�73�R}3���3ܮG3�,4[�N3�{3�Qa3(�3��*3
�3a��3�13PA3�3��3�E]3/1I3�r�3�E�3��3?V�3a	3���3A�/3���36�3l��3Ǉ�3��4U�G3��$3�K3dAB3r�3|�3���3��3o��3+�4xU�3�Ė3η�2���3?(o3Ш�3,I�3�JR3|�3�q3�J�3.e�3j�B3�w3��3x�3�L3ǜm3�tX3{�]3��`3��3��3��3�L�3�V�3`��3�r/39x�3�5�3W�Z3��3��<3�N3��P3��3 ƽ3SZ�399F34�'3���3!ދ3�3� 13�Y�3}f�3*n
3i�\3�O�3�1�3?SW3�@3ԑ47l3b7�3��\3��;3rv3��(30��3_�+3A13A�33�N4���3΀3�]^3�L�3`0o3�{o3�C3�;\3�[X3�O�3=H4Y3�*3�~�3�3�3)�	3ŀ�3n*3-�53~;3%��3u�03���3�[93V~�3#c3�~�3tl�3��3��H3z�M3��3��F3��3O�3�]�3.��3́�2+�k3�(�3��23���3=ј3��3��43�k�3��3"�u3��+3��%4���3���3���3t�s3�y}3t�3g��3�%35��3z^�3.�>3��3���2�tq3E~�3�/3�r3VV3fO�3u)3�J�3��3�]�2�13@�a3nSD3��13�&33��43�_;3�l3�*�3r��2��i3%"�3ʜ�3��3�%@3�o3��R3�3�g�3�83��33��M3c�3Œ93�3	�,3�Ȟ3-4�2/?o3�"3�ރ3a��23�I3�3�d3}P'3]�3�=�3,13>Z3��V3��[3&5�2�m�2R73KY%3O�33��3��?3h�Z3B5+3,L�3�83Ⰺ3�'L3*�3(��2u"�3�k3�P3��3�N�3$�3�3Nt�2 @L30�	3���2r�3�,3#}U3��3`�3�?3�K3��?3�Z�3��<3�d3��3��3�3I��3۩3sd3}$3Qt�3^3>l�2�	3�}C3�3��2��63��	3�ǉ3'�2��U3s�Q3&3��?3h��3i�2�n3�#/3��H3�F31OG3ph�3�� 3�D�3]��3�z3x�3dy3ҞF3�3�3�>3�G�22�g3Ak�3�\,3�ޏ3��2�ի2��#3dU�3S�3��@3�y�3�d)3�tk3�%3_�~3Fd�2WN,3���3��3d�k36P�2�\�3���3Y��2���3FM�2^3|v<3#�3w�3B�a3R�`3�!�3��)3�4�3�,^3�3���2�~W3Hyr3v��2��f3�e 4c�f3��<3�9'3V�3��3X�<3c''323�g3�3�޻3Ŭ634�*3�2D��3!1b3c�2��#38h/3PV30�\3�˗3��.3B;/3 8�3wh3E &3*��2�`c3�~;3�5�2#Q�3�3-�3833��/3U�2�3"7*3�d�3V83�u33j93�@3��3��B3N/3v��2e��3�r�3Cф3ۜ2�c�2+�;3V8*3�G3�R�3��3ϽR3y� 3j\�3p3�2?�L3�&$4
�35x>3�&-3-E�2���2�3Xf3z�3��3hX�3�+3��t3��3~3}p3V�r3C�<3j�E3��3l�3~"u3n13#�2?�3҇�3,r3�D3�h�3�a3��63��3ֆ3�3T��3��3���3��g3Z"�2b��3�=N3,43���2bP3�>83ަ'3��83��	3r�47l�3�84�[�3�3r��3�t4��3��4?�64�3;�3:4�ά3G��3���3ߑ4�J�3O�3���3���3b=4`oa3�u�4�C&4M��3+r�3o�54�^�3M%4�D�32��3V��3f��3Tc�3�e�3���3�!-4T�4u�	4̳N3�)4x�3C�38j�3�iW3�`�3��v3��-4��3�r�3|�m3�;34'�3��3�I4��3��3���30��3�(e3֢3i�`4�K4��4H��3Z
4UY�3d�3���3E'�3S48�Z3_�'4l��3�G4^}3�Z4;��3=�3�4G��3���3)m�3�F�3��3-o4�zh4�'4	�38�3���3�`4�3���3}��3�:�3a�3c�?49,�3�p�3�4ҭU4�"�3�b4�'�3.M�3��3]^�3Z�64��v3���3k�14*�(4#��3��3��)4��38	4� 4�ř3�v�3n[�3�	44?Y�3�E�3���37�64J�3%�3�?�3�K�3���3؋4��3Yț3���3�164��3e�3��3Y8y4�m4�ۻ3�4L��3��4ѻ3v�4L�4��3�#�3'�e4H@�3q-�3��%4I4�_4���3�4(F�3��3�AY4��4Ҿ�3Y��3���3a!�3Q%�3�g�3fܟ3���3��l3�sJ4xը3��3�h�3�1Q4Shj3`��3Bj�3���3{��3y �3�+4Z�3'�4�C4Go4#�3c�3O!4��4#�3��4�� 4��4*/T3�=�4��3��3�|3��4gC4p�N4���3��3̇r3��3Bl	4�ʏ3��4(�S4)��3�44�=�3�x�3��3��3���3�{�3Y�Z4�n3��j4Pw�3yu�3(�4�/�4��3��4���3���3���3T�3{�4�U�3��4���3TZ4V7N4�9a3�4���3�,3��3wE�3���3��3�J!4m��3Ɏ3�Ė3A04�B�3�7�3��!3��3��E3�T�3�V�3*��3�ۍ33��3��s3�5�3�ta3��33�3��3��3��3e|v3�wY3�
�39�3K�3�b�3s�4���3N	�3�@U3�4�3��3���3 ޹3`xe3
�3���3���3\�3��"3�{�3�`�3���3���3���3�@�3�U3̋�3D�3�h3���3��4�z3@n�3�3RK3el03R�3+d43��3���3�3�3���3�~3/�3���3,.�3lW@3!�w3#t3���3}E^34��3c�3�T�3�k�3_H4߈{3^I3BR�3ݬ3��3�Qv3�@�3�@�3t[�3���3�#�3`��3�3��3��K3:�$3� �3)��3��3(�}3�Z 47u�3��3:/N3��B4˹�3�e\3*%�3|�.3�.�3m�3o�3}j3��3�/4���3*:�3��B3
n�3�S�3S�X3��3t��3���3�n�3��O4��,3x��3�1d3��64��x3vA�3/<}3T?48��3)F�3P��3	%�3(��3��3}J�3���3v��3r�37<�3YN�3��[3[[�3��3��x3M��3%7g3�-�3��3�$4��3
��3J�93��O3w_W3���3qղ3M�3���3]�*4}ӥ3��g3�H[3�8�3��3��93&�3�LA3�Q�3�4�3Q.#4���3@��3#o�3[�O4�)�3̈�3�3�0�3�!]3��3�a�3�'3%5�3�O4>��3Q�3��(3~a�3�x4S�3{<�3�13��3�3g�4;��3D-�3#��3�"�4���3L(4�/�3�Ԟ3�u�3��3v��3�J\3I�3��3��4�!4֬�3)�3t�4x�b3�
�3��3:>�3�|E3��
4s/]3B)3�U3~��31�N3�3��P39�3�#�3�y3Aw�3v�{3��3{q
4���3�X3u�\3<�4r8�3L�L3���3@��3y� 3���3���3��31�&3���2R�G3�S�2[�-3a��2[r	3�.�2��13P�2�8�2���2�[53�r37�21K3�X53�:�2B6�2,�20@	3÷3J<�2SCb3�-3L�3��2��	3���2X��2�u3#ʯ2��2?z�2�93��2��3�C3H��2Z 3S�2x�3x��2%Y3�3��2���2T�3��83���2խ53��h2\��3F'�2it�2uk�2���2<�3�%�2�$,3���2G�3�?:3�3��2��2.�3O�!3T��2��3J$3�43覻2t�3��2�(�2��2��^3S4�2PQ�2��3��2f��2/�3��3{S2kV%3vpf3'H3A.�2��l2�,3��3�ǃ2ed73�Z�2�
3Z��2Wi53�%�2;�3�aN3��G3��3E��2tي2g�03 �2'{U3�/3�V�2�<�2�|3��E3;�*3l{�2z�E3�3��2�%3.�)3NY3�;�2,'F3d��2��23)�2ć3��2�M�28�33��213�<U3 �3� �2��32le3��%3�B�2���2\#3�[!3�a3U��2�}�2�lI3�[�2�<3�q3���2'x�2�݄3���2j?�2�* 3�3p�K3��03�a31p�2
x3��x3�Q�2���2�D3��30>�2�م2k�3��2dP3k˷2Ā3>��2���26F�2Nܔ3O� 3J��2���2�(�2�3�^3��3��2N3> V3�� 3��3Y��2K�3�]3&}�2k
�2���2�?3�o�2�+m3�%�2��2�\�2	Z�3z3I�(31�3?=�2f��2 r23ۏ3a�{2���2Ny[3�$30��2�2r�
3��2a��2.�3��#2�63�̵2"3��34��2P̳2���3�Z�2J��2���2z��2~��2(�3z�@3�D�2���2��3J��2�� 3�0�2�Y.3Q�2G� 3F�Q3�@�2>,X3��31�3�r�2�+�3��3�is4�'�3 �3�c3xtk3O3���3�?�30�3��3К4��e3v��3���3�D�3ApS3��I3�i�3`A3&�}3��K3��	4��3���3u��3,
>4�b�3�KN3��3�!�3�+�3��4��3<�3:��3���3Ч4���3��3�(�3b~�3�`�3ƛ3v�3�G�3�ю3��4��4��3�M�3��"4vۮ3���3���3Q!�3�,�3C߄3��3��3ҡ�3�_4�%4���3H��3��4=��3��$3�$�3/��3^��3�֍3��3�K�3���3I�93���3�i�3v��3��p3��3�1P3 ��3�#�3KF3���3A�J4���3�\p3HGU3�3�H�3}m3�3;G�3�q4]3�J�3�N�3�Oc3AF�3��4�ժ3��b3���3���3���3�Њ3$,�3Mi3g��3s�Q4.4Y��3��k3�e�3��3u�3���3g�=3{B�3���3���3��374ٿ�3�;E4��N3R�3��3�J�3��u3A��3�-�3���3�� 4{X(4�=	4k��3��3կ�3GR�3:��3�7�3���3F��3�ܼ3'T�3�2�3���3��13�Ղ4���3�T3��3,}4�B3��S3I_4}�3Z�3�{�3���3ѳ[3��\3{�3�s�3�<3�3��2*��3/ n3��4Z�h39�3�t�3��4j�y3��3���3~ػ3���3���3va{3��3�3R�4�t4��4��_3�~_3�i�3�lm3�3C-f3��3�
4��3��g3j�n3@�3��14kӊ3㉷3�J�3��3�Y�3�R3�W�3
J3�3Rh�3�3>|3��53c}3�3�R�3��3o�3[��393E34��l3
IZ3+�3O��3 S;3֤�3�h�3�S�3�_Y3��z3&�3.s?3���3P1�3�̸3E"4�dh3��E3�� 4h��3+��3}3�[4��r3���3�_�3���3��73K��3��X3	�3A�o3=�u3�(3�t�3vڦ3|`�3�VI3E�M4\1C3���3J{�3�4�3�1q3���2�+35ށ3`k�3�33�E�3��3���3�(�3S�4Gk�3�3`w�3I�3�>3���3B�4�/A3�
�3pe4��4�g�3O�f3̏�3��3�xB3���3��3E�3�3;u-42dV3�َ3�OI339�3#j3`�3_��34y�y3vj3Ѯ�3]U-3��3#�]4�e�3�q=3B�3���3H-3�53��3fv33�|�3��<3t�4���3�z�3(�3P4s�3�i3s��3R�3��3���3�F�3�I`3���33V4�� 4���3�t3T�3�X�3{n>4*%�3?a]3;#k3cD�3���3Wj�3|jr3^�I3�#4�W�3��3?�3
�^3��i3�h�3/n�3�oG3�0�3]�3���3u��3��m3Ո�3�i�3�*4��3m6+3݆�3~(�3��3��h38pf3��e3�54d�T3xO�3KA�37�3�R�3-�3w��3_%A3��3	�3h��3��3�(j3� �3�]�3��u3#�37R3���3B�3��w3�[�3��3�E3��a4��3E�3�J3fp^3.J�3]�3c��3�V�3Oo�3��3î�3�=�3�uN3壣3�O�3���3�M�3�GV3�^�3	�|3���38n%3Ɔ�3�B�3W�`4�m�3��3~��3�dZ3܋3+��3#p�3 1�3�۪3.��3"]�3Po�3��>3 ��3���3B{�3v��3�u3��4�M�3�)4X�c3"Ϯ3}�Q3��R4�3��3�3��u3
\3���3��3��]3!g�3�s24)��3	G�3��~3���3*��3^�3��437�3'�3��U3��4给3XVA3섂3�j"4��c3AJ�3�}�3���3�|�3Z��3O��3��2ki�3u��3���3>�3-�/3�2�3�L�3��d3z �3f3���3�Q�3���3�93���3II3��3 xR3S�2r.C3��L3�cA3+cd3�gS3Wr&3� V3�E�3�t+3��M3F�3��X3Ma3h�e2�:33�3�_d37�3��|3���3ۮd3�_�2���3�pA3�=�352�3�+3�ׁ3���3���3\@`3k=n3n��3���3�N43E%3O��3}g 3�o3&�R3�L13���3I�G3���3?��3�63�y+3���3�D3o%3��u3��3R&�3tC3oJ�3% 3��.3��p3ks�3ꦊ3�=x2!ߣ3̗�3���2���3���24A3�;t3��3j�32^3.߂3{%�3V�J3��q3�	�3�bw3�!f3cT3}s~3s-.3��3��3.{3�RT3q�3��b3EJ�3yA�2��v3;�]3%��3�@$3���3`��2)`�3Z�<3P�3��3��>3w��3��3rh3mۄ3�):3��s3�K3.��3�.3��!3�{^3�xA3s��3�Ӱ3y 3�|D3��U3�=f3z3Pt(3t�"3�6�2��14�z�2�?03�ec3@�3{�[3n�3Gv3�Yy2�$�3�~�3�g�3�yj3��2K�.3jg|3cf[3��I38SB3�oU3ȁK32I3�X�3�J3�e�2͢4��^3�r13�F3}G3�#3�K}3(3��<3�3��3U
3N�B3  3�r�3�O3��.3dʊ3�3�Ն3Xu)3y��3o�#3)U3�'�2��42e3��330�A3L3�đ3Vʩ30��2�6�3�C�3+Bd36>3W(3rgQ3�*�2���2�^3j�m3�U�3%?'3���3��s3��13�f3E��3}x�33�s3�L�2�
a3 �v3��3��Q3���3�}�3�L�3Z�)3O�53��/3��38�E3gm3�/)3�"�3�Z3A~�3b?N3a�3k344�3 b3�T�2a�<3By�3WR^3�W3��3��3�$3��.3pU�3�(3M"33���375a3>�?3;|�3���2��V3��%3�$j3�ς3V�F4�4�3�P�3�3�ġ3�`3�@�3�h#3���3Hˣ3 �3 �Z3�148�36��3إp3���3�s3e-3�p-3^�3c\�3J3�#4k�y3N�3[�m3��4��33.��3�i3��3:b3~��3��3l��3��)3U3�3�0�3�C�3A�3*ڴ31T�3{xo3�p�3~[3��3?�k3M�3-3�Ό3�H�3te�3�U�3Ԣ3O>3pJ�3)�3�E�3��30�P3:�3�$[4�y 4pQ3D`�2e9�31ܹ3�u)3���3�;�3/��3�F3dS�3EJ3~;�3�S[3��4>p�32�^3���3mu�3,��3+l�3z��3�3EN�3��(4���3.Ga3-�3,�}3{7%3�k<3���3P6W3��3+�73��4�^�3.:3�3�A&4rʒ3���3�b�3t��3�>g3�Z�3Շ�3��~3Y՗3$��3�4[�3M!3��4��4�Ң3��3j~F3��3w�3hǷ3���3�1Z3��3`4���3�0�3���35�h3�33g7�3��3�V�2 U�3-є3��3'?�3);w3���3:i�3�3Er3��13�~�3X�s3�
4�|�3���3��3�4'��33Q3�Q3��3�3Y��3�˸3���3	��3��4JZ�3Qw�3�#3��35M3�S�3��u3�u73A�3��N3���3��U3�p3�Z3���3U+y3�#h3�3�}3�	13�a�3a1�3Ǝ3�K�3p��3�G�3
Xp3��3s�3 ��3M��38�M3q�M3y�=3;7a3T��3��C3��3��X38��3~�3�I�3���3��R3OJ3�_d3pxc3��Q3ܟ3m�4xe�3�/�3B�3�#�36�g3I;�3H"�3I["3S��3�L3!�3�ˉ3�� 3�i�3�h�3��n3�r�3>��3?�3^ƃ3�²3���3QH�3`�4�r�3�E�3
�4���2��3���39�|3��3=�(3��3&�33WV�3o�3Hdo3���30[�3Hl3�H3:�3��3 �3Ub�3��83�d3�D�3�Î3��z3�T3��p3�C3}v/3:�3�c3��F3��@3۫w3��~3�"3�83IMc33�3��^3jLL3�/P3���3�433��t3��3��z3��533�3M|3 ם3@�;3��=3�q<3u�?3�,:3V3���37zK3�z3"�3���3���2�qy3<>�3~��3�;3(�x3-;73S��2T�M34:��3��3��{3��j3�633Sف3��S3���3d,3}i�3y�;3���3�b3�m�3�3�3-�M3�tc3ʃ43#�2�ۥ3��2��34�k"3�M43攳2.�\3��3K��2nc+3�տ2c�3c3�4N3�pF3?�%3u�=3��4��z3�;}3��303|3`3�GD3��-3y�N3[�3�i3W�-3:a3ؕ3<;/3�j/3�]�3+�/3�fX33��2��D3��3D	3V�P3e>�3t�C3�P3��"3>�\3Hz3�q�3��`3+�2��%3x��3d%a3%13�3�26:�3g�3��_34��3/�2|�3@43v�^3ZwJ3�F>3;�3�S4�dY3�m(3�b�3��&3>�f3�ua3�-_3��3B_�3u��3�3K3�_3/�37�3�&Z3� �3t"3�O3_Z.3�3�W53ųP3��31��3>rB3 �3h�n3�(R3�3Q3��D3l^\3FiA3	F�3�x�3B�3�ܓ3�`3a��3;��3�3��3ԭX3��3��2�L�3|�R3�=3o�Y3��3��3��3�ԃ3�L3��%3�~i3�k&3v�3���3(r�3�i3���3�o�2���3@�P3x�*3�~3G83-�|3���2%�3X/l3��3M�D3�0�3%V?3��s33cv3 n!3�z3� 63�!3��3���3k��3�q�3�3&�I3`�3c�3�33���2<�3��?3c�3�]�2��O35q3��s3�#3�<?3��3lg�3*��2�׈3�C3��2C��2�d�3��V3�&}3��3r�3�5�2�$-3���2/�\3��`3_/3˟30*3�OC3!�93�C�3�`3�\L3z=L3B��3��J3sBJ3��3\�3kk3��3���3$\3��3�.T3�^3j~�2�w+3��,3mZ3�(3b@�3�3[�3"3�h�3�� 386<3λu3s�3��*3t3dm3��3OT3Q��3��C3���37e�23hN3;�b3���2�D(3��	3�ԩ3��W3�;Z3�9<3%wR3��3: 4��3��
3�_�2�B363�z3u�c3P�3�(3�x�37R"3��2I��2��3ZU3��Y3��%3p3=�3V� 3�JU3s��2�'3l�R3�Y�3ʃF3��3Ǔ�2D�3"f73i,3D�L3V�3��F3��D36��3�p3��2(Bd3�sX3]��2Y�33��2 �83T35=m3,�v3��2��3��3�H3v�M3U�3C�Z3���2�~3c	A3��23{�3NZu3�c3j&(3�3�3�j33S�2�w3�U�2W��3̃&3c��3Rs3�+3��2ve�3d?3�3Ƽ3�N
3�~�2C�E3�@3Tv�2!O3�'�3!B�3�� 3	��2i�53T�D3�83:� 3���2���3=�3_��3*�3��3�
3aw�3+�3��H3��3P�&3�d:3��2��n3Q��2�_3���3��b3�)3!Q�2Y�J3E73���2`zD3��3匃3��3�Y�3��$3�yu3�Y3�L�3��o3��u3/>�3���3���2��V3P�r3c-�2/)G3Q��3�3
Q
3�33��3��2�2'l�3��2Q�?3ͫ�2�=�3Cj	3̲3Sv3<�(4`:�2�A,3��3��3��)3��?3� Y32�2�f�3�L`3jT�3��D3{��2�f3�]�2'� 3��3�Z�20V3�?3���3��3�:3EWR3#Q�3J\3g��3�aq34X 4��o3+��3�~23%�3}3���3�r3�=�3�k3)��3��D3�)83w�3�E3��3+�!3��3��B3��3��3A�4�3�E3��63�av3��R3#�3n�3�a3�v�3�D�3��,3��3�Z'3���3Q�3zu�3~��3���3�3�^K3�{�3�L�3;�K3��3[7	4$3W533$63G۞3��p3�:63��3�T3e�3e2�3)4��3��3�j3�7�3Yv�3f�X3�Y30B�3�`;3��3M�3��36r3W(�3!|3�Hw3��3s��31�V3CLq3v��3�oI3ro3��3�~3�zZ3*�#3C�3��3�3Оv3��[3t��3��n3!ȑ3��T3X�J3�D�3�z&4A323��t3ߨ<3��3]�Y3^�i3kNw3	*3�+%3<�3��3p��3=�W3[�3�WS3��;3^��3�'M3��^3��_3O��3+�[3�3:3
�73��3���3d4�3a��3[��3�3�g3Ϲ�3KA�2���3Kh�3 	�3�ZJ3)�M3_Ĭ3�#�3��3�R�34�E3Ζ�3XG3��4��j3"v�3�3��3�J`3P]�3GLt3ц3�Ǩ3Ϧ3���3��H3t�G3[��3�33Vr�3��:3DMW3.=R3�*33��3�W3�	�3� �3� 4�3'd3n��3:�04�$3�ʁ3$��3��3=083E��3%�3 ��3��3 '�3E¤3�6�3�!U3"3�3|Z;3�_�3�ƪ3�l�2K�Z3&�?3�3���3]'3�+3�$41-T32�3 Ԓ3�K3�3��4MQ3�3/�~3
�	4��3��3� }3�
4[3�'3Hs�3�_13�3u@36��3�l�3�$03]0A3Sٔ3>3�h^3S��3��r3,�i3��31��3�y3��F3��e3&�3&��3�V&3���3��3��3~H�3 )�38?�3eE3��}3#H3�
4��f3v_ 4#Uz3}v3#m{3�uK3vH)3%>3:'�3�$3��b3B�
4ܵ�3{ޅ3��3��3;̜3�L3�l3is3F"�3t/3Ŕ�3n�3�9�3@M63�24Ӻ�2���3���3�3}[_3��3�·3��#3��o3 �3Ih�3!��3|F3f#w3\��3�3��13y�I3��3�ן3?�30�3��3��30�3��73��I3�!�3Dz�3nG3�&�3��3�r3Ks�3k�"4pT�3F3�<@3|im3�u3qT3�!�3�53,��3��?3뇖3S
�3y7p3�P3,l34��b3�o�3Y=�32�03�3��3;�R3�~r3+�38��3�q�3�i�3^�2}��38ӓ3ws�3:Ύ3ﾅ35��3��3!��3Z�I3��z3_�%3�$4���3?'03�ڗ3�l43!�3�b�3	��3s}7322�3a��3��357�3 �.3��3q�c3t3�D�3M�a3N[�3Џ3�T4]V]3�7�3CG3q��3+z�3�Җ3bN3a��3�lt3_��3Ȗ�3��2n�3��3��3!֜3��B3c�3i�3�43��3ѩ<3Z��3=�V3�Յ3�E_3�<$39�3��3Ȇ3�i3f�K3�G3 �3�k\3�"�3��@3�ڿ3���3�]3��34Z3H��3ڰB3*�83@�73�KQ3!�34�P3�8�3��3��73JL3�h�3i+�3�&�3 =�3�@�3�	q3k<T3�Ԙ3��3 ?�3��'4�3Uf~3N�3�S�3�JN3�$R3:�m3_bF3�ģ3�G(3WC�3�fc3�~D3��3���3��X3t�y3G�3��r3���3Y4�3y7�3��T3�j�3W�3�B�3�4�3b?3���3�@�3WmU3�]k3��L3��4V�v3��3�y3:N93��3�4U�X3,�j3��3�p:3��*3�i�3Έ3+�3<��3-i�3�̛3�I�3�-N3	g3(�3ѧ:3�g3x�R3~*�3��R3?
�3�k3��N3�X�3W��3zS3�D0383A>�3b*%3�Ǆ3�$s3N�L33\d3�k�3H-3�'K3�)v3���3N[3�33�K3�Zb3a93��93z;�3�{3��3�e36��3��3��T3 3�N3}��2�q3�َ3T��2>��3e��3�eZ3�y3�13��3��#3x�3 d3�f+3�_�3os%3�3�3]�R3���3���3;��2��83��43��35�3��Z3���3�l13�U3�F�3�NT3|�53�93b�3�lh3"x�2��:3
3F{�3�<3��3�<R3+��3QJ3��4��2��B3z�#3K�"3)
3���2J�83� �2p�_3y4��3}��2��2�o�2qE3Ё53��;3"�3��c3�0�2 7m3� :3��3���2�G4��]3�+3CU3�'A3f�3q�3�P3��2�T3x�d3���3�U�2��3�+3�G3�!�2��63;��20�P3��2&un3ȷ�3s�3)4I37^�3��C3�83�	;3�	3�X�2nG�3��$3i�3'�3��3�O�3l�33�

3~]38T�3	��2��`3���2��I3���2�$3&�)3c�3�k�2|�3m�53�I�3	3��3ٌ>3�/3	(3��=3;�(3 &�3�_I3zgn3@S�2�u<3�_3��13�(�3�q�2+�43c�+3�z3t5<3Q�Q3�m83P*�3��F3��3�r732�53�p3.h3ߋ�3���2��3���3�vZ3��o33g�G3I2,3s;�2�֬3�o33��&3�3�v�3�383j�f3�s�3Nʃ3��S3��{3%c3b3_�3A�p3R�
3�3�]�3���3V��3Q3�9j3:3�5)3���3)>�2}��3��-3��h3�v3���2A��2�4-3��2T�g3f��3=��2e��2GF�3`l3��W3S��3���3��*3a��2i?s3�IN3$3�FK3�`�2��z3k8�2�Y3��13��R3z��3�+�3`,3��]35��2��3P�?3G4�3H�?3��3��63),3��2]�3��E3]M63�E3�3�3jP3J	G3`,#3f�3i�(3��H3�23!��3�f3�93JfT3��\3�3`�"34�m3'�3�Cs3)��3�Y�3EtN3Y�3d~3y�{3u�W3��3��3gF>3��]3M�3��3�[3���2�)�3b�3l*d3�yK3F�"3F�-3ꕈ3mǁ3�33�D3+4ٺ�3�� 3̠�2�	�383٪3�3^3�23� W3�J3ع�3K(3[�3�\13g�4�[3�_3���3>�3I�#3�yM3ݠc3�=�2fD3ě3b�3 ds3d�3Vo/3o�Y3[c'3\�.3F��2p�3�\3�҅3��3�~�3C�3��3�r3���2��3�[H3T�=3q��3�w�31+3��3Y��3x8�3F�H3��/3�i3!�3��\3˷�31�3fڤ3.0Y36t�3��G3��3��3x[�3�:l3��Y37	<3R��3��2H�,3���30��2��M3�9�3v$�3�v3B�/3��3y�L3�/3r�M3�]�2�V3�3��3��?3��	3 b3�o�3%d73�j3f�j3�p�3�3Od3�l3��\3�`3�r�3��3�ށ3��3�3�3�83Y�3�z3��:3�'w3�M3��3��73�q<3H�23�~�3S�3w?T3Pm.3Z�i3v93>@r3&�R3]�+3�dT3VR�3�!3���3�3��3�;63�23��3N�93��3z+3Ad�3$�T3�z3�$�2'�3�%3h3,�3�g3�>�2C`3%�-3|��2�}I3��3��93r�3�� 3̳k3K��3���2���3�>3�3���2��3A3�~%3+�L3`,43�#3�zO3�H?3w�.3_�X3J�=3ײw3%K&3��3X��3���3�t3!��2gp�2��437?=3�q3b�2(͑3��2Ǧ3	f3�?3e�2�O�3D�V3�x+3�X�2�@3�Q3X%Y3vH3s!3ݓ3��R3�53��l36��2�J3b�:3���2L��2+6-3Yl3̓3��3�Ӄ3�@3L�3�Il33p93$�M3-�c3ǌ�3h53AU$37�f3�S3�Pa3��3��3J�83ㄪ2�
3�f�2Ջ!3��]3� $3i	73eN3�{,3
b3q��3z5-3�y�3SJ�2AQ�2z�b3�%3[��23<]3�3a��3G��3V�q3c:(3���2qRZ3�yp3YX�2;%3
�26�L3��2�D�3��3��b3C�3Z�3�83kT'3(3o�@3� 3��X3�A3Ԗ�2��[3�c�3��3� 3A��2:�F3�G3R3��`3�$�2k�^3�3�*3���2VP 3�  3���3�j�2�%�3֑.3�3i��2I353Z3GX3v��3�n3M��2
�2��t3"�A3^�73c�i3�J�2�U3���2fԡ3(r�2-"3\�'3sP�3�*3y�>3��2��D3+�
3�li3��3@D�2�3Wok3���3B�$3
I	3K!V3��83O3'�3�+3��-3�;3e�f3TQ3/�Q3��3b�b3�3X�Q3�03M*36�S3b�3��3�z3e�f3յ�3�7z3G3���2�@J3��2`3l��2m;�2W�q3)d3�,23z%33ԩ53�v�3���2�?;3ͽ3�3�:�2uj�2��03Z�
3`EM3y��3�23�x83_��2��]3q73�U�2D]j3���2#\X3��-3���3���2r��2d3%!�3Q-�3��33��#3�V�2s3¤3�\+3E��2T�3�� 4Ut~3��2�!�2��U3���3��3Î
3�7�2�T93|��2p%v3��H3�3=j�2��3��2�r3�%3�(3�&:2�3~��34��2��R3Kƫ3�v3#�X3���2�Y36W%3�2�2�-$3�S�2�y~3���2)�3`i/3~ˮ3��2H��3�(>3 
)3s��3��:3i��2��'3��'3[��2Q�Y30Ŵ3(��3�K3�3�a3Ƒ-3,�3�>3�4Z3�v3^N3q9�3��M3&il3�@3�)U3��U3*J�3�_e3�23͏�3�BV3�1�3�@]3 nR3���3��3:K 3�A!3�P�3���3y��3�ݧ3�OW3$^3�3;��3"�M3^�u3 �!3B$�3��3O/3sz_3ٰ�3��3��3��3X��2��V3#>�3�E�3*�3�Y3�y�3KnR3�31��3��3�Þ3��>3�3�`3ej~3��3�v�3!�3�_�3{{�3�<L3z|^3<�X3�`3�3���3��^3?�3�F39l3(9Y3~lh3�J�2��R3�T3#D�3�'H3��3�
*3�?3|�3CJ�3�H�3��$3:H3vY�3Y$3���2z�,3u��3�[�3W��3���3���3&��2Ca�3���3|�2#�`3��3�rh3�v:3*��3_3��h3�z�3��3>�3��o3��3���3r�-3��h3*��3v
�2�g30#�3#��3Ffq3�43�9*3ǿ�3(�C3��3=��2{Ad3Z(3~U3��3�H03���29��3+;3*�'3��@3��<3ϔ-3�G<3�ك3��3yQ�3��3�ю3�̎3�(>3 �w3�Fs3lIi3�Ӓ3Z��2Q�3i3P3S�3H�3zF3��r3��3��v3��X3!!�3٤b3�f3�9R3�eq3�63��]3~��3���3� z3%�2�j$3(1�3zg39z3(}o3Z��3&3�t�3D\3�'3K6U3>�4]��3�/w3I��3��386s3v��3�m�2�?%3�]�3�3cn�3;v[3�d,3w13���3��O3���32�K3��i3(X�3�ˎ3j�E3���2n.�3�9�2�J3�߂3|53Ҥ�2���3��3m��2hi�3�>n3}å3_��3��	3�3�3�ʐ3J43u�3z3j�3�.J3<�3d�^3���3��H36*�3��"3�30�G3��%3�<3s�3O	F3�:36�63���3Ծ�2�2�3���2�5�3ŭP3�)�2��3Q9^3.�b3���2r�Q3C��3JFc3f͌360�3�Rc3�I3��%3�`=3�j3��h3�$3EYe3��I3R�d3�3�3�93�@3֬$3��13b 3K,3p�k3F�3��J3�`3̀�3�c 3[�03Loy3-4K3+�2��O3�Cl3��<3�ZN3`�]3W�k3�ci3e+�3��3s�Q3���2
��3��|32M3}v%3�N3��Z3��2�ux3�O73o0�3SЂ3)�K3���2JI+3�-3Wmd3h�*3 w3�|3'��2�[3�L�3���3Q�3�C3�Ů3ȗ)3��2W��2�'3�[h3Q�3�$s3�^3�� 3�t43Z��3��3PF3A�3�	3LJ3��D3.��2�3U�>3|^i3�L�3�3]�w2���3�F3��35=y3��3JK%3n�83Xe3<]@3k3=3]�53�u�3<�@3��V3��T3��43U"3s^i3\fL3��2�3V�4<�3�)3��
3�Ӌ3І3#K-3yJ3�LZ3��T3�^3�U?3�)�3��-3���2j��3,!�2�13: �2~�2�=-3{)3��P3R�	3��&3S��3{A3��3�G#3u�&3��3B��2�NU3�c3s�.3t>3�vv3�G03���3��t3%��3��3�&@3!:83�K3��"3��U3�+d3���2�8c3�_�3%k�3}�3.3�i3�<�2|�&3<d3m��2_�T3!�2��3�`�2L�3w"-3��3�#%3: n3+'�3f�E3f9�3��)3:aa3e9!3��z3�1�3~��3 n_3�_�2�zp3�bG3�oA3V�~3�i�2�3(23�u�3��3q��25��2�#]3 [%3��E3��	3;�O3SE�2T3� !3�`�2��*3R��3�83�{3� 3�T3@
3'��2QXW3̰�2�9:35��2c�3�3{J�3��3��37]3��3���3�3\Wh3q��3z��3^#M3��3%�4i�3t�3��T3�c3洤3k�3'��3຅3��3��A3�2�3�A�3T�3e3~�41z]3b=�3\3��3B�3���397�3Y/3�7�3�:�3��3���3
G3���3κ�3��3�3-�e3CX�3!��3:P�3W�3���3�HT3��4ȕ�3�E�37j3���3�`�3��3�׫3��35��3R)4|��3]��3�3�3��3��h3f��3�l[3�a4!*=3l��3Ɩf34ϥ3�L3/;4bE3j]3��3��3��-3�^�3t��3��|3���31.54Q5�3O�3\��2�W�3���3ck3U��3�r(3��
4�J3ţ�3E��3�<�3Ÿ�3�� 4+ς3�e3��3~Ni3ܞ�3	F�3���3�>?3�v�3�z�3���3�3B13�P	4mg�3��q3��3~�V3Ӛ�3�G3�Ŷ3�y�3��3��\3��3���3i7�3��33 l3<H�3�ܨ3T6�3r�3�di3\�3,��3H��32�+3�4
�3ee�3�x�3SH3/>�3_a�3d��3���3� a3%�q3Ҁ14x�3k}�3N��3O�U3Tj�3�F�3�K�3cX�3���3�D�32m 4l]�3��3���3� �3D�P3{]�3�e]3���3`��3���3��3��73��t3z4��3�0�3؃�3j�z3滂3?��3m��3*��36d�3W	C4��3��l3z�3d��3a��3��x3�C�3�e3�5�3�I3b��3��3=�x3��3��$4�a�3��3Q��3�Ie32�3g6[3ARs3�=3rf�3"�3�m4o��3�8�2E^y3��4<	q3,J3�3 �3Zn3��3��3:m3�� 3��-4WIh3&��3 ?�32OT3*�:3I)�3��3}A�2A��3�,J4���3���3r�>3��43�3ˌS3A��3�3��3�jd3CU�3}�3u�*3y-3uΤ3U|�2��3Cw 3Q�"3�:3��X3�30qP3�B63�Yz33M)3*3�3�C3�})3ah�2��3r?3yVT3Ž�2�I3-�C3��C3���3_4ٍ�2��	3_(3v�3X�>3�l�3qȁ3��3	݂3��3��E3s83=i�2�g3oth3���2
�38�@3p'>3��e3j1�3Ql�3�i3Xmc3��3��2&6;3�13�fH3�03>�+3�K\3�93�І3bi�3*�~3��R3
5�2:�I3:�P3P��2��;3�3�W3�3�u�3?XK3�g33f/_3a4�3�.\3��O3|	-3�J�31k+3X73X�3f�3�Dw3�3�3�=3ZRN3�c3��^3�S�3�:o3�E3}	3�O3�"3�7�3��<3-�_3k��2A�3QlA3��:3=К3AW�2}�q3�n�3�RU3'�2��,3���3ӏL3��Q33�a3	�83c��2滄3΍3�|43ST3D��3��N3��#3}*3���3\�3�c3\93A��3Q~3�E3��c3��2p�3Z�3��3��(3dG'3F�>3�J@3��37�3|�3;�3��V3{*�3<�"3$��2��[3�ۗ3�;3)D	3�Ue3"��2@3Y+R3@ĥ3��#3l�3���3�S�3m� 3k>3��:3�D3,3x=_3��3��3�@%3�n�3,!3�D3}
U3*Y4�]3xPG3g�F3�� 3~=#3ysG3�~c3��2Bl/3��3}�3�lZ3�3Xh�3^�3�N+3�;3�A�2�b]3��3��3��"3ւ3h�23��3g.3���3tz?3�43[Es3�pw3�Bq36zq3�=V3�|3U�3¸Q3�,�2��3�a�3)F�3��G3���2B�=3]��2@�f3�X�3k��22V�2��3<qF3d3�?�3Zu.3O�03\43��3�.:3��3~9�3*w�3�'k3��2r�"3 ]�3B�83�$Y3��2TB\3�<'3<�w3o�3��3���2ܐU3�l�2�3!3��2�F�2��2�a�2Ԏ�2B$�2+��2�;37�2_��2��R2�3���2Iټ2�D�2Y�2	��2�jJ2� 3�43;N�2�T�2��H3i��2Cu3�3���2-�2��2��=3�@�2�A�2�pX3���2���2��x2k3�2|��2��2��2���2y�H2�Q3�l3�P�2/_3ik]3�3�2���2���2)�F3�_�2Q��2��+3��2ˉ�2T��3�f	3!A3��g2�?3�<�2��2w�3��2{�:3��2;4x3l�	3�\�2�L�2�ng3`Ka2�g�24�3���2D�2�V�2t�3���2̴�2�)�3k637��2��u2�3A]�2042�3'�2!�3���2Z�3�e�2崸2��
3jhV3!9�2<�2.��2��2�1�2)�3��43d�2�M�2�Jh3���2N�2?�E2.�3Z��2 z�2Y�2���2�H�2Mx31�&3L��2�3�82
P�3��3�33_�3��3�3-53���2��2x�2y�}3���2|�23͗2Fl�2<=3G��2�|�2V�2'�#3�E�2 533��3���2nGx2��K3o�2�h�2c�2���29ذ2�Z36��2���2M<�2ez\3��2S��2q�2.	�26�3���2O�N3�!�2�3���2B�3�`�2���2��53��3�`�2C��2y�2�۽2���2m3�M%3pٰ2.V3<'A3q�%3���2Ŏ�2���2���2��2�e37	|2�Z!3�/�2|,
3��3@��2Đ2FΎ3:�2{��2Gg�2��2U�w2��2��3��2(Lo3*�D31S�2�3V�2p+
3�}3�9�2;t�2��2�83봒2Ț�2�8�2��R2J�&2U3<��2
\�2�"3�z3lU�2Y�2�"3V�2���2�@�2��2�ٸ2O��2��3}x�2�qp203,��2`��2C4�2!�2�-3�?3I983�Ȗ3o�j3m�b3���3;�3�-33�3��3��h3['3(G�3���3i��3#3s�3��]3��)3��3ēV3��3�y3���3���3Ҹ�3��.3���3���34�38�3R3N�f3v�23�/i3
3���3\^�3���3�k}3�3mX!3���3A	A3�u3*�x3�3�0;3��3l�D3FĐ3"3�E�3�?g3��l3 9J3 ύ3��3UL3�c�34|�2�W3��3�[�3��3�=
3G�p3�r�3���2g�3�3�۬3HT3��3cSI3�!^3���3v�3V�d3vO�3��3bOF3��3�`3b�3?c3�ZN3�v4��3$�3W�2A�t3�Qu3��!3�4�3]n>3�7�3/.{3�4�3j�<3}ϋ3��13P�3Ke>3���3D��3��3y��35��3���3�53j/Z3�g�3�9�3��T3E>�2T�u3�_3t;3f6�3%��27�3�730D�3c,D3�h3�y3�k�3�G>3,?3_UN3�{3�|3x�J3��D3�3D:�30��3>�3\y3 �23T�3X��3 �3B�3��Q3ڡ�3H�h33�3�3��e3!�,3^�H4`�]3}�Z3:��3 ��3�O3DI�3&y�3ܕf3	��3��3�g�3vNM3�$3��3^3(37�3sx+3�63R::3�(�39�}3r]?3��3H �383h��3~��3���3�rK3+Ͷ3r͸3��3�/�3z4�3��3	&36(3
O�3�Ҕ3�N3�3�=:3�ٗ3YqH3�M�3�z�3�'3�yP3���3��=3�$f3A[�3Ҵc3�`s3/&[31��3^<3��c3�m�3�3:�x34�63�_o3]��3�`3&�A3,c33�Y�3g�83a�3��B3��23�dA3�K4�J>3�q�3���2��_3XZ3��33�`3��S31ٙ3�6�3b�3P�3'/3��3�3�t3�c�3I3�Z3��X3��3C^3S�3��3˸�3��M3�J$3�3y `3G�3�<#3��i3�j�3|�F3��3�>3�c 3(�3�	a3=�]3�O�2�{3�[�2/3�#�2�6�3��A3O�3lJ3ߩ4�73*�3�338��2��2���2�w
3'��3[�2�F�3�`@3��>3r��2�c23��*3
<3��@3��F3/� 3�E�2�@&3υ�2�8M33o�3��&3z�3Dr43Rt�3�O�2	3�@23��2F`�2,i�3�X3^z�2�&�2Ŋ`3�Q3��3(v3�(J3VC3��2�
r3y9+3�W�2.M�2�d4#�3�S83�S3�P3a
3�=3��C3�2*W3���3��$3qma3B�2n�}3%�3�-3$�z3c_*3�Q�3�>3E��3.�j3�[,31��2��%33��f3.F3h"3B�"3�o�3��!3�P3B�3o��3�>�3?��2HZ�2|CT3,!3?f3��3�-3�P3uI33�Ň3��m3>�w3��2H�3��H3!�j3 CX3:�3�#
3��3��3
3��P3�o�3�n�3�!�3)B3#�V3�5�3�]�2&�+3��93v�73�O
3��`3�73��3�,�27h�3@�n3��^3x�3^�2��53��y3�($3�~3�#K3iC3��38(3���2I=3�*J3�ڮ2�AX3� 3�!35cQ3�3?�3�<3f�3 ]f3��26�2�3�_3���2�
3�SR3v�2r�3���3�]�3!v�2��2�xe3:3Ú�2�3�0�2�3���2��Q3=�
3��3�JF3���3b�3��=3��3
�3>�[3b�3�t3��2ZT3,��3:9�3��83�n�2G|�2�4�3�h93�,3)0�2��;3�;3/c�3��:3#��2)�3߹4�#3Q)3�cY3`13�D3fa3p%3�P�2�+3���3�3N�2��2'q3_N*3s�3\�83AF3���3u/�2R:�3�BW3��3Z37	�3u37Z43J�2�X�3��"3���3��43x.3�h#3 �3��3��3�� 3g[�3��@3�W�2d�3��B3�s~3$"�2nx�3[nI3H�13�3t��3��	3�>#3��h3Q��3ԣ�33�3�33Ƴ3)�3wƔ3H�_3?�.3w:`3/b736A;3Ppl3"�@352�3���3�F�3�iy32O3��2��3��	3��63s�H3O�)3���2�+�2S�j3XF�2��2�c�3�\3�E$3S��2k�R3��d33#3s$F3�a3�-@3I��2��3�33�R"3U�$3�6�3�!3硃3��v3�za3�W3��3�J�3~�2|m.3�Yw3̇p3��Q3Z3�r>3��2X�k3�g3��W3�vi3,37O�32f73�B�2�X3�1�3Y:3��.3̔3��<3�8�3�h�3|O3�53�N-3
�L3��3�މ3�
3	�?3��T38��2׊J3a

3�3,�
3��3�#3��Y3(|)3�ӕ3L>3;_�3�`3��]3�3�3x�3�?3Ye�2�"13�L�3�¨333\3��/3��]3V�
3�Ly3;�I3;��3Y@_3�)z3��3�P3-�63\��3}�2�=/3���3�IS3�=/3��93r�3���2کX3#4Q��3*gX3B�3ʕ�31;]3k�3ĄE3�%3^�$3��3�f�3r 3�3� 3��3_�j3G�33�:3��3/i3O9�2*�3���2��3��3�xz3;X3��2"�3�RC3_E�2N23��13Tp*3��3$p�3:n3�av3�3\e�3t�3	ߎ3��37.3��43�&3dā3�I�2�`]3D��3��3���3�3jsh3��3�3�/Y3���2p]a3x8a3�p�3?�33�$3 \=3SL4��3'�3�3mC03�3!�`3g3��3
��3u;�3&�O3�l�3�D�2��3�	$3&�3�Xi3�.�2Ы�3�33�iD3
xv3!�3�:�3"�=3�e3V|,3�A3�N3B�Y3:�63B3&23Տ�3p �37m3uC3P��3}�H3���2��3��J3�M�3b��2+��3�3Lݔ3� �3%�3�.3D��3C'3�B3�73���3S$�3=�/3���3%JO30�3��3��2�3��(3
K 3�y>3�i�2&s93	?+3֦m3[��3(�3m�f3��3�l3H4.3�M,3�̈3�\�3R37��33��2�1b3�N�3���3�
3J�3H33�<3De3D3a^�3)��3�*3ݭ�3	B3Op"3�|E3�z�3�`3"�93��-3�wJ3l�235�@3�
�32ǧ2��P3�dt3�N�3
`3@��2��g3��30b3��)3.s3�1�3���29P�3!,3U�$3!�3Yh�3ي,3It<3X3�E3��e3>l{3i^�3��2{�k3�03��w36��2]�2?��3��73��2f��3�23vb3�s=3��3c·3W2R3��q3$1�3��3��3 ��3Aog3*�63ͿW3D)z3:�3�;�3�ǵ3���3�<3��2��3��g3�m�3�P632�3��n3NZ3�x�3w d3��E3F�$3�i�3�03k3�%3!�I3�j23�3Ӟ33{�36?S3�<�3Y8J3��I3��U3��,3�3 \3k�3��:3��35��2���3Q�s3�Y$30�K3�)4»W3W4&3�23t�3��33�S�3�D3���2'�	3�[�33�3hzq383H3�3�fZ3y
3�9O3Y�+3q[3�g3���31�h3�
3�d331Y�3���3%��3�ϊ3X?�3]{83��_3�{�3Z-3F��3U\�3�0�3E3P3� 3R�I3s;.3�3�I13ݑ�3�Yc3��3���3��`3�GB3&�#4y�3G�}3�	�2�%u3ʻM3��3D�3O�C3q �3!�3��3�(S32#3�K�30�3�3��34�-3v�U3�x3a��3e] 3��3�h3�ș3MJ3)�23��<3dM3�p3�T�3+�3%�:3��!3�3�#�3��t3��C3��3�wB3.�354�3$43o��3��3��S3O�r3���3M53�3M�$3U!3$�_33�Q3��	3*�)3��53���2)��3���3�`3#�\3-�2Bɓ3�A�3��434@Y3��'3�[?3���2R[�3�M3GHb3j�3�.�3S183�[r3�Y�3��3D0,3/��2│3��$3�`3D&�3S|3�C3j
3Q(D3XGG3�X�2�d3�t+3��N31��2y�3J�k3�03��3Ę�3���2�83�s�3�T3z�?3�"3��o3�(3�(%3��34�3]�b3ڽ3�6/3�R3](�3�"R3[�#3��@3)LB3���3�E3���2�#�2���3�33�ZV3@A3�[U3��T3��'3�8E3��3��=3��3HF3<Љ3.Ͱ2��`3��j3��23�6�37�B3�$3�C3�R3v��2j�3�E;3$��3T��2���3,��2}�E3	3PN3�/3��29Q3yl�3*��3�Y3��3�l�3`܋3��F3쭋3j|3���3P~3��3�S3+�M3�$,3f6�3Dt23<�3BUY3�s3PU�3~��3�/3Q63 �E3c{�3�%K3��3=S3Ye3t0�2� 3"&�3�߃3�MU3��+3ITU3e�V3׍U3w�s3�.4'x3(��3��K3B35#3[T�3E5/3(�(3��W3�3���3�MO3W.�2��3`g3x/3�5�3�$@3|�b3\j<3���3� 3�.3��M3�{�3�(�3�|�3~[3���3�b3�cz3���3�|�2�n{3�ճ3(H�3��D3�]3E��3�ky3)�3B�s3���2N�31\3S�3�SX3��3���2�_�3�s�2 �'3���3,c3�r�2��U3��3D3�Nb3cH3�ݨ39�m3�6�2�^3�38B13�93K�2��{3�Y�28�F3��^3���3?�3���3�bn3jd3�:3�G�3 G3��3ɱS3 ~3�{W3��3å~3p�R3�D3���3f�o3A�2��3{�f3�U3�3ߖ�3 �y3��3�+�3FQ�3�3o�k32[x3Lʖ3�3�;�3a=�38,3��332��3��3'�3�@3�1�3��%3�K3m��3��P3��3%3�ɵ3��]3�JE3u� 3U��3���3��@3*�@3}~3�>3�Y3��z34f3H�%3^N�3�}3r03$�21�3���3�$3"D�3]f/3��;3��3Fː3��&30wi3`�o3V��3K.�2ā3�L3�#3��U3;{l3g�3��2<�3+��3" �3xY23���2�!f3G�3��3�"\3�'3�3f''3>��3��3�3:�53-�4�L3]|!3.A3��)3�w3�`3��3���2��@3no3L3�3�;l3�43b?;3%�3�:�2ni3�΀3�br3RxP35�Z3n�z3� �3C,�3�C�3�W.38ۥ3�W�3 ,A3�T3-�k3^��3���23�a3�T�3B�3؃3��3i�3�B�3*ۄ3�T3�3��K3<�K3D��3�&�3�q.3(�l3V_4x�2�w-3>;-3�3l�	3(�q3�r3n��24�:3�-�3��3�{h3m�*3��3�U3�I*3Qҗ3�n3s&F3�g3�Cl3xA3�3��M3�=�3ǰH3k� 3��3ݻw3sȥ3�C_3�8a3�XE3U?w3x��3�S3�m73QC	3�%Z3�<3�3ך3�g�2�$3�[�2�A�3N�/3� 3zB�2��3��`3�T3"�3J3	�.3�*Q3��-3�E3�M�3���3�Q�3�N�3߽�2BvC3���3s'3�w�3��K3�X�3н
3�[�34�g3���2)�3��4xb3Ϻ�3�o�3�F/3�#3s��3[T3�5Z3�hX3��3��`30��3�3��y3_3�)-3�-u3�P�2,��3U�3	"t3Oʓ3`J�3úT3"A4,�O3S!3Ӆ3�5b3�I�2x�C3�9`3�S3��X3]��3�l*3��:3�53?�r3�f3�j�2�?3�M%3i��3���2�K�3�
D3\D�3nq*3�=�3�ԉ3��3��3Y��3�i3�z^3�~33U�+3�s4l��3~�3IY3��3��J3�Z�2�/@3>�43��3�r3�3h~�3!�2>�@3�x�3�9�2D�33t¤3��@3�9�3�K>3�MO3�t 3�V3�u?4P�3nBm3��2r�3��3���2~�E3��r3�)3�3G�4\ @3t��3T.�3	4�.3�8�3h��3�P3s�3~��3��483d�3���3Z��3��p39�3.E�3F�3d�i3�N�3 �3�\�3���3~�3Eщ3�b3i��2�3�0M34%`3��3�P3z�3��3�$�3*"l3��3�5�3V�3�g3��3,��3�ŷ3�Y?3?��3#n$3:�3�d3d�3��&3�039	39��3�3�JJ3O�4ڸ�3ʆp3��\3���3��73��E3��3'L}3tǀ3+%33�3�"b3ָ3�%x3�S.3"h3�2P3�[3昘3�k�3HLa3�4��3Nr�3_53&��3>j�3���3�j�3`�a3�l�3s5�3�\3,X�38�3w,�3V2^3��$3���3j3I,�3�~�2���3�$�3��@3&��3A.�3'k3�+3��W3��3�N3�~O3��3��V3O�53��3�ͩ3#'b3��3�)g3��3R/3��3��53�	13c?]3��3Ǳ3v�3�zD3.�4��~3�NK3�3@�@3�.3��-3|�3�r3��3�#�35�3l=3��2tU3��f3-��3)��3�>E3�}�3��&3�:4[Pc30h3��3&�4VV3�;�3�mp3k��3S}3]�S39R]3s93GC�3�S�3�4c3 P�3�'�2��&3'��3z��2��3ڑM3x`_3W�63��3��O3�3�Z53�j3I�{3��3"8*3��E3B�3HG4�a93xnR3�%03R�3bC�3@�3�5,3�Ko3o53h�3��h3��:3+" 3��j3�m�3��3��j3HS33�3�Lp3g3��X3\e3)
4g�d3�2�3OS�3�7�3�}�3��~3X��3�*N31��3��M3�3�@3��~3;+�3B��3R��3y�3�N'3}�3%I�3'�23@03s��2��j3_c3�LH36r]37�3y}63��3�	b3%�_3Y�2,�_3:�3�q
3ѾB3�l�3��Z3{��2�U3=f�2sQ83`83�*�3<��3}3�ȁ35473�m3v�-3��3�3��93��3Yho3��D3���2��%3mE^3��P3V�"3�=q3eq�3c�2p�3X�I3(�-3X��2r�3�Q�3��3�3��;3O`B3���3�c3_�2�|h36�3���3;;[3y,�2�ߕ3d�R3D��2�%O3���2�33�>53N;�3�Yg3�33�{d3	�4��3�l3]��3���3�P�3�b�3��3hf%3�uv3N��3s�3�J�3�Jn3x��3A�3o�3�J{3(3�<83�$3�Q�3��"3ЈX3F�3��3�[f3ך�3+{t3ah3ӎP3s�e3���3A�3
Z3~�4(�;3��<3�D3R�*3��23�3�7�3�$3^d3� -3�[�3��S3Eg�3^�3�4Xu3�sv3�'3K�63,�b3@/�3���3��3wuG3.�3E6�3oU�2Tz�2��3h�3�93}�t3q~3��3l 32��3�%d3��2��H3��4��r3�[Y3��<3��E3h�E3o�V35y3=03�.3rͷ3^Q�3��3Ů+35vJ3��3ҍ/3:+�3���2?�3��3��3DӉ3آ3��3.�24tw\3��d3��3�3�KV3!�:3ڝ�3�3عt3���3a��3L�03�|3G�3/3��3�l�3���2�s3.�13��3@3N�3{�W3���3�b[3,�23��G3�S�3���2'�{3_y�30�22T3���3v�[3Ӵ3Ԗ;3}ہ3r?3�
93�'3��3�Y3��2�,�3�\3p�3O �3��3Ջ=3��3w�s3O93���36י3���30��3
u3�U�3���3q�>3T�3��3! p3�3� �3�b�3|��3N�M3�_�3.��3�VX3��I3�L4~@G33@�_3� �3��.3�b�3=]�3���3=�q3�z4�<�3��l3G�2@��3+?y3^\3��t3!q�3�æ3�`O3n�3�6�3��83{�}3%64�]�38\�3�k�3;̀3�u�3���3&*�3h��2�)�3�`�3W��3c��3I83K3���3-��2E�Y3�d3ֶj3�Ք3lS�3D+�3hY3Neh3�*4�=g3'�_3��A32J.3Є3)'h3�k3a��3�0v3�4�{�39|3I�O3�ޅ3x`�3XG_3�%�33w{�3��A3vr�3�u3,��3��3p�4��3W��3g.3i�3�Bs3#�3�X�3	k�3�TO3=4�E�3;F3�3��3&̒3��3���2�23��3�3�j�3G�3��G3�?r3k�41	#3�:3�3�|l3��T3i/c3O�3{�3�_3a4{��3��|3N�:3��[3�u3cQ�3�uN3>�2΀�3��(3��3��O3d��3�K3#4��3N�3*҈3x��3V3y�3I�3Nt33�h3v��3~g�3�� 4�d93�}�3�,A3]E3��=3�3�e�3�U3�ƹ3��3��3�53�^46ѐ3�0�3Ǌ�3�d�3��3݂3\�d3b�I3���3���3�'4>��3��(3P�3�v�3H��33�#�2�uK3���3�Q3kY3��73��2��3��3]%�3�G4_̮3Eu3o]J3Щ3҃�2Tw�3�r4��3ِ�3L��2T�3��3,_3n�3M��2M��3fO)3�V�3��53E�3�_3z4��37��33Pĸ3>E<3t�3-A�3
z3��3�B+4%�4���3���3%�3oH�3EHL3 �3��3Y�3ɨG3�4�4���3� 4�A$4]�3�V�3o@�3�y!4��3�	4VZ	4r��3�>4��3��3��3�,d3AH�3���3~93̾�3�s3L|4�Ջ3�#54Fۼ3Y��3�3��/4�Ѷ3�d�3O#4���3�B�30�3k��3��3��3��'4S��3
��3b8>3�̾3�A�3�#3f�4��4��3y�}3�44+Н3�U�3餵3	F�4͙�3j{�3���3�?�3C_Q3�)-4~�3�N3�Pk3�)Z4��3fĥ3k�X3qA4���3_�q3�n�3�Ӯ3ӑ�3J�83ŤS4�ټ3���3Y�3B�	4�l4���3}��3� �3-r�3�"v4���36)T3�3��3�(�3!ܢ3PVp3g�*4y�3u�H3��54�3�"�3R��3��H4F��3y�3�S4J�84�O�3�a�3�f�3�	4萏3L�3�t�3�6L3��3:�36��3�ɕ3��3O4krM4���3�m�3D%�3P]�3m\�3�o�3+&�3�3گ�3�|{4q�3.��3���3t��3���3���3���337�3���3�,4��3���3xDf3�<4�[3䎊3{(4���3��3՝�3�2N4��3�
�3�R�3��q41H.3M�3�;c3<T�3��3���3+y4 ��3���3�w<4���3�~>4-p�3�v�3���3�֝3���3:p�3�W41�3!4g�3z��3Á3�AL4OΎ3��3��3+��3�/�342�3O��3��3R�39�`4���3��*4�ߗ3܎3���3#�3�q�3�\j3Ԓ%4E��3��3o�3�SI3�3a5�4�"�3app3��3TMp3O�63e��3�[4uN�3��3;�3i�3�]�3��D3_�3Ũ�3V��3N��34Σ3��39�3�g�3�#�3#N�3R*3�פ3g�3�A3�}`3��3؞3_3a3ϧr3K�+3��2<:�3�Sx3�.�3�
3��3=��3k�333�Q3L�&3���3��
3��3�0"3�p�3�x�3��3�*-3A�93���2P$63��3��2@�53QV�2Eƃ3T9�3!9h3��3�z�2��B3�)3�O3k�3��'3�/U3?;�2��3�43��3�Z3��4�;&3�"3��Y3&�3�|3�:@3|�,3i�3�5�3�E�3�39)3�b�2�G3ʜ3.��2DF3a�2RP3�q30�3�5E3MW3v�03c7�3Y13T�35Be3
�03� 3T3��J3F�3��{3���3�>z3���2�6�2{+r3�`43&:	3!�3�3�SV3��3Bg]3e3�%!3a 3�A 4�r37E3�{3��t3U3\@�3S�$3��2��C3;��3T)x3��s3��2zQ`3{�2��3�U�30c+3�(a3Q$3a̿3�R�3��3"�J3w�4��d3�/63�=3#/39��2WK33�13a��2xO'3
<�3��3��z3�3=np3p;3�3�+�3�I,3%��3�b93���3�T)3H7Q3_9A3�/�3�!3�`�3�J/3�e3v߃3	�3�l3t43�0g3eΧ3�ni3��2��03.c]3���2��3mEo3$)3C�3��"3��3��k3doS3uT53i{�3� 3��735��320q3mE3�A;3�Ӗ3�?�2��^3N�3/�S3��f3P3R0J3!��3��.3���3��O3�U3��3Q��3=�%3���28{3��4M��2��3$}39�33$N*3L-�2�K3�5'3wd�3}\3?jP3�or3�x3��:3�b3� Z3�z+3��33YEp3�135�3h�m3g�'3�T�2�C-4#}�2<`3�� 3ׂ�2���2~�"3��O3Ye3��c3]3!g]3ǁ3��2��3�,3�.3U�d3!��2�d�3ߒ3��3/:3�a3��3���3Z�03��13��3��h3f�	3kͧ3+3}3��h3���3��3�S�3��x3{i43ߊ�3��3�Q�2mlR359�3^�W3�3��3��3��3�w�3l�4�L`3Ds�3׆�3�]�3O3rZ�3a�g3
c3i>�3��3��p3ཱྀ32/3���3�R33��W3���3��~3�ki3���3���3t�3��`3qǨ3���3V3P�3
�D3m��3p�3w�73�.93��3k��3�f�3���3��3T��2;�23��w3��R3�I3�Z�3 �3��3W�3>T3�U	3<#73.��3&*q3�ք3��3軴3�@�3u�|3�t�3t�2C��3��3��3� t3��2��y3���3f3%3�B3�_�2��3�H3��{3cQ3��13I<3d�4u�3�8h3�H%3�O]3�%W3Q*�3L>3�03��&3���3�IY3WU�3��'33��3O8�3W�3�Χ3��J3�vn3!�3� 4��3��2*%�3���3���2*f3-�V3;�73XK�3�3�3�)39̵37s�3mT�3��c3�d�2���3��3�\_3���3�[�2ｆ3o��3��4�9.3�13 �$3�2^4U�/3�y37
�3�vr3Lb3�d�3H^3(|o31��3##4�]3�ź3�3 � 3�>f3<f<3J��3�*b3=�3�_r3�q�3�3	3">�2�n4�fR31O�3�3|�a3��H3�-�3�ߊ3& 3$Ã3��31̓3�3�^"3L��3�t83�h"3.��3�3#Ba3J-e3��3��G3�T3��3�$�3��53}�b3��o3?L�3��^3�5g3"k3X�&3��J3�?�3�	�3�ߏ3�c3��3��3�e3��?3C�q3%�`3@=3���3�I|3l43n�N3:�4���2	�3�U3^3�U�2y&3�m]3Ed38n�3m��3�de3gǛ3�3O�30�q3tjl3� �3�3��3�U3��3a#m3��3TI3�3V"33��
3(<3TA�2b�n3�|;3�?3v�3�5�3A�137a3��28�r3n��2��2�-�2�-3eo3+��2(
?3Y�,3K�G3��b3��f3�'3{�2��Q3�'O3��2�?3B�^3��2]�R3d��3�^3�3̡�2Y��3I�@3��3��Q38��2��2��3��e3��!3��3N�3J�3�@3�&3�c3&%�3��2���2=��3yz3Z�3cP�3��l3�Q�2 ��2\�.3BZ*3:��2=e63��!3��3�2�k3�
3+�3�n�2��q3 ��2�3���2�y'3|�2d3��3$/�2L�3nm3,?P3��;3\��2�X3��3^:3��+30�:3�3��2��3%3�2�� 3J�3;a�3�ϡ2��83=��2<!�2*��2q2P3jM3�43�zB3�k�3��f3g�3�� 3�!X3��>3�53�(p3V�L3�;�2�l�2pܝ3��2�;3@�;3�3��3��3���2a�3H��2��33�,3�[3
�3\zj3�53�^?3���2��j3Wi�3R�2}�+3V
�2�W.3���2��3���2��x3˻�2n�3nZ�2��.3!�B3�3�N�2�3�K3�3Yb340�3�K3�"3j�2��e3Q�>3cb3+e.3��3b@�2�a3�^�3��3��
3M{3�3$3(�2(3��E3 (3�|�2�3��c3v��2��%3��G3�`53��L36�3�C�3�GD3���2��m3��2F�V3>��2'N�3��03N3K��2s3�?3%��3�[-3"a3@�R3ST"3Ʌ�2�<�2�m13$~3,[�3�n=3_-�2l)3̘N3���2cVT3)�2�3*�3u�N3��H3#q�2�<3=u�3Ǟ�2Um
3h�K3@3$ל2D^3��93���2 �a3O�3d�3��3ȳ�2�]v3��E3�	3a(=3b��2�u3Ҥ2��x3��R3��3`�3��4��3jf�3/�3��3-�3א3�{}3o:�3)K3px4CQU3�Y�3*�3�3$�Y3�(�2k�3�J�3R�<3��93QM�37U�3j�,3�_m3�ٙ3F>3+��3M$#3|d�3Wד36�3���3�|"3<~!3@��3�̧3���3��c3J��3��Y3	b3�D3�kf3?�!3��3<j�34ٌ3+VK3+U)3�"4X:3��D3>�'3��g3e��3�c�3f�3�Hn3�^\3>��3�֑3[3P�13F��3q153�NV3(3u23�3�� 3��4rW�3+AF3�;03��3�93��3
Q�3.|B3���3re�2�ځ3Ƥ'3��H3?W�3KA�3`��2�g3�Q3�S3F�93�ѡ3®V3�L3V}:3Sb�3�	[3�23 �F3p��3�c3wD�3C3'��3mA3.gG3�݆3*�$3�8r3�	�3y��3�3a$!3�|�324b3g �3b�P3�C3��J3�dp3��\3X��3��3mYW3g��3xPK3V�3��E3.��3\�R3��-3Ѕl3��2.n�3�	4�\�3�Z3�� 3xE23�3\�F3�+y3��(3���3�:3lT�3#�3�؇3���2j��3��v3��3h�V3�&3%�3Ucn3%t�3��j38�]3,��3�?�30.,3��2[�3teE3N%3t�3��h3:�?3�TA3��3��R3�8�3�32�4��]3�d3놅3^>�3-F3�H�3V(�3��%3�Q�3�*�3B�3�o3�13���3>��32ċ3(��3O�X3�3=d�3	)�3ܕe3Oz`3�Y3z��3��e3&��3<ʔ3b�{3G��3���3�0q3y�N3�~3���3{��3�:�3��53���3�3�x3K�3��>3Cj�3�13�� 4�T�3�
3�0�2��4]�3BF3�ܪ3��t3��(3��k3|o�3�43�N3f��3F�J3}(�3f'�2��t3n|3�w�2��3��3���38�B3=�3�13�4�3��X3i�4�ç2H>3<� 3[�3+�J3���3�Y3Fn3�/�3�=�3c431>�3A!73#d�3�[3t 3�ы3#�63�SW3��3�@�3��r3�3�4�3�}p3�,3��39�w3��3�T3��R3��3�[�2)��3,C�3��3�� 3`#3�q3�ym38r/3�)53��3�{3"nS3�s3��+3��3��g3�c�3r'~3�s|3��+3<CF3���2�BI3��3u~'3ʺ�3/&�34(3��53�E3���3�eS3�]3�&b3o_3k�3!�3�
4wY3��q3��T3�
�3�cK3�f^3�p3v/l3��s3 ��3о3��3�3���3Vp3�WO3sP$3���3I�3�^33�X�3�0�2�˴3s�3�J�3���3ouN3V�3� 4֬63�3�%3�o3?u�3��30(�33a3�6�3<|�39of3�oN3_߈3܂�3I
93�I=39-�3� 33�&M3��*3MFx3�
�3��,3���3{3�	�3�:�3��3.�)3V��3O<�3��3��\3�9�3�,�3� 73.)3��3tN�3��2���3U])3�C�3A^3�ߊ3�?E3�w'3��%3K8�3���3�y~3a��3�`3[ǲ35<>3h��3��T3#��3W��3��x3L��3�$3��3RN�3�u3"�L3�ɂ3��3Y3�\�3�)�3un3s�)3���3�H3�h3�m/3�ns3+o31��3��3�h�2P�3�*�3�sz3�ޤ3��)3{�3�j�3u|31/�3w�3f��3��z3^�3|T3�3��3A43rn3�D3�w3�UY3�B3�q!3��3K3�El3)?�3}��3��3[�.3��L3��3��3���3�z(3x�c3�#3�13�a3&T�2mQN3�4�3�{3�~�3�c�3?ϰ3>ڞ3��A3G�m3�O3��3�N�3�Q�3�bv3�D�2��k35�M3��;3þ23c�S3b�w3�(3��3b	G3��3�2���3�e3=3��>3�%3�23#��3�!^3!�83!3	�3�j3P�3]8<3I,�3�6`3ܚ�2�mM3�3N��3#:/3���3�H!3VЙ3�W�3�P�3���3�D73Z�I3_�3c��3M13�[�3#�C3[
f3%G�3j_�3��B37�g3�R�3��3�v�3��w3���3¦3��e3R�R3��33��F3מ)3x��3�3�6C3�U3��c3��O3P�	3��Y3��2��g3Z��3� 3�	�2���2��3�z^3��	3��W3=^3픲3�ח2��3/�A3;f�3��2<�4Eu3͟3��3�{3��2�|3�C�3��2��H3&�3y:3��93�� 3`�e3�� 3�W�2>̅3��63��N3���2�h�33xh3;��3���2�+�3m3��w3��53��I3~�r36x�3�m3��&3��i3��3*83��W3�V3"{�3l"3�=<3g��3ca43��23]�f3���3��3�/3+o30s4L�Z3/?3c3��>3�3#=�3��R3>263��3 �3�0�3�5�2��)3�t3:aB3��3a�3�"'39�83�3���3�@3��/3/�3��
4��+3�o�3:8M3��`3�38�o3�]3�3#3��r3�|�3�l�3�L=3UH3��3�nC3y\3��3�s	33h3^$3���3��A3��3�LV3��3�zD3/�3�3��$3qS�2�� 39�3���2��p3�-4;ԇ3�L�2�<3��o3 E3 e3/�3Ic#3��3]3�=�3B�83�d36��2U4x�38 w3V��3;{3�� 3y�3KG'363��}3��o3n�R3��3a��2�ֈ3�|O3b۟2���3B_�2���3;K=3�E3��E3Lj�2B�K3��4�X3@A/3*�)3Tk3��k3�o3���3cy13��d3��G3bOj3Ĝr3ث�2T�`3�^D3&�3�{3Z�2�|3�!3��y3-D436F�3��3���3�w3�S�3̮3�3o��2�(�3Эj3��3�J37	�3V=�3�
�3�K3��g3�!o3�C3M�3^��3��a3ƀ�2gԟ3�r3��3̅�3���3�3'3��X3��3�M�3D�[3Wߦ3㐑3b|p3 P3��3MW{3��3��(3�3"O<3��53��3�+$3ጏ3Tu�3_��3�b3{�-3�
3���3L3pqe3���3�h�3�u3�o3�nJ3�x3r��3��3��34�p3|� 3 ��36�!3KS�2��3!@3^D�3J��3��3��F3�<�3��3���3d�d3�O+3�"s3�H.3ռo3.�j3���3J @3�&�3�4K��3��I3��3Y�3�z3��3�É3>>3�F�3/n3��3xua3�13*��3ň4"�)3��	3sMj3���3S�F3��O3g]3O573{Ѝ3S�4D̴3-�3�X35,�3q@N3��2��H3l�-3�{3я�3��3��<3�KY3xT=3P4��}3jxC3��T3�d3d503�RJ3 M�3b?�2�VR3��3�;�3Л93v*D3���3~�~3�Z%3�G3�3=�3��U3Y�3~r3�rl30�3�� 4�\�3�)3Lmg3�J3G%�3q�-3M��3�|3 ܑ3�E*43�3QP�3*H�2���3�g�3*>�3]�3'aC36�Q3gZ3$�4��e3�E3?�S3(C4^��3�iJ3)��3�̘3GW3�FB3v��3�33��W3[��3��3.��3���2W��32:�3fF3v�3~�93�0�3	�t3��3�.F3���2yE�2��3G�.3{W3��53�13�K?3t��3g��3y]_3�*Z3sϺ3���3�b33�03��3��l3nz�3�w�3�DZ3���3<wX3+P�3��V3_�#3��A3]i<4=l33�\i3��/3�ӄ3~3��39Q�3�"'3h�3b��3�Ĵ3L�M3Ԥ�2��?3�`"3���2���3�2Cэ3�b�2��I3�2�3���3���3�4'�3�\q3��S3\4X3�93O�3��Z3k�3Eq�3��G4�V3�3�3ۙv3ъ�3�R3��3�23C��3��3�<3F�3f��3<��3m��3lr?4/Z>3�)�3�v�3X/�3;�B3eA�3�
�3� �3I��3?��3��3���3َ>3�
�3�|3��C3zu�3�D3��3�� 3��3���3�9�3��~3���3�o�3���3��~3��p3T-v3��3F��3ˤ�3��(3�?4�N�35Yf3��?36��3��g3m7+3��3��q3�n�3���3���3��3�Ҟ3f;�3�L4rv�3�ۇ3pZ 4��3�2J3�<3��3w�*3(��3��4N}�3v��3QÊ3V#l3�4L�3��3�3S�3�Y3��3?v3p,3�<3��43gk�3�Tp3�V�3�a&3�3��3�83+��3W)�3�h�3kaD3,��2��3}
�393{��3��f3��38;3��3*si3=�3��73!n�3���3̠�3���3�Hx3��3�ߊ3��3�*3-3�4��3̤4{��3~ 4��3�n�3\��3Ff=3���3�R3F��3p�3���2�B-3�j4���3��3d�[3�j3B�3"h�34��3KM3t^�3�2�3,?�3IL�3б\3��3�a�3)C3�g�3��3���3��3��3O>Y3rs�3���2�\4�3	��3�7�3cݧ3�[F3�*�3÷�3�Fe3MX�3U�3��3\5{3�Q]3��30��3fN:3��3#ǆ3h�3S�E3��3m��3_��3�+�3�M�3u;�3�|�3X4�P�3r�3�o3<j�3}|�3_��3i�[4��4��Y3h�I33��3�L�3¦�3���3��3���3�M�3Q454LШ3��R3�b�3�5�4I1�3���3�m3;�34s3λ�3�4�3 �'35��3
��3�"�3m�4ő3�ci3�O�3��3 q�3��&3=�4W�3��3}�]3Byp3�l�2�i3O3�3�93[ 3�� 3o�,3b�<3�,3*VR3)��3Ht3� M3�73�/b3J�a3GV�2��37 �2�B3��3-�x3�g�3�,!3߱{3@�4��63��$3�r3���3g=%3�p3�O73��3_4�3�3vR�3�1R3!3V|F3��'3��2�093��3�NO3:�73��3'*3�s63�h�2
�4
}Z3n�3+{c3W�3y%3�;3�}3t(�2B&3���3&�3=	Q3��23��J3Z�93
f3_am3|��2�q3��"3|�3�m�3n�3�Z3d�49*E3�pY3:*Q3�n34��2��~3��%3���2��3C�4�)g3�:3c�2(�B3F�33}��2�u3�0&38Q�3e�3���3w&3��q3�t3i�3���2�<�2).I3-�3�)G3��3˭x3�°2�=3��S3��q3MF/38W;3B�V3Z#J3�h36fI3Nu�2L�Z3��*3j��3aD3�}\3�3�
�3�H(3��>39<~3v^g3i��2`O23ՏI3�."3ܞF3�ۛ3�E}3�)3S��2�In3�g3c�O3�{03���2�eA3�
3�B?3 �3���2��3q�32�)3q!p3]�*3d�3A3��93��E3L,3E�e3�ʛ3��t3�*31��2z֜3�r3�wA3��3��3X]3��P3XK�3��	3h3�^3�X�3�R$3��O3B33��I3L�(3��3��Q30�
3^�J3��3Hb�3w_3$�2�k�326d3��f3m�3=�23IŒ3��3<l�3�rl3��!35�E3_	�3�&3��h3cp36-F3	Ԅ3�D(3sKu3hK34�$3ui�3ܟ�3؟G3r�3��3Y�3V�h3�tJ3���2m�y37D�3�.3 ��2?�2�3:��3z3�C;3��3u�&3v�	3���3B��3ݹ3��	3_��3Ie"3@�a3M�3�Z|3�r3kl3�3W��2�J�3k��2T�t3�'s3��L3z��2�@�3\�2�53
�3+�3	��2oj�2�3o3+�3�3`��3�&�3�kQ3�k3��S3F��2��2�_3�f�2%{3��2^�3��e3ٍD3`�3M7�3"�!3tI#3�q�3^ى3��3��P38+u3�e�2��+3���3�#o3�hN3���2�]3�3'��20�3��(3��T3��3;U�3��_3M�@3I�P3z��3�H3bL=35�!3GrV3g#3�{�2L	G3�[�2�C�2��3]�3ß$3�M�2 �31w3�$�2��@3KԿ2	�b3�2/v�3��3��3A�M3��363���2��3zU�2��3A�t3+�3�&3�Nu39؆3|D`3|x3��3�63J&3P�3��z3�I)3�͇3�S�2��3�#3/�3�UE3X�4+uh3��
3k�3�<3s�x3u�3�3N3
�C3-'�3��3��3�&3��3�>3��3�)3=43�(3K>A3.��3���3�V�3��3�3�b�3���2��t3�[3�B#3��2���2k��3�\�2��f3�Y�3�S�3�,43V�3t K3"��3��E3]L373�+�3��"3"R�3{533�3�ĺ2���3 5e3�f)3Py3�Y3cVX3>-3���37� 3u��3��I3�f�3��M3��27�j3Ü-3[v!3adv3��03�#W3_�3%��3��u3��2�u	3�.�32BM33��%3�!i3�3�r�3LH,3�s#3���2٠�3�!y3Ʈ'3u�2��34�h3h3�2�6a3dj�2z13���2P��3%�/3Z��3���3 P}35]3	��2�/C3J��3ľA3o�g3�y�3��-3�_3z�}3�i3д3}�B3��=3��<3� 3�}�3ӯ\3�3�3���2c�m35�3��3�0�2]K�3���20R3�ޟ3�\13��39R3b-X3Y[�2Y��3s̳3*R�3�9i3Z8�2��|3)6.3G�=3H*3�
3s͌3&�2WɄ3��S3I3-3e� 3Zgg3/3w#3��2{�\3M�3e3�G:3�G�2ؼ�2*�\3�l�3�?>3	��2q�3n�E3!#�2��33�/3��@3Nj�2 �[3z�:3�b3Rab3��3���2֏P3�`43ʲ�3��3d�*3n�.3��+3�H3��{3�9�3�W3$B&3�E�3�}3Ԏ3�%B3�V3̬3#$3� ^3�F�3(�43��)3��3�	3�n�2�?t3��53L�2�*�3�(�3'	3��]3��l3�833�Z�2��(3d�'3/H3``�2��3ʴ3�J33�z�3I3�3��3�z�3�a3q�S3,-03]��2��!3�<3l&3�Ŋ2��3�ob3�1_3
�2���2�J37P�2�3��3��3��3�Z3���3
^�2��3{��38^�3��,3`3�9S3�203��3�E(3
�3��$3گ�3-��3�T�3��U31�2��3@`]3.<�2.�3�'�2��s3~_3�'`3y}3�T3�B
3�ܤ3���2�Q�2�SU3�DB3��
31�!3n�93�w�2�N?3�!;3Ah3�@3l�2��3b�3���2�
"3�?3:\83�:>3�Z3k��2m &3�1@3�]3;E�2k	3e�s3�/�2'�z3Ǔ|3sB3��2?\�2�˚3�
�3s-F3Y`3�ؔ3"�3�N3�zI3�`*3�3`DC3 �3���2l�E3xn'3�u�3��3��3ޒ:33O3J�K3t�-3��73q	3�R'3��	4*��3��3�Q�2	�(3Ջi3P3H�I3���2�s-3��13Tp�3�o3?�2�3T��3l�R3��3�73��2ٚ53�3�cM3�3��!3x��3Mͬ3G�/3���2�w�2��3��?3���3A��2e\3O�43�a63k�3�ު2н23\U�3}Yo3��2�a�3W30!_3�$:3�mm3�s�2l�3�O3�>�3��z3fV�2̾3Ap3,�730m�2�%3�3�M!3q9�3�[3*36�43�&c3��3�"3;@3��#3�"&3B�%3��3��2ٖ�2��P3�`3��I3���2�r+3��3JN 3j4�2@��2�>3B��2�3�Cd3F�3��2i�3���2h[3��=3m�3�33�3��O30W3�Q-3�+b3�F3/�2 3��]3|3sG3c�2 �3��3	r3xn63Č�2�p�2�c�3)3�03c33���2QU�2#�'3쯲2�d3��Z3�,M3�=3�g�2;�2�.3`U�2��.3j�33K-3��3�W_3�p"3�"3��633��3U?�2��2L�$3�}03K��2x�34<Z3�sr2�a.3g�c3�,3�"3b��2A�2�I3���2�W�2��3�g,3ޝ�2g��3��2Uz 3k.�2�Xr3�2E��2�b3���2S�2OjP3�/�2�n�2��.3�3\�3�.3���2 *3��43��2�b3��2��2�f3�)3P�3�3I1�2n+�3=�2��3�3<73G�3��33�3��a2�$3��3��i3v3R3yY&3_�:3 �3fq�29�3:z�2���2�h*3`��2�A&3���2Ԯ3���2��/3���2]�3�\3.#3}w43۰3�3���3���3(^3�2X2�2�)�23�2�(�2Ya�2�#038@5363ꈵ2n��2��3��h3��2��3��I3Ù43:��2�f03X�'3~}�2f�[3r��3�|93p��2�9�2�d3�V�2�ݖ2�I3Ϭ�2#��2���2�o]3��,3���2\g3�V�3�3�34�2��2��/3�:�2<��2�Z�2�73�؍3��y3�&�2��2|��2,�83�x�2��2�,�27�?3\�2� A3�b�2#�2? u2�E�3�L3��2�J3�3]|�2�8�2wk#3�lx2z��2�J3�3��D3���2EU#3�I3���2��
3���23S��2��V35�3���3��t3�4�w�3nͷ3a��31��3�E3%��31��3�Í3l�3mj48�3�ɨ3^Ԝ3���3!�3�ڼ3W:Z3���3��4g&3��4���3?�3�Ze3;��3�E�3�Ղ3�S�3���3O�3'\�3���3�K3���3``#4���3��3i�N3���3q�3�I�3�4�3�I03�]�3f��3�ݼ3O3��3F��3�M4��=3�)�3�J�3��3��3�c�3!�3�*�3�R�3
8+473�3���3�E.3���3�p�3o~O3�t�3���3T�3���3�3ɇ�3�x�3@��36�54Ԑ3S�3��53{ �3�H�3��3B7�3*n3n��3z�3a�3ڧ�3��13.$�3�zf3|`�3j$4YJ�3���3U�f3�-�3���3y��3ff53�64�(�3�zU3���3Ƹ�3GG�3��h3���3,��3���34h4X<d3�s3�4�ƿ3/��3ʖ�3�m�3��3 3�4Ϙ�3���3�z�3@�=4<F�3V��3�/[3V�3"�s3u�3���3�A\3��{3�w�3���3�N�3�D3��3P��3)�23h�3$BU3[�3d3���3	V�3kO�3N3��o4V��3���3�p^3��34t�3���3��3�[�30ܹ3�4�ќ3�i3�*�3[�3��r3VZY3�K�32dR3�!�3dC3��	4�<3�˝3�4�3�]4��h3���3�J�3kP�3TG3-ߺ3�04aF@3��|3�3�B4b��3�gm3�,�3���3�;�3�4�Nd3%
�3��3o��3���3�ě3vp3�;[4��3���3W��3L]�3�h�3l��3���3b�p3���3�)�3��V3`!�3�ɷ3�^3��3 ��3H�3�cs3�Y�3 53��4��3#�:3^�'3���3�p�3R�3Zp4�|�3(Щ3+��3.I�3��&3?��3�_�3��E4���3��3q�4��3t��3��
4[2�3+m�3�Kh3T2(4���3�e3F�63j�3Q�l3��C3�y3�S 3���2M�%3K�3Ӻ3�|:3�ӕ3�!3�$3W��2�4,3�@3B�3�	3�e3�$3t�2:��3��H3ä"3J+3O��3��3��W3�8`3+�3�3<�L3�cO3��t3�?3��"3̪3� 3�w3BZG3n�&31+�2�f=3kA3,�?3^��2���35e�3�.3:�Y35v�3��P3��3͇3��-3�;3�3��3�U�2��'3�h�3ZV�3�� 3�d�2yy)3�3B3D(�3��2lZ3��3_�g3{73���3� �2�^�3�}>3�[3,E(3�EC3��2�z�2��3➉2�n3���3{�_3��3��2F�i3�93t�3υ+3��3,��3��2�93�*;35q'3FE#3Rx�3�)3(3`�3bB�2d83�a3!�y3��)3D��3?_�3Q~3aw3�$3�k�3i�43�D,3\�3@133�3X#3�"k3�'3AKG37I(3�א3F�3!�93�E3"�3�;3Lgz3�3��2��D3�,�3���35�P3�F 3�FZ3��p3y�2[	63(�2U�u3�<3�m�3v 3 �3��2���3g�3|j3\q<3F�H3'�U3e�3'.�34�m3���3e��3/�3}�2��2@G3�VV3y=63C3 ��2���3?�U3��y3HW�3;2/3���2��3�;3�u\3��2�+3S�-3L'3�Q53��3�!3�e�3TqP3��93�)�2Y�p3w,d3��3��_3ڬ3z5k3�3p�3�qU3-�E3�`3�� 4��W3�r37R73�F3��-36�Y3h�]3�.-3��3< �3S�3&��35��2BH�3�Wy3O�&3jg333e3��3��3e��3�733�p3ʂ�2^5�3���2R�!3%��2{-:3o3��f3�43�N3�03�R3M$43�3;��2�<�3�J%3_(�2�Y�3�3�Y%3eA3Ł3���2U�3?Q3;�3�#3M�3�@i3|�{3�,3ћu3w`�3o�d3
�T3!��3,��3�/4��3w*4�8H3��R3ӄ�3�z�3�!�3Z�3Z�3a+W3�3S��3lڬ3�53�Kp3vnn3B'f38�3�|3A��3�|�3ii3��3!�z3383@�32��3��r3@�Q3�fE3��13g/�32�23&Ƃ3��3oXv3�1a3=�3&""3��3�h�3:��3�A*38F�3h�3P�,3 y�3��144��3\�3%�2�x`3X��3~3\3/I�3�/!3,�`3��3�ݔ3�~3��3Ý\3'FF4Z
x3��*3kB�3w�Y3�,�3E<p3
��3qE3\8n3��"4�\�3 <�3�`3V[E3(��3p8/3��3]Z3M�3�#3���3��@3��3�Y3m��3s�3T7�3��d3<~:3d�3�3��D3�_&3?Ь3̎3��3�3�3��/31 4�O�3��3��3��3<2�3(�/3ߝ�3�E�3�{03�*3�H=4�	H3��3�`3�ھ3 V3T�3��p37Q3t,a34�3�ȷ3i˫3�3��3��3p�3�̨3O�Y3�Q�3�>+3�G�3��33�5M3��/3N>4ݼ�3q�3M��3Zt�3��37C�3��3�r;3�!p3��4�3�|V3e��2!��3��q3�\D3���3l�2�Uv3�Ѻ3B��3�2�31��3�OR3�R�3�K-3ةo3]�3Yt3?7m3\�k3��3L3�G�3N�3{1�3*lO3�sD3��3K�s3%T3��_3m�3�_3�>!3�@�3�{V3�8b39\d3�#�3��`3�F�3��3��3�13�M3I�3�i|3A}3k�4��3��3��W3H��3܇�3��K3���3��^3%�3b]3yq�3_�h3�[L3&W�3Q">4 �73�4�3��3^�3xE3��3��3�$63Z�4�	4ʟ�3���3A2�2I�K3�
a3��3�[13�]�2�ʸ3Қt3��4�^T3'��3X2�3;�4�x�3n�37��3��04�|3���3���3�:�3��3�/344�e�3{�3��4̓�3�X�3�(�3�m�3�4D�300�3��e3P��3��3��%4��3"�3-�3��3N��30@�3�:�3�!�3�̤3�4�K�3^��3W�3:��3�f�3��3?�X3+x�3)�3h�a3��44/�3&��3��3�h4d7�3PB�3Kv3�[�3�j3�w�3���3��3h��3��	4Ǐ�3Є<3���3
í3�3�3"��3�!Q3��3�-3k��3�3�3���3��t3��D4y7�3 �3!8�3���3�44�c�3�v�3=
�3�d�3R9`4�{�3tQ�3� �3�d�3�B4��T3FG�3߈�3 �_3H�3��4�Ƅ3��3���3��942:�3��4�3��03Pq4�x�3y�3=+�3�#4��3H94�Y3vv|3��3�r�3 �3��4�Z3u�4���3(�3 �3e$�3P�J3��4�ȩ3}�3��3?4	�3e��3\4\[3�F�3�,4�4�=�3i�R3<��3���3Q�3T��3O�3��4&r33̐�3yy�3���3��3��n4l�3s��3�g�3�H�3�N$3���3k�4�K�3�<�3Ǥ4D�4}=�3ew{3�4��3hަ3�;�3�� 3�g�3�q3-�3��3�*�3�4�3�u4��o3Ri�3qK�3>ʲ3
�3S��32�4ޜg3H�3�gJ4�Z�3�o�3R�|3u)4	}3��3,�4�D3cr~3��P33*4�}q3�O3(�3<��4�@E3���3�4&sC3��3x�p3��3��Y3?M 424o��3���3�nd3U(�3�470�3��3�[�3�K�3��3'��3͟�3�QK32��2��?4�3д3GJ�3r��3��o3�CA3��3���3ZU 4��3َ�3�6�3�O3y�84h�3~��3%��3�Ć3���3%v]3�4Tw�3�u3S�3���3"&3�3��;3�2�33��2ΠT3��34�3��f3R�4��3<��3��3�j�3��3��2Ե�2� 3�a3���23+�3��Z3*c{3�3h��3�/
32�3tAZ3\?�37�>3}<;3X3�{3�3)��3^��3A��3`�3�3��3X�)3��[3/=3��m3k�3_�3*��3��3[�23���3P,�3V3��t3��3��
3��3��_3���2��"3�4�3� `3n"3s/345z3���2�[X3�;s3���3z��25��3�^%3�7�3�}�3@��3`?3��A3"�.3.I3x 3(��3�$30rG3!�3��3Y�3�23�93�o3C�3c�3�K@3���2���3�~3�ۉ3��e3�CN3�,,3�&4Q,3?�r34o!3��.3�T&38F=3C�P3�,3��3tuk3�T�3W�S3��3��i3S��3�Q3[��3eV=3�/�3+�B3���3��Q3��R3ze^3�@4��s3os*3��!3�nJ3]{03�bw3�m3�3�<Y3ke�3��y3ŋ`3�13��3CX;3N`�31J 3�23JU^3͊(3�4U3=�}3U/�2��2�T44 �"3Or{3j=3���2n`3< b3F3<R3Y� 3oV�3�ٌ3;�,3�3e3�3Y3�,3�E3p�3�Q3x3 �_3��3�|	3���3-��3H�3�w38|73�2�3�<3}�3 �3���2k�?3@K�3>ڋ3��Z3]3Y1 3h�3�}%3�mx3��3�#3P!3K�3.�3r*h3�J�3(��3��3	�C3^k�3i.C3��=3�D�3�X�3�mE3F̟3���3	�|3�GD3}hC3�U�3�fo3��	3�L�3!�,3І3Qq�2�p�3�T3�@-3�yI3�` 4�q�3U�3��i3�i�3��3�B>3��o3�'3A�*36
�3�ا3Nxy3K�3F�83.�T3�4O3�ƛ3��3���3C�03��3��C3�ؕ3��3�%�3���2�~03W�2?��3��2���3Rl3(S3r&i3Ri�3��83 M3s�3l�O3S��2���2�3G3��y37ڢ2 ��3fv30�3z�.3�d�3��#3+�-3�h�3�33A?=3��:3��i3\3uA3���3jh�3�y?3�`3�3��3�.(3Ϲp3�h63�w/3�gv38ޚ3t�U3�E!3���2ܬ�3��-3��+3�y�2yh3�/3m53���3G�3� 3Y�3?Z�3%!3��2b�N3c�V3U��2L�k3c�j3�A:3�N*3�xL3O<3T\s3�3\��3�3�=�2�l3u�63_�_3�\L3hE3t[�2�I3��I3��3�Z3���2��R3�,3��%3,1+3gF:3���3��3���3��>3	�@3|�i3���3�L3��H3Rij3��34P�2�	m3�O_3$O35c53/_4G73�Qe3���2�=�3'**3���3�;�3]� 3p�3%@3��3�3a�=3}nY3���35,�3��k38b3T�43%3fK3�r}3�2�3�z�3�P�3���3���2/ �3h6v3��r3��l3�l�2���3�G�2�ބ3�3,�M3l�2o�4�� 3��83�b�2��R3��r3V_3�ސ3�3`3��z3}��3si39�[3�s3r�3�2}	�31(3��y3�-�3MU�3&��2�3v�3@��3��303�/83A�K3�O330KW3#�m3��3��[3I�m3�]�2��13��2�UG3�HG3.�?3���3���2���3�,3�E�3=�3L�3�3;X�3|N3Lԃ3�l@3�x3DA3��I33�3�,3*=3oN�3��A3��s3�x
3��3��3:�3�h3�Ƒ3(��32�3�[3;`3�.3�\�2]��3ްx3q~U3��3O^!3�V	3v�M3y�33���2&Bq3Q3�/�3&�@3��2�(3�"$34�:3�s�3�+�2܎63Y�3s�>3y�73!��3��3fR4�pr3�u�3ZEN3.�|3��s3���3C�3��3���3O�4M�3�"�3V�R3;��3���3�^M3*�3&��3�d�3.�_3�v�3�\�3�L�3��3�b4k��3�ߖ3{+ 3S1�3���3N!�3��3��3���3�l4n��3��k3["3��4\A�3A�B3�>�3�3v36��3bY|3�n4�(�3��3���3��)4�3>�o3���3DI�3$"�3���3�{�3~�v3N�3��'4#34�L�3��3i�3�օ3��O3M��3�q\3��3�΅3y:�3zR�3��3�k�3W�f42�23)�E3��3���3�a3�63���34�83C�3hQ	4�!�3��3lwz3a�3e_�3"k3��3�r�3���3ɒ�3���3)-�3l[�3�x�3oYH4���3��3�K�3�{3�\�3pu4���3��W3��3_��3�>�3���3�zM324�@�3y��3 8�3���3�\�3Z��3���3��3��3�՞374���3/��3=��3Y��3��d3���3>�3�Z<3v�3Rz�3��30G�3F�'3I<�3I �3�6�3��E3=�L3A�3�xv3Tǉ3��D3�+�3��k3([>4v�u3Q�3,˸3*��38@4t4�ɱ3)ܼ3z��3�VR4�z4�U4�(Q3ר�3�D�3���3G^46�3� �3�*�3�t�3��v3Py�3כ[3�]4V�3���3��z3�M3�130�3���3O>=35��3���3�׭38g�3��C3h�3*�S3CdS3	r�3�F3��3���3��4�\�3���3�ff3V�.4A�4k��3��3�o}3�b�3�{�3���3<Kk3'D�3A4w�3%4�+3h�l3e�Q4v�3�q�3t��3&�3�ˢ3	�3*�3_�<3�C3�I4�~�3���3F.�3�lK3�3�3g��3�E�3%��2��3�4��44�[�3R�33 ��3��3�
�3��3z�M3Խ3�Ń3E3 4�{�3�6�3���2Z��3��83�w/3�� 3LT83'#3���3U'�38tB3�93��3�.V3�H3�;,3i��3P�,3��3Ԉ33"w�3��3���2��r3d23x	#3�e3B�3�W3*3�x3S�3�d3QJ�3�s[3��2I��3]2�3�U83�	�3�#�2K�3�123��3�3��[3-�A3��2���3hO3�3�U�2���3� 43�fq3.�3hA�3u�2�`3:Tm3�1a3Ave3l��3�R[3S83:��2%��3�Sb3���2S�33k�2��3{
3�`3��3��23�`c3l�3O;3��l3`�x3��3E�T3ޢ-3�3�e'3�W 3[��3�
�3&y 3w�3�g�3U�3
�2��L3�M63<n3��3
�3�!$3_��2G2P3�̕3�m�3נ235)33M�Q3�A�3w�n3N4�3<�/3�_3�B 4��K3<�3���2�p�3��3^�53�-�3�3���3~�n3��k3+3U3.3�"3)|4C�2�@�3_�53Z�-3��@33R�~3G`3�!"3�q�3�/�3��3�~.3㧹3ND3�E3_lM3�g�2b��3=3Z3���3��S3�'�3Q3
,�3��3v�3/��3�"3��#3n&^3\�3� �2���3���3��3��3=�=3�c3#3�);3[Ta3�d
3=|3�|�2d��3�6r3h�3
8�3��3��p3�DR34#�3��3c�K3�<)3�_^3Z�3Xp}3�B�3�	r3�303�i3��3���2�)�3�A3\_3�n%3σ�373k�3R3�z�3$}E3�=�3��N3�3�r�3b�E3oZ�3JcJ3�43z<�3�_3Q�T3���2V�{3�1B3�i!3��3Ͳ3 ��3��2W�3��D3Ď�2�t�2��Y4gc@3283Ӗ3{]3l �3�?3{iv3�43��3���3J��3Q�3�53g��3�j3�H,3=g�3):$3��3�)03n`�3��3���3�aS3��3�̃3��3�g�3	@�3�P%3�q�3+$�3���39�3�P�3&��3^�3743.T�3��3u�s3ƃ�3u6u3��|3_e3nT4���3	��3j1�3��3a��3Vb�3a��3?�3p��3a��3E2�3�H3J��3:43��3Ɛ3�?3�ލ3Bg�3���3�[�3��3���3n.H3�c�3B� 4�`R3a�$3��4�Q3v��3`*�3�ڬ3\HE3��3�ȑ3�sk3�c�3��64���3���3@#
3ݭ�3�4�NE3�܎3{�3�P�3�
O3���3I��3�}�3 �>3�4Pҿ3�\�3±3��3��	3��3d��3��3�n�3��3��3�i�3M�3)��3�s�3
�w3��3�]3��3{�34�4�p�3�|3Wqo3G�P4`�Q3Ϡ3��}3uu�3Ș=3O6�3c�3�|3��]3��4�24���3�D3c��3
.�39tc3Q�s3��3���3P�d3�3�:|3���3�D�3S^4=d*3L�o3Q�X3�N�3��R3��3`�`38M3I23)��3�3��3ɍ�365�3R��3��3�x�3�8]3�F�3%�3�B�3w|73<Z3��3l[4-�3 k�3��i3���3?N�3=�3���3��3�g�3���3�N4���36)3�3a�3�Ae3!Z�3Xǩ31q�3�2�3lf�3�8�3u��3��3,�14�3�3q��3�k�3<�3lA3��3��3ڀP3",�3:,4i{�3�P�3(CX3獀3v�3�q3CR�3��3W��3�ɔ3^�3s��37�;3�aM3�wE4��334��3W�3�j�3���3\m�3
_�3wA.3!f�3H�'4Ơ�3T��3'3���3n��3&��3���3�@d3��3�Ԍ3V9�38I�3X�_3�^b3�b4�)-3��3鑴3:'�3o�K3�E3{�(4��y3/�3�*�3,�#4�8�3*B3p�3�	�3	 �3�3��3si�3v3/[�3���3Ah�3��L3���3�9�3?�3�'3Nļ3}�W3��3r��3kJ~3�P$3�2�3��m3��3;�\3�ɴ3�Q:3w�O3T?3��3�6�3`�V36�3Af3Ѕ�3�-p3��3�i3Im_3�<�3�6v3x�]3B��3���3yl.3v��3cR/4�J�3�-�3s�L3���3cЗ3Dr�3Ⱥ�3��3O��3M,n3ە3ޠ3�63��3���3>�%3�K3�S3,��3.�$3��^3G�D3��-3��\3Z4q��3�X�3��33��3}�73):3ߜ31�3�8�3\�G3��4���3S��3Y�O3a"4��X3>3��G3�3��,3��13A^�3<(93���3o�J3�A�3`��3o��2<��3 �3�9P3��r3��S3�R�3��S3c��3�p3��73��3Oa�3)��33ྔ3�A3�t�3�"�3���3z�53W_3qޖ3�ڑ3�3vL!3�ڥ3!6�3�K3}Q�3�J3I�3��p3��\3�x$3&<Q3�I�3���3�KY3�z�3&y�3(v�3��K3�f23��_3G3H�:3-�3���3�u3r&3D>^3Sv3nN3ҕ�3��33��3/L3���30S3�g=3M?3���3JS3��_3���32L3��%3�/3
�3�<3)߲3|�:4dP3#�3Y�+3x�3��g3�3'f3u�3�K3�'3D�3���3��U3��3���3��f3��83�D3�%�3�*3�O3�J�3���2~��3ȃ:4��3Y�3zV3(�X3{��3d�:3'��3a3�6�3�43��+4��=3�H3,@32�i4o��2��3@O3�3�II3p�t3�37j%3,��3�3�3u�W3U�m3}�c3�Մ3��3��A3U:�3�+3mL�3�yc3��3:y3�.73�O3y�+4��33�7�3�a�3p��3�	O3��G3F�l3}n!3�3�c�3���3̀4�D3���3�Ԥ3�633~�p3+��2���3G�3�M�3�B3��3�_�3�41HF3e�C3h$e3־�3=�-3lܔ3r�3>PS3�&e3dtx3�w3;��3�M3hL�39L<33�'3f�q3�<�3o]�3J��2lb�3�#�3�R�3�|3�P�3B�]3��3 Bi3�Y�3�x�3��3̡3��3�}Z3��3CZ�3ߙ3�3�fG34�b3��3*�43c�28Q3�ڥ3.�U3^�&3��3��3�t�3��63pЙ3v�32�o3_�R3J�43S�w3��Q3�W33���3�u�3%�^3D�$3E�3}w�3�93�{m3x�3��3�C3�H�3ώb3D�?3��t3p��3e�2�U23�3HP3Ԟ^3�'c3۹�3�13��z3eQ3�c3�3)O�2.�3_z�3a6�3��N3��R3�[3�d3��3��a3G�s3��3IJ�3��26@3��Y3^3�ǁ3�l3�vv3ϒ3 ��3�G�3�ۆ3<��3*�2Uo�3���3���3=�3�3 ��3;�3��p35<3p31DT3���3��35Da3h�3ne33��J3���3i�3ծ�2c��3�ƥ3TQX3�3383I0�3:��33?P3jB�2U{3i�O3��_3>Y{3⡰3$׃3�U�3��3gs3�9�3�?3p3#�3���3H`�3�&3#�3B"42_�3�*?3�ʀ3ɔ3Xa�3A_3��y3��53��93_}3��o3�T3��E3��T3��3G�3�gG3���36Mj3oQ�3��w3Ɦ3�E3~i�3[B�3dd�3R�A3=3>3�ڽ3��s3*Gu34�j3h��2��3%�03�U�3��|3	N3��@3��4�s3�!3\w�3mZ�3r�S3B��3Cf3N7�2Kц3���3UCv3C�}3��2�Np3"]�3x�3/i�3�+$3ۭY3�M3�û3�s3�-T3�~(3��4F�+3/�3��%3��-3��3�`'3"�V3��
3�z3�ƨ3>��3�ͤ3�q93҇3A@�3*w030�D3=� 3U`Z3�63!%d3:&3��W3u:3b�3��2�{j3.��2U�2~�2�@3��33��M3�3�i3��63	�d3P��2�W3��3.i�2�3�*�3�&3E��2��k38�g3L�u3Z�2�i�3��3� 3�3�B3NG�3-�23!rS3��3�(#3w;�3$��3��3��3Ri3n3Wl3��L3�D3�Z3G��2T�G3�k;3�q3�+�2���3?�[3�q�3P�+3�:3CY�3�Ɠ3m�3C��3�23hu�3�Sz3e3Y�2�Jg3HfF3�"3o3���2�%3>�3�C�3�_S3���2:��2���3�03��3��3#�}3M+3�� 3tc"3E3dl�2-3�3��,3(�M3�n2BB3��-3)��2�G3DUl3���3���2̜k3�]�2�^U3��3ti�3Q(�3N(E3�v43O��3�3�m�3.�3?'3��3^�s3�3T+323g�B3C3�37��2��3�3�t237|@3���3l�!3��3le�2�3��D3��"32m�3BP3镙3��Y3�b83S�3��3@1^3�˖3��3�2�jM3�5p3�
3�	)3_��2�n3��o3�3%�35�83I�2�`�3���2@��3@D;3��c3�;3Nl3P�@3���2�	p3�<�3�)h3s�3`�2���28�s3J�2�j 3���2��R3Ў�2�V3�483t�3Xu33�
 4\��2�6�3p�E3T*3��3���2��$3���2�V%3��3��_3�7*3=s�2⒂3�� 3�m�2B43YÈ2�:3YI3�qG3s�2�� 3�.3��3��38��2+�v3CyV3)S�2��s3��|3��.3ZvA39��3ʕq3O�3���2�t3��P3�W53�k3o�f2��r3��2���3��2�~03�B�29�3�F$3p��2�\L3��3��2Bp�2(Qd3�3��3���3��3��%3[-�2
X3�>3�#3�р3K�2��*3j)�2�t;3 �J3=�402'3��/4��3��3�3y��3$~[3bA�3�C4���3�3��4�D�3�4�33��3z�3��j3��3F�G3��4Ƙ3w��3L��3���3�4�3^�4�jO3��3�Ֆ3  4��3;M4�Y�3�]3��3�'4�C+4Bn�3"3�V 4᭰3�3���3�o�3�!�3'3���3��3���3�h4k��3b�3_��3��3I��3�n�3��3Y��3@P3�Y�3Ó4�'�3�Ҕ3)NM3t;�3Α�3�Q)3_�3>��3�o�3��I3�V24ǳ�3aH�3�c�3)�4�q3WҚ3���38X�3�jk3M��3Jt�3�p3�k�3�4�\ 4$�3	]G3�n�3��3OĚ3���3纂3���3��i3v�3�J33� +3}A�3�1"4.�4䎼3a�3�3�3���3Q�3���3�!�3h�3��3���3�Cw3P��3�x�3U-�3���3�Q�3%4"�3��4�7�3��3*��3�D*4<��3�Ƭ3��63��3�x3L��3Il�3!�&3��3B4���3�sU3�n3���3�g�3�U�3��3�k�3J��3�a�3-4H��3z	�3H�*3fY�3�*�3(�3ӝ40ݟ3��3i��3���3��3���3��
4�
4���3�V�3ܰ4|R�3	�3jP�3�.!3n_�3��3��3��3�]3�n�3�4$�3sG�3KpW3�b�3Y�3C7�3!ѻ3Ო3ܛ�3l~h4���3���3qV43�:�3�4�3�J�3\a�3���3��K3z�E4`��3�F�39~�3n2�4p�3=݉3sp�3�L�3ؕf3GW23~b�3�y�3�>�3 ��3F��3I�d3��&3��3��3[_�3w��38	3���3�r3���3�fk3�I�3vZ3��i4�M�354�Ƀ38T�3��34��3d˹3��(3�/�3f4a��3P�4B�33�u4L��3�R�3��3]3A	�3Ie34p4y+J3�m�3�7�2;G03���2%39�C3g3��2�
3te3:G�2�Y3�j3���2|�P3���2EN3���2�p�2���2�N63��3{x�2�+�3�3��A3�h3���3L��2�f�2�l3��&3��'3��t3�%�3	��2e�2�30�23r3b��2,5I3�̰2���2q3S^�2z�3
�36�L3��'3��J3(�2�f3l�3C�24�2[[3�%�2�3P�J3�l�2�P3�qc3N�V3���2�q2 S�3��3�o�2�623W#�2��?3h(3i�>3�2b�)3`&3m$�3:39��2�:�2<�2A]3�B3>��3 �2��I3�M�3��J3�h3>�[2�
3��3���2)�)3���2�S'3�ۘ2�953M��2���2C߉2���3oI�2��2��3�6&3�4�2��?3m��2��2[�!3DH3�_�2�3_ѯ2��3��p3�D�2�}3�0�2�3x��2j5!3�\�2��2��3S3~��2cXV3��3T�`3�< 3H�	3���2�6�2�3�"�3�03�!-3j.�2��,3�H3��3�O43��2_�3'�2�(3d�3��R3)�2҃�3���2��,3�>3mc3�Y3D?'3ժ(3(,�2'923o6�3^b�3Z�2~1 3 D3B�3�?3�i=3S��2��3�3�B�3q�3yq�2���2��3��31�`3�q�2ؓ�2g�Q3s�3��43��3�]H3@�3��z3�3��2ł63(h3��.3--#3F;�26�&36��2n_3��s3�3��2�B�3��2��X3�I3�x�2A.3b!3��(3u��2�X3��3mGI3s3V��2�3k�\3}K�2T&03���2�R3���2Pm<3�~�2�3A�2A6S3���2a�3�,�2Ү�2BM�2g93�zr3��v2F�E3Iߛ36}T3��3���2��K3�3�Ѵ2�u	3��2��33�`3��R3�#�3���2z�H3��2B8|3q�s3'k3|3�2��]3��&3D�%3�	�3�D3���3�3�>3�M>3�s�25�2y-3ZI�3�x�2_��3Uw3��t39��2��3�3�@43�^s3�>3-�2��2Q73�H3��#3nX3o'C3엟3�QS2�w_3��2���2�l�2Nt$3 �3���2��]37Cm3�\3�Z3��3�(3��3��3?g�35�73�D/3�53���2��3W�3Y�a3��3E�2=?e3��:3V�2�523�}3�%3Z�$3x�393�W�2)�]3׾�3�3��2�k3�$3��3�uF3��P3��3g�)3$P13�܄3'�3I��2YD3�)53�e�26�3��3A3[��2�'{3�,�2�W�2��'3C<�3�>3:53���2 �)3� 3J�<3�L3�.43��%39�3��A3B#T3��3�H3O3dC�2q�3�:3+33e�3֊t3�3�^3��G3�ð3�W�2�#%3_u�2^3� �23�>3�Ti3W��2EH3� 4&\�3�x�27�?3ͅe3?_30A�2��3���2��[3[f�2x��3��,3��2.�;3r�4*�83̋
3��h3�?�2w�2��3�oP3��3�(3$`@3�P�309$3r<�2�3BK3��/3,�3j/�2��3��2ٷD3Z`3[3|]�2��36��2���2�(�2�*�2cg3��23�� 32�)3��?3֢3I�C3D��2��2��o3�}3�63wS�3�3�K3l3޳�3�>R3��3]��2#+�3�^3C�3��`3�[�2���2�H3O�X3��2�Z3l��3�Il3�.s3N<�2Ԍ3#E�3�m3���2
��2��g3k�2��3�3.��2I�2 ��3��S3.�g3�� 3� �2Y�3,�3@3W��23��Q3/�o3�@3���2�n3\&�2�=�2�u3U�32�"23d�2$e3�XT3���3��]3�x�3�(v3���3#�3�'�3Bej3_��3��}3^53�0�3Q��3 ��3���3)�3�^�3,T�3�
3��3�Q�3�0�3�N33:��3�6�3cƺ3LIt3�P4�ɭ3���3�ʕ3���3��3ѷ3��3$1�3��3�V�3��3���3�Q�3�9�3EF�3D��3�c3�	S3�3�JY3���33��k3u0�3��(4圕3�ؕ3��3]��3	�S3k�388�3N�3{j3�A4t�3=�3��?39H�33��3t�|3�Ct3��?3B]�3m:�3j<;48`3���3&�#30�o4[�+3|3|O�3J�3D�3�g3��3Åe3:a�3v��3�+�3C�B3Y�3Q?�3M5�3��i3�:�3`�3�\�3��3�|�37VS3���3��.3 M4�}v3�8�3T��3 }73�_�3��r3t�3LO3ܙ�3�X4%��3WU3�3Q��3t?�3mp3�3�͠3l�3`r�3��3�@�3m�x3�~3$M�3@��3|Y�3���3yݢ3�N,3��3(��3
�P3� q3ɯ�3���3��3�ш3ˉ�3T��3g�3i1F3Y�V3g�_3<�C3���3���3J�3�r3#�4���32��3\�T3��3nq3K�L3m��3�(3��k3�f4ʛ�3xw�3s �3���3W��3��3�z3A�Q3�E�3��z3^��32`w3-ӯ3��3�/4��<3s_�3��33�n33�,�3@�3��<3���34�3�3_y3ȥP3䓟3o�3���3�1�3��73.��3�sn3��4uaA3*�f3�E3'4N�Q3�?s3甇3��3>��3͓3���3D�S3��3��4B�4�v�3�`A3��3�)�3�?�3uȠ3:�83C��3/�U3��3EB�3�Z3]� 3d9�3��.3��3���3r�a3��3�b3�Q�3BwP3Tó3��3m�4D.z3ir03��3v��3��B3�H�3�4q3��3���3z��3U�3O�3s�43Ij�3�3v��31�3�"4=h\3d�3 ��3�~�3,Z3<��3ʣ�3�O�34�3�T�3e��3�9v3	v�3�_3ι�3���3�ͫ3���3�c�3_;�3�<�3%�o3�$�3=�3� �3���3�3>��3��{3�%�3��
4gv�3]46�E3	��3ɫ3��$474�3�73�.O4�3E˻3���3q�3��3�p"4���3� �3o�*3�q�3Q7�3�
�3�5�3絎3�9�3k�	4х�3q�3�e�3a׺3nm�3��X3ޠ�30�o3v�34���32�3lش3=��3�?>3K�343�8�3+ɿ3���3��H3U��3�e�3��q3V�3y�4=�3�q�3݌13N��32�3z	�2�H�34Y%3Y��3��z3ִ�3@F3�i3���3c��3/�e3�*�3@�u3��'37��3��3�ݿ3��3i�x30��3>��3RY3���3�	�3\z3�~�3!Ӥ3O�3��3�&M3On4���3�0�3�#�3�n@41��3= �3|1M3?�X3y*�3��z3�3xW)3���3�7-4�G4�A�30$D377�3`Ѐ3h̆38�~3�KK3d�3�m?3]I�3ֆX3`�3 AE3�g4YCc3���31��3�y�3���3��\3Aږ3]�s3��304���3�9�38C3!�3LC3/�3K�h3$N3���3���3�D
4�j3�ӊ3~(3�g�3�y�3-��3��S3�ć3Z��3r0�3���3�W:3�j�3V}�3~+4.�3�63�y�3�Qv3��3���3�43��3�83���3�r38>3�3��L4Z��3᭜3鐥3I�!3x�3n��3�4�3Sw3��3J*4��3���3��K3l73�,�3��3�a�3��3)��3�VZ3q"�3��3=232l:3�� 4�C73 n<3@n3��H3�
v3��534��3��3o�F3^��3��4�+�3��43�*�3�3�3H7�3_i4�ML3�)l3��2���3ik�3h8�3�73a��3��O3^3u�3��3���2.8�3�Ѣ3۰W3o[63���3g>�3���3NpS3�y�3ߺ�3�d�2XT3Tq+3�n3>13=��3x~g3�y338��3��4c `3[Ƭ3N��3>�3A�*3���3La�3ҰD3�$�3g��3.�4ټ�3�/3d��3�,�3NY�3V��3���3 �A3��U3�ͼ3�o�3:��3���3"�3�ʼ3�k�3�\31�4iR�3UB3g �3*,�2}�l3��4�[3i3�J43٫�3�S�3�=u3o��3ƃ3gШ3��31��3�*�3��3BM3�9�3�F3�3�8J3���3F�3ּ3A��3ԴO3ap3���3b1�3I83�N�2�m�3h��3-�13T�3�k3��3[$�3��3>�Y3r	�3��X3��3B�3VK3E�+3|��3T��3ZQ3�G�3@nz3�h�34�	4�^�3�dd3���3J��3⽂3�:�3ic�3~�3t�3P�3uR�3־%3��3��_3
�!4C�53?��3�v�3Մ�3x".3r�3$�_3<�R3&��3�74gX�3FW�3^`B3�?3R�v3�983y�3$g3b��3*�m3D��3e�h3��n3��;3��L4���3���3��H3��Y3/\3��3���3� 3ź�3��3�k3*�}3̪3��g3/ �3<�%3��3�=_3��3�]3���3#�o3�TX3�hZ3�U4v� 3 $3�N3n"�3�03���3��3)�3�W�3��3Z5�3�b3C	3M!�3�օ3E�3���3C�"3V�3&Z3*j�3�v3_��3�e�3��3R3]v3��3�^e3���3��3+��3_�3֖M3���3(^�3�ѕ3��3�3fv�3Rќ3Eɟ3��\3xL�3�E3qئ3/�3�{(3ǣ(3x��3��73hX3&�d3�&j3'i�3%�38	�3!33({3P��3��4&M3p�2��3cg36g3�ge3��3�31"63:�3�	�3�z�3ҋ3Hj4��X3cS{3*5�3< 4�*L3��3p��3��3�R�3��54|��3$]4�&�3��4�[�3��"3V��3��3bK4x/�3�`4��3��3��3�f�3��3m�l3���3�2�3��3J�3���3k\3[�3���3�L4�l�3{�E3ӕ4?<�3u��3�S�3F`�3��3�M3���3��3�9K3�Y�3�@�3_�3���3��3�3��#3J�3S�3C�e3��3�Z$4��4�q�3�V3Ņ�3��3l�3���3�V3�T�3C�4Dd4YS`3��3gd3a,�3���3>��3��3|`�3���3vQ3��3���3	�3��24�S�3:�4�MU3z��3vڟ3�D�3�3��'3V��3�3~c4/4z3R�43��23�<n4�B�30�Z36t�3\f�3��f3��32�3|3�6�3�!4�^�3��3Z�W3G4``�3�.G3u�3K4�3W�3��3�4��3��3��3�4��3:j�3Ŋ�3�3�3-�E3#μ3*�3�zy3��3v{�3��3wN�3�dK3��3�w�3a��3�L�30at3ɚ�3�b�3F]4��|3W�l3{m�3�n4x�X3�j�3��B3�0~3kA�3���3��3,Ro3�NW3��	4�y�3�q�3�d�3��3�i,3���3���3�^m3t��3��3���3��3~v�3^��3��'4	�t3���31�3�e�3���3,��3�s�3%�=3��3�43�4B�3?d3�Ԍ3���3�(�3n�4~3�ۉ3SF�2Ji	4o�3�A�3�43̿?4���3^S�3��3��_3��3	/�3�v�3��t3]��3��-4#��3�S3c�3jܽ30��3}�3���3e`�3�N�3�:3sm 4��z3�q_3J�~3��4��\3b��38�3�N�3yG3J�~3��3U3:ȉ3I64�+C4�\�3P�03Z��3��3��.3��3�:3S<�3%}M3��4˪�3[YK3ؗ3}}O3��3�(3˦2� 3|��2
[3j�,3�3���2���3�3��3$�3�O-3�-3�*�2�{2��H3�=3���2�:3��)3��3�7�2�e�3][�2���2��3I�33A�2{z3�}�2̩�2�/3��3��3�|;3�[�2�@{3�tq2Jس2�%3\֚2��2�*%3���3ҥ�2���2
�2�43D��2-��2�q+3��3��2`l�2�b3HY�2|3!3O��3��93VY�2HK2^�C3���2�|�2l;43l��2�=3���2�IS3��33[3p��2��3���2�d3�h�2b��2��2W��2�D3��2�2Q3��3�y13u�3v1�2t�#3�o432k�2�='3��2��43�թ2�LQ3�e3L�63��3O!�3�q�2�23l��2��2ރ�2��2v?�2jh�2q3dV3&�i30�2��2P_3��2��3��.3+ߑ2�.3N��2�3$��2{S�2e��2;��3Ov�2.��2�63p��20��2H�2M�3FX�2'$ 3�e3�*L3��3�6�2"�x3��2�۽2��93w��2��
3!� 3��'3B�2�&3-�3��N3k�3GT�2�O�2 ��2ǟ	3�;3�3��2�53
��3�=�3k3�͊2�؎3�Q`3���2��'3��2��%3B3}A3���2`>�2OL�2�CG3�?�2n�3�� 3}S�2�;�21rJ3)Pk3?��2�3TDP3�M73�(�2 �2��O3�C3/̆2LM 3�x�2��24`�2	�f3;'�2�I�27x�2��3[3o�X3��3c�23�3��,3��27L3�
3�73-XS3)��2�� 3� 3a�2ބ�2qW�2A.3m\�2�e3�=�25�&3�j�2���3R;�2�ya31��2�m�2	�2m�83��3��P2�6S3S3�W3V�2a��2g<3Z 3���2V"3���2A~3$]3�p3|w�2a�3�َ3���3��3��Y3�b3Y3833ʉ�3Z4�3�r@3(ō3��&42��3[�3a�(3Iq�3,g�3(PW3�oG3��3�`�3A��2�V4��3�3�g3X�4�{3/A�3��3���3�z3�X�3�H�3h�3���3�ѓ3��3u��3 3ӗ�3Qk�3�3g�v3��g3��43IH^3��3�^3��3Q_�3H-�3&��3	�_3�S�3��3#|3�23���3xh3 V]3��3GG�3w�i30�$3��}3֨�3% 3�)p3�533���3�ǡ3\%�3U�i3�YW3"݊3���3�ڀ3˿23�e�32(_3A�-3�B�3\��3��2Ν�3C�/4�3AX83�3zc�3%=3 �3�=R3%�23���3}?3|D�3�B3���3 k3C�F4�W3̐�3N�g3�[[3]L=3��3`ϔ3h=o3pԳ3=r4�Ѵ3��L3��T3x�3���3��;3&�3^� 3�Mb3�0#3ǣ
4�r�3�3��]3��3���33�3&ľ3�ծ3�+:3�%3��3W�/3�$M3�}�3��3Εe3FPb3��3��3��n3ՙ�3E�3���3z�3ю�3x��3G<3�<3���3��f3��3(�%3mJ�3U�3�ɢ3w]�3w 3�~l3�I�3��3��3΂(3Z�j3�!�3̆3��3�"83�_�3�H13��4-�f3�ӷ32��3�K�3J"W3)��3�3�J_3v(?3��3ə3=��2~ �3�4\�3?'�3|�g3:�3���3�3>3β�3��3�ؐ3��f3,2�3SUi3�`j3Љ�3$!�3EmB3/d3��i3��3y�d3�n30H�3��2W��3-b3Ze�3	V�3�3�'�3M�]3�3�ˮ3x-�2٩36(Q3�F�37';3��43�KN3��3��n3*�3"�3��3]3lIV3�u3�&23O��3� �3M��3�v�3�E3v<�3-��3�#3�ô3��30�X38T03�6g35P�3��(4Y	�3��64/q�3��3&��3���3r��3���31�4�M4N4Y�84���3��g4�֪314Y�3��3T}3�}�3�
�30�e3�=)4�L�3��3�)�3��4#�4�w�3�.�3�*s3���3)4c��3/�3?L�3d2�3?4��3�(�3r��3t-4e�4���3*�3g��3�3��R4W�3Y��3�H�3j�4��y3i�3���3�5�3�`�3��3��3@�3���3�pX4cw04��3BW3���3H��3Y��3T��3�3a��3�լ3�W@4�E�3�y�3\��3�;J4�M3�@�3/�3~ 4M��3�P�3��3�J�3��3�<_4���3 `�3O��3�L�3��4v@�3���3��39��3��3X�3RS�3�3�3�b�3_�24rR4���3vi4 5�3���3�e�3}��3俀36��37gZ4�}&4�|�3�X�3��4
4�4Л4@�3�3��3���3�s�3��}3�(4;z4���3��31l�3K8�3��3
4B+4���3Yӳ3&4��3J��3'S`38541%�3#1�3�A�3�c�3^8�3[�3�*�3�
4��3�є3E�x4Y8�3!8�3خ3K��3�
64@�3(��3�7�3I�4���3�9�3n1�3�v;3���3�+4d}�39��3��!3X�3���3L�4�Ú3��3z��3��y4��3�"�3XG�3R�3��3��3 :4J��3��3��	4M��3�v�3s3V�4� �3qm�3�4�s$3+�37R�3�94�T�3�p4��3R�"4�e�3 ��3�*4;ǅ3'ۡ3�c�3���3zX23� 4n4�t�3~34�=H3��4�c4�d{3;*�3�S�3��4Ҁ3�Ѩ3&�4���3�K�3F�Y4���3�J�3���3���3�Zq3Rj�3��3��3о4+k=4�34�k�3�9�3o��3�j4�f{3b� 4��3԰�3���3@�|4K8�3�O�34�f3���3�6|3��3,1�3��B3.;n3Y��3�53epi3�,3���3恡3 2T3g�N3���3 B^3�G3_O�3qw�3�'r3�3�&�3	�31-�3��3��3i|L3��3�]U3�_�3�>�3�N>3w~3U��3U|�3ԡ�3va'4=�z3?-3��O4��3ϧz3�[3Rx3��3��3�F�3��3 �3[[�3��
4�'G3Z'�3��Q3���3�Y3%2�3>��3HM�2N�~3�cu3��3�L3�3�3�3zX�387;3Α�3v3�23�"3�Q�3
��3G~�3x߬3��3N�l39B�3L]�3��3���3�;�3/�4/��3Ȳv34}�3�Hw3H��3�b�3�ȯ3~y�3y&x3��3~�3���3'?e3.��3ؠY3[�,3hn3��3'd�3�093���3�"~3��3���3�``3�F3ײ~3�$4�z�3w~3��*3�Ǖ37	�3 ��2&��3�GR3t��3Z[3��3ߖ�3WQ3��3�?k4���3B��3���3�U34��H3���3�1�3���3��m3�S�3|�34��3�}\3m��3cm�3)��3ix�3L2_3�*4}W13���3@I�3�)D3�G�2�Gg4��2��^3K�3���3|D3vw<3�A�3�\�3_��3���3���3�0V3y�3�	�3o�3�G3\u�3��2��a3"*.3O,�3�Ɍ3<r�3�R3�B4e�$3�SH3�733^�3f�'3���3`� 4x��2��3�$�3��3i�A3�.�3`y�3(^03��b3#�R4 W�2B:�3	v�3Mf�3���3��g3��Q3C�4_�93Fl3��40��3oF�3|c�3��3s{�3xJ�30j�3β�3���3{%q3�3{3�*�3��3u�}3��d3r04óq3%�e3���3*�$3=|U3�)L4��3J�q3aY3��M3h�y3|�m3�%}3��R3|s�3K;�3���3�~3�P3���3��{3�(g3���3l/*3`3��3Y��3-(�3x��3GnZ3f6�3�|�3�Q�3�@N3t3�u.3��35b�3�B630�53h��3�ݓ3�`�3�B3��3�}3}-M3y�3 K]3xb3:q63꿽3��[3z3mZ\3L��3: +3�u53�j3-��3��2��3�C{3��3t�i3��49CY3Χr3Z�2�a�3�D�3��t3_:�30V3FF�3��3c�3՗�3m�3��2��3�߁3$P3H��3�2�3@//3 �C3�@3��?3�]h3s��3Q�3(�3}��2]vW3�~�3>!34�m3�_3�Ş3дG31�l3��~3�>p3��63��	4r�=3�3��P3�_3.;36�3T�3�23�B3�a�3Tpb3g��3�O�2���3���3N�R3e��3w%3��s37�+3��3��3��F34�k3���3ѐ�3�]_3�v3fFO3���30�3�#{3I�\3��3ʵ�3�'�3o3 4'�P3���3+(�3%I�3��3%�53fǼ3���3M��3���3]��3�8�3s4':�3�Ȟ3�P�3Uz3�'3�q�3]�3钗2�*93NV�3m�3^�3�d3��3�Ɣ3��3"e�3�ג32xc3Y<)3���3�.3ȅ 3��I3��4O�`3,�3�I�3�ȁ3:�3�3���3+�N3/6�3�C�3�v�3�6�3qAi3h�i3W�g3��3��3Ci-3��3��3M.�3ٵ3
�!3�{�3���3�B3��3�Ê3u9�3\`�3љ[3��3�yE3U��3���3fɚ3ҵ63΁+3管3��3�q�3t�3�mA3wg+3.�N3���3 �c3��`3	�e3�74��#3}��3�7�3��%3�ݐ3j�_3�3L2�3M�3c��3�/�3_n�3�B/3<�3���3/	�3�K3�iV3=�3P��3<��3m��3	�93Ъl3�=�3�Y3��f3EJ�3�E!3 }�3n�3��3P�3��3,�3Ѷ�3���3U:3�1G3��>3�#3h�y3�}�2���3� 3(��3���3\�v3��3���3�� 3}�"3��!35� 3�t)3��Q3��3�Y3�$3ۨ�3��3�e#3HRD3�/�3-�r3L^�2��d3��@3u�{3p
3�9�3~`<3�h�35kj3��3�$3�3Ê�3�u3�JV3 '3�C3p3�Å3�'�3�3p�3��3D�3$5O3:�.3�'3Z��2��G3|F3�D�3��?3v"�3*�3���3�H3=
b3p63�lB3�l3O�Q3,�l3�2��3�؊3��3RM^3U��2��A3UN3�.3ь3��=3��3 ��2�K�3*3}�X3��3�=4l!M3�V3�L73T�T3���2jGq3Z3�93k�L3�>�3Պp3 �.3/�2T̚3f�p3�4�21p�3EP'3�13�1�2`!�3�~3|�2�.3Q<�3�DM3�]<3�03?�?3�{a3't$3i�^3��2*nq3���3�I�32i3�`�2�3�'�3�P�2��p3���2E��3�u3�܆3A��2f&A3�a73�o�3�3��3��{33j~3Ԫ3�d�3Tc�3r3�&g3=݈3�Jz3Wq�3o�3�q3�>>3J�2M|3y��2�Ң3�X3E�13<�^3H��2��u3P��3��3�3X�U3��3 ��3�\83C��2?��2_�<3o�3�Y3��B3F��2�i�3�(3�E3��83S��2��-3�3-�Y3>�3C �3�>93[��3J[�2��K3��=3�?'34o�2�=p3���3/�23��:3��4t0�3��k3��3u�N3�"3 �B3��@3ǊX3�8�3���2��3�q+3�3C�\3���3`P3��^3	gN3rr3
213!3�~38~3M�S3��z3垪3v1]3���2��t3A!�3��Z3 lB3C�3�c3�2W�3�3��3��)3�~�3�!33d��3���2��33	}93�8357�2�Y�3��f3��3G#�3�\3�w<3�b-3�3Re/3���2hƿ3g�3�zC3��a3/4)�p3���3�̃3ǐZ3�63-[�3	3�Ǖ3��3oe�3�$3�	4i��3��3P�f3p�3��z3'3ޞ`3��i33d63>�23��3�Sl3]�p30�344 �3�0�3�3���3ѫ�3B�h3�a3�͎3��3ܪ�3���3G�3ū�2�a�3/m3X�63ߦ,3-�;3��3k�3x"�3C�k3ԥ�3yO3:�I4�eg3E�3x�23�)B3(L43 �3b��3k&3��73��3-Α3�r�3��.3^��3�"�3�2�2�b3�A3}��3��R3w�3�΀3�{3�t�3[��3���3��3��3���3��P3��3��Z3���2�Y3۞�3�7�3�{�3���2�}Q3��"3Q�B3oS�3\73��x3U�:3v|3^�L3�[o3���3"�4��@3�u3�E[3�Q�35l�31�3y�3�:;3(�o3x3�3��34�$3O�F3���3~8�3n�q3�0�3��[38�3�>�2�G�3�3�3�;3>B�3�
�3Y	�3ݍ3�3	�3�(E3�ʇ3c��3�M3<2�3F|�3L	�3'+^30QV3�3z�3%��3:�3�V}3��g3F�x3t6v3�+�3N473}7X3�T*4V�3��a3�i3M&53L3���3���3:N3.|}3f��3�c�3�`3>�2�Z`3��3ko�3gr3��3��3�U�3��3~�3��d3~�=3��%4m'�2��3��2j>3fI3�Tp3�T�3U0�3Ι3��4y�36�)3C-3@y�3�=3}��3���3�B3R��3�B3}z%4��T3���2s�(3�x4���3�731��3�e�3�tt3��=3L-�3��\3���3i}�33^4h(�3Q#.3�'�3ߑ�3ʫ�3�c�3�53AǬ3��R3���3�W3LG�3�}F3�y4z�3��3n�3��|3�D3}~3VZ3}��2�ߩ3�Y�3S�3�v3	U3�R�3\��3��<3�6�3qJ�2\�3+A3��o3Jl�3���3��2���3��3et3��?3u�f3�g3KR'3sJO3"36E?3���3?��3ū�3��2�Հ3��[3��3��3{}b3ƚS3"F�2�:3��S3|�3'�3ż3Tx3'V3�*3��Q3�{�2�N3/(3 z�2��e3!�3h�(3П�3YE�2�jT3�X33t�3]�2��W3��2-�3��N3�A3��/3��3å3E�x3FH:3P�3�G3��35!u3Z��2�3���3�o`3��3��2��C3�_s3;L�2p�:3,�2dg�3U�3�Mk3i�3�Q]3��83L��3���2��b36�&3��3�Q3�xa3O�;3�Ɇ2��R3߻�3(D�3P>34��2��h3>[3�a3��43�Z&3��3�a�2��3ȇ*3wJ3��3�=�3��3v�&3�t!3̾3��,3�,�3(��3���2Q�:3GY�3���3���2׸�27�T3�h3�^�2�D3e�2��U3�A13Ӈ�3�*3���2v�3T��3C3�(3؞�3�Y>3���2ECg3�L]3���2t63L��3�C=3�3�_ 3C�f3���2Q3�$�3|[�24�03_��2�R3��v3���2�� 3���3��3�3��3�*3i�&3��3#�p3R.!3R�a3��3a=*3�R3j�2Ƃy3�Y3i�\3Z=u3p��2�3�E�2ˈ3�U�3ڿ!3L�3�?�3{.$3�F�35�I3S3��2.�f3hl�2��2H�23�3̓3݉�3��#3�)<3�3�m3le[3S]3A��3���2!q�3�S3��2���2 И3��n3Ҙ43�Ù3iN�3?�3��h3q��3r?3�@K3��3k<]3��73L5P3�IK3�3��2;�A3�f�2�/�3�3#�2�\"3��2���2ڪ3��P3�H3��z3�3�O,3|�?3Pa36�$3�rb3	�03�C�3�Q�3���2<��3�1y3�s�2���3i�2'ц3�)$3�3V3G3473��3�H3���2�;�2<�3
5�2I�2��3I�3�3��3�3�"n3p�3���2�C3�C3*�D2��2P�.3䲷2���2�=b3�3�$3ҏ3�/s3���2��\3�j�2��
3ш3W��2�z3ԭ3*3D^3 H3b�3V�2� 63�
�2��2�"�2�3+�63�ש2dk3��R3T�3i��2�Y�3;��2��2+n3�(39��2o�33Ъ2� 3�3cBP3�-3f"�2���2.��3=�
3+�2�}3@"3+n3�
3��2t��2^�$3WM"3�X�3Mo�2�3�H3U="3,3U$3�	]3�|�243�Č3��]3�s3�־2�33J��2#
3��3��i3s��2y�3_��2(u�2��3���3	�-36�3�b3i��2Ud�2�.�2jG�2��2p$3kXs3C�m3�@�2�2|2a%Q3903��2o�3�3۸�2�2��u3�,=3)%3v}�2���3O\S3@� 3m�O3�&3z)3Y��2�X3k��2�pL3��3v�	3.� 3�f3|�{3�O3��2��+3'�2��39��2^[;3��3J�30�3	m�3.3=�G3��3�)13���2��F31^>3��2�KO3��_3�#r3�d3;}�2��K3(b3���26�3B]c2��3���2'Z53�e(3)�D31�'3éz3��3q.3��d3�aB3�5�2��3�)E3�I3+�q3���3��W3 �\3X&3Q�3��3+��2h�=3xj�2�3^d�2uR:3��2�b�2�3F��3��P3s3-��2��A3�3�3�eJ3Z53�+3�Z3"�21�3c2�� 3��036F�2�)3c�	3dT�2È�2k)�3��35�2�Y�2�@3���2�lL3��2Vt*3R?�2uI3�3���28W3��Z3��-3��*3��2��\3˶�2>J�2���3���2@Y)3�F�2	�<3nF
3yk�3E)32�$3u��2Ⓦ3cp+3ML�2�A�2T393*<3�l3��3��c3�3�2}��3T&3��3-��2�-3�n�3�f�2&�t3|s_3�o{37�3�N�3��03�V3�yD3m�3� 3>�W3	cR3! 3�/_3��3;��3jUM3�
3 �3��G3�:&3��)3o�3��43_�E3��x3¼R3��2&3��3EU3!j93%�'3�Y3g�W3��3G�f3olH3�F3)۩3��3<3P3���2��e3��3"Ϸ2rы3���2Ba3h��2�a3��2��3Č3���3aՋ2�#3��S3�И3v��2���2��z3�
3�1P3�9�3nx_3��33��3�b�3�
<3�|�2�j3���2U�R3'�3���3�b3��13'�3�v�32B 3\@�2 w�2�|3��~37͌3)�B3���2V� 3��3���3oG3�}�2^�h3�p�3&�,3yH3�4I3F)�3bM3�Sx3ݧ�3sL3���2v��3��73�YS33�t73�'K3�]3��z3s"35Qs3RiR3�Z30ʂ3�+3��=3���3��2�e38�&3H�3L�3.�'3��3UC�34*3���3V3"�Y3�>�2���2�}A3��3�53�3L'q3���3=�v3�63��93�P�3��24�3��i3Q.3��H3z13�3�r.3�'�2��3��3
3@0#3�M3˶�2\V3��3&�x3G�2��3��3|[�37�P3�D�2H[@3��a35�J3(O�3��/3�w73z�3��3!*3�%37e�2wv�3��3�S3�sX3���2�!3�~�2<?O3���2ko(3#7�3���33��2-'�3<�A3�3�^3=3v2�3{��2�u�3�3�y�2=�2���3��03���3wZ�3�0/3$�3�T#3��3Y��2i.3D3��e3�Rx3Z�2�n3�N]3{�%3�R(3T�2�l3�"3��F3�P3�+3�#"3� K3C�U3�6�2��>3ش�3�<83�2G3��o3"�A3n�2�53iNF3�3
B53|EC3*K3���2R�43���3Y�J3���2f33p��2�Vn3�xP38��3��D3�a3��H3$�3 R,3i*3�P3��25(3q�&3�=3-�i3b3�D33H�%3 *�2��)3&93�}.3�>�2���3~�}3��Z3��J3���3��,3MON3��2q�3��3ݴ�2�/`3�;3W+3��3���3��3�r3T�k3�aY3�3��%3��J3�qr3j3F��3�3��23�V93�4^X�2�3pBB3#�^3[�2�5@3�g3;��2�3���3b�y3�ʄ3��
3��H3n��35 3�&3���2)l�3��T3��w3#�3�23�M�2Q�3�P%3۩	3�
3OW93q�2X�U3��L3�>T3$�v3�x�3%H93�3���2ï�3#�[3��2.83T��2�53i��2�a�3}c�2}?j3C�3�3�3��3�;�2C�3���2�}'3	f3�03Q�'3N��3��}36�b3#��2�BI3��3��2�}3v�3��3T�@3��3O�F3vgh3n�3���323b+o3�[13K13	3<��3q]�3���2n3*�3�3O�43���2YeG3�XF3�b3��,3�2h��3��37v�3A�3[��2�-3�߭3��3Jd~3�|�2�M�2���2sq3��.3�3�s]3R�38�U3U3�7�2��e3�.3��2�Cp3j��2ǩ43k/�2��v3�`�2�Y3��63���3ڮ13�>�3�V 3��3���2�d3�a�3��3Z�B3���3�83�=33�)�2��O3hY3�� 31�b3K��2`��34%�2��I3�}3�23':�2?.�3�	3���2���2Y��2Q�2(�E3�	�3� 3��G3Z��3�/43hF$3���2��G3�F�2 �_3%�W3#��2��3���2�&`3h�,3�93��P3/��3�M�3t�[3kk�3�M�38�l3�L3VIx3�ϊ3��3�ߖ3���3)�j3��/3��3@�	3h�3��Y3�Ѩ3��I3}R3�]4u�>3�Љ3ا63�ǭ353���3� s3/�3E�3�ˇ3 �)3��3��3��3t��3,[�3���2u,3��03�73�R3�:+3�3��M31P�3��3%;�2*tE3E��34U	3Մ�3_+[36��3,[3�\g3Q�P37q3�C�3��3�G�3��3|��2�3X�C3�� 3�'|31�
3��R3�>@3d��3�m3���3��e3X��3�!<3�M�3=dL3G�G3��3ȃl3{N�3��3T�B3u��3cˬ3�i93k�J3^s@3�/3eb�2c�(3��
3J�3��$3W��3"V3E%K3�/3�L4q83z{3w3�q�2��$3x30X�3jS3�
�3P�3��K35Cl3�3:v�3�n$3�i-3��>3e�2�k�3W�3=��3A4y3��33�K3)��3���3|�3��3�L3ۈ�3��3h�}3<��2��Y3��3�p�3�P3�uF3R��3��3�w3p�3��3���3�3zt�3�|3��34!3��4�&13 53��x3�ݓ3H'3%&3��i3]3?�U3�n�3t��3�!�3�3�=�3f3;~63z��3��V3Hƫ3RI3L��3Y�3}�93�3{w�3�$:3��	3˙33F�Y3�QZ3dAa3��3d3�x3�8�3�
�3��r3��03��4O 63��2wʓ3"3�,3��V3ݑ�3��Y30zl3��}3�}�3�r�3z̓39�3���3a�c3o\3&T�3���2?�^3���36�3��3b�D3��x3ۚ�3�B3��j3<l3�L�3�b3�b�39{y3W��2g�2��4�:37X3$q3�.3|�2.�3�63/{�2�e]3Ї�3/K3y�73��2��3�1u3)� 3c}3�S&3��!35j�2x5�3l$34�3Fm�2X](3�Ĳ2֛/3$3��2 8�2���2��3I�63v��2�xW3~C3��3kۻ2��33I��2Xd�2�à2ө�2�z 3(.3���2M��2��W3۟03z��3U�2�2�v�2�^B3���2�C3�X�2٭3D�2"�E3�S3���2��2��63c�	3���2:�(3ل�2��3Gg2��3��2�:3�Q�2��'3�\�2��3|�2�
3��23�O03�:�2
�2��3˵�3��3~�o3��2:X�2W3Ö2b��2�?�2=��2�3��3";�2:�2���2��3%q3X̔2���2E3��2s^3�j�3�N�2���2�w03���2b(3%Ǵ2�t3l&,3��2s3O��2>�%3�f3�A03��2Q_�2L��2Se3ky3�R3��03�O�2]�3:3�M�2Fi�2�[�2N�M37l>3?|3��22��2oS3�Z3cC{3Z��2W�2f�e3�p3���2���2� �2�}V3��L3M�
3��/3bR�2��2�i3k�Y3�؂2���2
��2���2	B%3b��2��3u=
3-"�2�G�2���2�G33�>3�F3�n�2�(�2�۔3�;�2*�)3��3f�2���2�L�2���2���2��3G*i3�3�+�2ug�2�C3hP3���2e�3��h2�{e3��3�K3��3bQ�2 ��2��^3�6�2��/3�\�2Mu�2�3V�2�*�2g��2�h3�W�3�� 3��,3�u�2�.$3W��2#~�2�43r�2�53��2��f3	7�2wSV3���2���3(R3�~3�I3���2��2_� 3kB3O� 3h�"3wt3�3�B�2���2��&3_3���2��2^L�2�-3H�25��2J�3a�2g��2"9�3�-�2y3��3���2��33"��2G�3�&3�23x�3ܧ�2?{v2��2�o3O�3+�3���2�S63��2�ג3���2E��2�c�2�/{3���2�3�d3^W3=�+3]13I3	3��U3���2�f3P�83�	3��3'y3k�A3��n28a�2Ï�2� %3���2Ho3�3x�G3�3�q3��j33Ŋ34��2%�3�l3��.3���2,�633�ؐ3m��33���2�U34w&3}!�3@+93s�!3!'E3j�2�&Q3>�"3l]�2��3D�p3>3��2H�3.�T3�36�j3`�:3�c�2��3VF�3��3��2h�2��e3��D3��2	g3e�2b2�2��83�py3z�3Īr3�y33ז�3%�2�
3>�_3��N3P�2�tB3�i3�8 3:�63c*3۝83��3�m3ͬ�3��3�i�2��2���2!#e3f�
3�|y3���2Q��2��%3��3T,�2[�3�3դE3��3{�73;#=3��2��/3A�p3hh73��3U��2L�*3�1	3��2ވb3�#3V'�22�3M�w3(^
3�+3 �3D
�3\/�2��3v�93�U3���2��3�3-˯2��3�u3-�W3�D�2S	v24|Q33��2z�3��}2�3�3�p3!��2vy3� 3�3�$3.n3��2��
3�3�2��=3srz3B�3
:,3v�}3w�^3"��2:4�2��F3�#&3-�3��3�S�2�kM3K��2"�o3"W!3e�3sW�2�	4=�Z3:�G3Ϛ3 �Z3@�2e83�03/��2�]i3z�3�~@3-�3@��2�Ba3�w�2�A3&J93�<C3�@v3c�2B��3q+�2A43�03=��3^�2}<)39�C3k�73%N�2�=3v3I5�2�r3O�[3��3�:3U�2�Б3>�3��3)o�3��2Q3f�22-�3��2#'3��3��3;=�2=�3G�K3;3T�Q3Ơ^3'I3�=�2/�E3=3-v�3DH43�[2V3�-3ʼ#3X�03C��2}K3��2�gz3!3vC�3���3�Z�3@36l�3Gy�3$��3�iM3CQ|3��3�=3	߄3�C�3{�3�~3�[K3c'�3��3�7.3��3i�3q��3;�3�7�3^|�3��k3Z�3�K�3n4�3qH�3g��3d�t3+3S�S3v�3�U3��]3�ƃ3��3�l4�}�2��G3���3X|3���3���3���3z;�3�Ż3ݹV3�C�3�?3�b�3�1@3
Ry3	I�3�M�3�kB3�Y3�373ɂq3q�s3��4B��3��*3K�3�E�3� -3��n3���3J�<3%��3m3�!W3#3iW53�m�3�*4n�3���3�0�3!&W3�E�3�؆3�3jK3���3o��3��3��I3�3/F�3*#�3"�	3;�n3 �H32�3#zK3���3��(3���3E�S3x�
4��P3�X?3__�3�3w��2���3=�3A��3{E3���3���3��3�X+3U4D��3谐3��3��3�Ƣ3���3�D�3xv3E�3ZP�3՚�3�ӑ3�Ml3�V�3r.�3΁3BN�3���3-�3��3�޴3��3rI�3H'-3ؠ3�{�3���2�<3B3.BA3�6�3))�3��k3��G3��%3Z,4i�3ޅ�3H�h31E3fIT3�/g3��3�=3��3�6�3]��3D3�d+3'�U3�F�3?F3�L3m%�2r�32U3NaJ3�V�3�C�3��3���3d�\3�f*3��33�B3�563��3"�3�K 3�n93=��3�L�3BO(3Ą�2Ʉ�3+3��%3uW�3���2�L�3+\3x��3[�!3d�;3��3lN4�QG3`L33�7�3�@�3R>3+�3g{3}��2V�3���3Ǻ�3琢3�#3y�~3[K�3a�?3�tV3�l�2��3��T3n�3t�m3��S3�	�2�|4 �2ա[3�_3�EU3U�3�03`>�3�!3��z3)��3�ֆ3H!|3�,3�U�3��3l�]3�K�3��@3���3��i3�h�3Ab)3*SI3���2�:�3��*3��3���2��R3�2���3�(3�3|J3�4�q/3��93��2��+3`3�e�26�e3v
3��L3s�
3�S3�%"3�33�4{3���3a23cc�3�D3��3�N3N�k3�573�3��M3�x3�o3�D@3�!�2g�3�^3&?*3fzW3@�3��i3.F3mdq3�9+3�c3əP3,֚3��C3��Z3��e3˞�3���2�g538�3���2��,3���3�t&3p�T3�T�2}��3�{G3([�2��G3?6,3�r�3P3翁3��D3�q3S�3���3G��2!c3�~y3��3:��2e�c3�!�3ծ�2�F/3Ǩ�3mz-3)�3;˳22�3�l�3r3?CL3��3`
Y3�d�2��3]�$3'�2-h"3��3���2'>R3M�3�~C3�=3�=3�5D3f�2?3���3~Z�3��a3)A)3�"�3[�&3R�,30�3J�2υ~3�V3<�i3^�33_3��3�^�3D�I3�~B3�c3�
j3m�2��I3�TH33�33N3l��3�(�3��2V��2ی3���3�P13��Q3��C3�BU3//3f��3FTN3�`3��3k~�3�*3�r3ך�3?�[3�2o3��3�I�3�23�=U3�04��x3/,3��3`�3b83��2�|$3Q�3n}23ٻ�2PL3��3ZG�3l�13z��3,�
3q3zG3�33Qsc3ϲ33�̬3�� 3��{3�l�3k
s3�l3�'3�H3�3�03��n36E�2�R3��2�m�3/�3��E3jC�2��4o"34�3��3�G83�4�2�)3�~Z3���2��F3�T�3�JW3�7�2��83�F�2S�3]�
3��P3X��2-Mh3��2��p3�}�22,�2�@3<3�3���2�[[3��;3��-39G13��P3a��3��2� 93K�37i3�|�3��2��S3[�,35�.3�dg3��2�C�3��3
o3���2�V�3�CG3!��3��>3��y3yr3܄W3�2�ޚ38�O3i,)3ͯ#3�>�3_�\3���3��2�l�3�ނ3��3��'3<��3�;3w.�2�,�3�D3��N3��3���3"�J3M E3��j3��3�<63F�3>Ҋ3&�53.Q_38W3�v3�{�3��3�w3l�o3I|_3f�,3�N3�d+3��13�7�3�O�34fu3[J 3��3��A3���3�3n0|3S3��03�Y*3�*�2i>3 ��3�0�3���2kϲ2�oK3{B?3��43nI�3��73Ae^3	��2>1�3YW>3��13
3���3�Q3��$3�Z;3Q�3���2�y3�k�3]Z3��D3�'�3zf�3�}93�3��]3F�3"3F3	��2��D3爧2-�3�;3/t6333�2#ԝ3��s3 �i3:�3��-3��$3#@C3z�3e�2��l3��4!83�3�R�2�ʇ3X�<3�2%�3\;3��K3��A3n+u3�3#tQ3��.36�3"T3aC3u�3J�@3�}C3m�y3h�3|��2�b�3��3n:|3(�D3s�2~�k3Ňj3'�93��3`�
3�V�3ICK3��3Xh�2��i3��#3���3�236�@34�M3�213�JS3�=3�Վ3�73���3{�|3��36�2���37֘3O��2��.3�"73֟�3��3 �3�K3X$3��A3���3�13v�J3O"3��h3]GK3V�e3��s3^D�2�<3P9w3�S�3��j36��2��.3g�=3��
3��3lv3���3��L3�53�m[3��W3��3U[4b��2B
-3���20 3��3��q3�)�3-3�?3��3�ڐ3\�G3Cp13�t<3H�K3��=3/'^3�U3�
Z3�0]3��i3hl"3:��2�E3��3@'3R3L�%3��3%=3��'3��M3:�
3�;�3��z3�\�3:n73��3v(�3��83�FI3�xa3�]�2��34��2x�<3*�L3ay4�T3�'�3LJ�3α�3��3>��3:3Z��3Lk�3$�R3�_y3�#}4w�3ƾ�3�R�2D&�3K��3��[3��l3A��3�e�3(H�3��4��33O�3>E"3��4�43��3�!D3��35K3+�3t�3a-L3bh�3�<�3�x�3��r3�i3���3���37j3b.�3��|33"`>3�,�3�r3�[�3�(31��3��3��S3u4�3���3Kv3��Q3��93?�z3���3��#4��33��3�\W3潁3�#537g3%�13S��3b�3N93cA4��3w,�3�Ҵ3�n4sOU3��3Lͮ3NJ�3��3�9�3ua!4;�3�S�3\�4�ƽ3��x3ܠF3�7�3	v3�U"3Dp�3��s3?M�3�W~3�s�3�3ߴv3\aL3Ȅ64��3�L�3�}�3$�&3�ѩ3Xk3#�3���3�X�3�9�3���33J�3:t3ƀ�3�%�3y8�3�$C3C�*3�-�3~g43l�3�|13j$�3i8v3{84v�c3��k3d��3�KP3�3f��3�;�3n��2�Oz3M<,4`�3ؕc3z�3,`3���3��3���3Y�>3�	�3F��3|S�31��3_t�3R>3ښ4��~3!�3���3%��3!<�3�3��3���3��4�m4�$&4�zz3��3��4m	�3I-�3m�3��>3�p�3�"o3���3��h3�x�3k[�3�&e4)" 4�Gd3�37<�3m�x3��W3��3R�m3�h�3e4WK4�|�3�:3���3^��3�l=3�4�3ޮ�3�z�3�k3?��37�j3䗠3���3��4�l3s�30T�3��Z3��3By3x*�3G�~3�,�3���3�ޮ3���3��r3��x3py�3�3B#4k|3�3�<�3��3d,Q3!Hv3.� 3�Gp4_k3�t�3K��3��3�A�3�Jn3���3�2	X�3�24�3Bm3�mB3��3�R�3Ǖ�2v?�3��
3P n3E�A3̦�3�+3�3�B�2��v3Z�73��Z3�	C3C$3��3"�3�3x@3\'
3!�.3xb3�*3�T3��(3��A3}5�2?�3�`�3(33��2��D3�`R3�-,3�,�2�,4���2�N63Ӷ53��3�3�+3$}	3��2�~F3r��3��O3�!3�t�2�w[3��3Զ�2�3���2�-!3��3�c�3R*3_��2��3v�3��.3@.�3��83� �3�t13�DJ3��}3m�+3�/�2�sp3�43� 3�c�2�/M3L��2Q�2�}D3[��2\�2��3�|(3h>3�ٿ2��2�kX34��2�K30v�3�3��3D�)3�3Z3�2�B3OH�3x�z3��?30�2��	3*�H3�cH34�3�k�2�6u3�R3H3�F�2�p�2�|�2�3�!43k53Ǽ73'-3��13lqG3y�H3}�2
.30��3zw3#X-3O\�20 3�3Σ�2X�<3�e39�3�WV3&3��2uñ2t3���3S7�2b30�33�m�2��2/�3E�
3�2��^3��3	]�2�x3���2��33ԓf3�^3��'3�3�[<3��3T563�3�2���2�g�3�3M��2A3�T�2�yF3�Z33H:3��2��P3�]�3|�I3=L�2>2Sm3L�#3���2�3�%�2D�U3Ҁ$3m\Z3�B3���2�1G3w��3yu3Ջ3V�Y3\��2�,3�O3�v3k2�2/]3�P3	7e3�Hd3��3n�&3�@(3%��2�u�3�3:d�2&23 �73ں63m�"3J|�2��3�e�2�3 �B3�E,3c3�
Z3ۺ\3x3�2��23L!�3�638Bh3G9�2��3��m3@}3�3oI�2�a�3���2ah3O3-�2p��2�M�3��3S�N3��3�73?��2nG3M�03U#�2l3](>3�XK303�2�3V�=3?B�2T,3���23LZ3���2��>3��3(4�3��b3�9�3Q�3y-S3/�63��36�3�3���3��,3]��3���3���3"�3�D�3���3�k3�K'3jE3�ڎ3�kt3��)3l3�3�U;3�p�3��y3�34w`3=��3��3N��3)|3�E�3^��3܃]3���3 J4�B�3��~3�_�2���3Ƶ�3n�N3�Y\3��`3�q�3�:3���3���3�5o3�u3��	4��\3�t�3��3�d�3�P33��?3��3Q�H3l\�3��3$�3'�S3]�.3Kwv3Q�n3q3
�P3�U3G��3�vA3
e�3϶�3}f13�%3�54-�i3q#3s2T3S�a3�7'3S�3[.�3�x3�=�3å�3s�k35uX3f�2��3U�93�Lk3H<^3��s3�\3�hr3�g�3tc3]�3�}�3�.4��3���3~Ү3��u3���3�y�3Ĩ�3TH3vE63?R�3��3b]�3�p3'J�3ǧ�3��3g�e30}�2�V�3��3Î�3;J�3��3�B3��3�<p3\(�3t,�3��;3v�/3D��3%�3u�*3n��3�u3���38��3M�3d'�3?�3�f3���3�'S3s��3G3 x�3.23m*�3�63m�43i3�u3��3��&3@��3�3���3B�l3���3}\4�eu3&A3v�=3��3G3�<|3g�3�l�3	3�!�3B�4�O3V�3%J�3�4!}K3(�`3�y{3��;3h*�3�!�3�̘3�D}3�{~3��3f��3�\�3��3��3���3^�a3��3�[T3�|3�m3˗4�^q3�P�3[�3��35�3�Z?3�$�3�k�3X�3)h{3ؽ�3oU'3�є3��74#�3>_�3�43���3�1�3�T�34��3��^3��3[7�31��3'B�3MaN3MZ�37"M4�Z73�~f3�V]3N�}3�' 33lx�3d��2��3��3K�3�b�39� 3킚3�+�3 gC3�3��3�5�3�/3/R�3�k�3��3��2�i30�!3@qI3'�3�/3���2�yk3<r3��2[�3�3H�3��3.>3z�;3�y3��2a53��'3�@3K< 3�[3'43\] 3�N3ZN3�[3�EF3030~3�23s�73��13y) 3�|3��H3��53/�2�\�2`3N93�.�2��V3�v3lz3�n/3E.j3���2��2��3L/�3]��23�3��43a�3��2N�3���2�93�a3�)�3=p�3S�2.�2�e`3�Z3�3|�T3��2+j30.3�}3��3��E3V�b3�e3=G�2�*3TG3�e03

3J�03]4J3�ͼ2�I"3.5�3��Q3uo:3gi�2��)3O.3�Y�2l��3
u�2�H3�4373�63	,
3���2Q��3�3��h3503�� 3��(3��3K��2��2�� 3?�3q&3:�3�e�2�23f�3��2���2C�2|}b3L3Rb3A33k�3�.3A �3~��2��/3��3�*A3{�2b�2VZ+3Uj�2T�?3Ȧ}3��'3Q�20J�2��r3�Y3���2��2Y��2��D33�13k��3l��2��3zn,3OL�3U 
3��*3:��2m�3l�3"�2S��2��2��`3�0�3ؐ+3�D3�ݹ2�bK3��3};3��]3�"�2�*3�-�2�3?��2�m'3w��2�P3!��2��2�.3
y3%�,3VT3��)3�3�`!3(o�3��c3&#	34u�2��3���2b��2"�X3���2�(�2�%3�F3c'�2�3I3}d�3hG'3�]3s�13��3	��2�C3&=e3j�2��2&�3P�3��23���2��23�C�2:3���2(�:3�&�2��3�l3�33O�3���3��+3I�3��2�R�2Y��2n�2��N3O\�2��>3B�p3歫3�pB3_w�2P*3��2��3@ޜ3�[�2��#3�?3^2T3�ld3�h4/�3~&,4ޒ3+Ӥ3O�3�W�3�B3n�31��3t��3�7s3BF4��3�ۮ3$�3���3<�3x"3�&3���3eNV4��13�4>D�3c�3q�3�M84��3*d`3xp3���3s�C3ϴ3T�B4��o3ʿ�3>�4�%4Υ�3�j`3�A�3*-�3Ql{3���3� C33*�3�W�3�=
4�İ3¿3�	:3�4	�{3v��3�5�3P��3ɿ�3���3	D�3�+3y��3	u4y��3�޽3)�3�x�3�Yi3O3X4�$3=��3@G�3�4��3��3[n3HbA4}N;3�c�3Y2�3ě�3
��3�޺3(�3ppF3���3U�4��4�I�3��U3=V4[ר3�jE3��4Xe�3>�4��|3��3}��3���3�!3F�4} �3@[�3@��3��3�Io3o�3{u�3
��3*�3i24���3n��3��|3o�4���3?>t3�$�381�3��4L�i3�<�3g��3�/�3���3�<4$l�3V�~3!ʭ3�1�3���3�K�3Z�3ϓ>3iTp3�b84Ͳ�3H��3M&�3}�3��3͇w3$\�3u&3��84eW3��3�|�3ޤ3�O 3��'4�q3Xu�3�4s�3A}3��3�34^��3g��3t��3k�3Tj�3�kv3!4�3�ǡ3e�3�͎3m�B3�<�3
χ3��3���3m�3��K3Z�,4�j�3i/�3���3_x�3�2�3���3�N�3��s3�4�3�R.4� >4���3,�3Q��3k��3ae�3,w*4X�n3��3tӕ3+�4���3&��3�l�3X^`4�g�3���3AҨ3!	�3O��3mG�3ai�3��3!*�3b+4�'�3��3,��3z�3툛3Բ3k��3@�53���3��I3Ĭ�3�@�3���3'�3~�)4K�83�#�3c:�3C��3So�3�4��4��f3�8�3Q��3�1�3 Z�3�Wr34�0�3�R3.��3"ލ3ɭ3� �36�4c3���3�O3���3��<35��3PP39��3��3��3,w3c��3���3cV4D��3�Y�3��.3w��3�(�3���2��m3iu�3�>�3Sg3�ӭ3F 3���3��3�U�3=�S37�30�43	��3ĒQ3LZ�3<8�3U��3V��3h��3SN
4m��3��73�"4�u3��X3�/�3D�3�yV3���3��,4�X�3?)�3�L�3���3��3:w�3���3��C3iM�3`�$3a��3�,q3f��3�sV4�ļ3\��3F�3.&�3��3ؾ+3��3Iˣ3 _�3ח|3���3���3:��3x�631 423�V>3l|�36��3CW3���3��4�� 3���3y�141�k3\�u3�73���3v*�37�=3���3cLG3�g�3%�B3���3���3{�33q�3diC4=�3F�3���3�B�3��3)�k3�i�3}�>39V�3;@�3{P�3��f3��63�Ϋ3C׃3.34��3̰53��3��m3���3��3h[�3�D^3b��3bh�3Ͽ�3T�3u6�3���3�8�3~@�3��3E�3�'4G��3>h�3�g3C��3��3��3LF�3E��3���3�f43��3��a3���3�3��	4zu�3gP�3��x3�d�3|�f3�4�.�3�|3B��3Ip�3p-	4��3ܲ�3N	�39.�3Љ�3P�3l�Z3�b�3�23ۏ�3��3���3|w�3��3��r3�S�3�	h3M��3�u'3���3C0�3d3J3ש�3y1�3c]�3Zl�3�w3b˱3k�3Q7�3ų3�8y3ڥ�3(N3	��3Y�93cZ36�J3�A4~,�3P*O3���3ݼ�3�˅3�8�3���3|bc3z��3���3r>�3_�3�y23s��3㊅3��3��{3Զ3%��3C�3]��3ա3��N38�q3F54��3=�3Œ 4 ��3�}z3mő3�A�3�*3^M�3���3��3�4�A�2ݟ�3��4oo�3�-�3��%3
��3h�3(�4]3�3�R�3כ�38��3X�3y�p3��~32�}3k�:3o��3'��3Ot$3�-3���3��3s�4�Vz3���37�3$43��33\3��h3�?3霘3��3V6�3Lp�36[�3N�r3p��3T��3b�3j�_3x5�36@�3f�b3��3�4a}�3Vֈ3�/�3��B3��Y3��Z3�I�3Y3��z3�W30��3cN�3R�3QK�3o��3��K3�Ӟ3�%�3��4Q�r3?�g3��36GK3�33�4��4�3�oB3ߍe3?g~3/j3�3_3�"�3�124gԀ3�
4:L�3O�g3,1Z3�'�3K�a3��M3?3?'�3Є�3���3���3��=3(s�36��3�e�3E<�3�p	3���3"�3��g3d(�3peU3���3�<3���3��3F�c3aP�3�4�u�3��G3&�73"��3���3��3an�3��R3��[3���3��3�h@3��.3���3�|�3A؀3�џ3��n3�#�3 ��3���3��3�!L3��3bU4���3YV3 #s3y��3�3�E�3�0�3}6S3B�3�4�:�3���3)[O3)~�3�K�3�i3��q3��B3��3��d3�{�3��3��_3�G3�N4���3���3�a<3Y�3���3�6�3��3��3�ٰ3k�4-��3x73M�,3(H�3��3�M3
��3.zc35j�3�.3p�(4ۏK3�7W3V��3S�*4�D3���3c}�3��3d,I3Ť3���3��p3�ڴ3wW4-44� 3�334�b3��e3���3=-k3J�J3.{H3�>4���3N43��3J�46$x3m��3�p3�4�36=3zA�3��3-��3��3.�3tJ�3uҘ3`D3{�3��3@{�3\��3�s�3���3e�38s�3ӣ73A��3Y\3�L$44u3y�?3Қ�3l0�3�L�3x.�3���3�v3��3P�_3;4n�T3��'3�m�3��=3&N3e��3�R)3cE�3eҀ3!E�3:[r3;�`3@�3o�4e43f�3�H�3�f44v;y3�$�3��3�0{3Q��3�-
4�3#��3��3��3��3�s!3w�p3s��3�*�3��h3�٠3���3�OF3c��3e�3�ba3ɒ�3\ι3Z��3��03���3Ȃ3��q3k��3.vR4t��3!�4�9
3,� 4K;�3掕3��3�׈3.t3{�^3W"4��13�O�3��3s+D4�}�3M^�3Ϲ�3c�4w��3Ņ3~� 4�Rh3xі3>?4��3+�}3�T3]�3~��3h��3��t3�'r3���3ɍ�3��3���3O�a3�h�3(�.4�``3vÉ3%ӡ3��3�Yl3���3`�Y3�ݎ3`��3}�4q
�3RP�3��\3C��3��3�1�3^�3gS3�7�3ה�3��4_HT3"�P3b�h3�R4˦o3�ق3L/:3�}3�Ԃ3���3�*4Ӓ�3x�3�4���3��3΢C3�m�3~��3�(�3�ݥ3�pB3 *�3m3d��3� �3��t35�3'�4��3δ�3��T3�m3�R�3�{�32��3OZ�2+�d3�\4���3�S�3�G3	��3k�3,#>3���3�x63K/�3���3]A�3�h3zx�3�v�3��54�Ȋ3wߣ39t3��3fq�3hq�3d�3�?�3���3�24��4��3ꊒ3���3��3�qp3���3y�z3��3ɴ�3�4��3��p3��3��O4q��3ĉ�3u
�3Vra3}�S3u�\3L�3s�3I�3���3�6�31\�3n�U3���3u��3�
g3���3�(3�ŋ3jXJ3q��3�l�3��\3�\�3���4m3�*�3�v�3�3773)��3�<�3�;�2³3�Qn3x��3٦�3�#43���3�T4V{p3/��3�H3#��3is3c��3�wu3F�3G��3�f+4"@3�3�#�3��3z�3�.�3'/�3r|�2U��3& �34V`4�m�3�D3XLp3H��3#�@3�=�3�](3Ԥ3	]h3+?�30�3Dod4��4u��3-�4Ct�39��3_7�3��p3�9�3�/�35 �3{>j3<��3s �3���3�!�3���3��3Ql3�4�3���3d��3�Ԓ3��4/^4k��3tE�3��)4���3�K�3��3"C4��3u��3��3��3�Rn3��3}�3��3$�S3�0�3~��3��3p�3���3C��3&��3N=4���3X$�3�e�3�	4�r�3K�3j4�3�:�3�l�3�n24fL�3G;�3-C�3��4m�3<^�3��3̼�3�l�3[��3�3�3�M�3ɟ�3(�,3Ƶ�3�Y�3���3XS�3{�#4�|33�3��4��3w"�3ŗ�3���37c3a��3�� 4�4���3s��3r��3r�4r��3�3,[�3P8�3O�3R(4�V 4�Q�3r�*3��~4���3�c3���3�p�3%F�3��4���3#{3��3@� 4/0�3�>4��3���3�o 4�f�3d��38�3T��3IК3i�54���3�[�3�x�3\a84�L�3#}�3��e3s�63q$�3Kƌ3	��3"gZ3
�3�\94�`�3$y�3p�037��3#�3��3�Lg3VZ3��4#�t3@��3!%�3;S�31m�3@�M4&�3l�3�S�3k$q3�}�3{�3�34���3���3�Pf41�3���3��y3B��3KS�3�4�g4��36q�3�\�3�y 4%$�3���3wc3% N4��B3���3��3{�\3m�3�L�3�P�33�q3JX4=Q4;M�3�n3[�K3�4)c�3	�3��3�-3N��3*�3��4��d3��3h��3��4(��3�`4S�3��+3�j�3p>�3|֟3f��3���3��4G�3��3�Ht3�Ӱ3�V4;]�3�Vu3��3��4]U3�x�3�J4*�33��y3jG'4�N83��3j��3��3�1s3Q�Q3���3)�?3oC�3(��3s�3�o3�L%3��3���3��3��3}�+3E'�3�)~3�� 4��3<�4'�3
�4j��3�*�3*��3]�3�{3��3��3i��3c2x3��4u[�3'}�3��3Ӛ40�3h��3vSX3��f3 �r3q�i3�˼3��3d��3�ʵ3��=4��\3�<�3��]3j�3��h39�3��3˽�3<ً3�/
4vH�3�Ci3:��3���3��3D��3�(�3̸�3�c�3���3b'4<kj3��3Z�3X* 4�[w3�4�3��3��3�΁3��3�%�3�:23�C�3+�4��4+c4+�93��3�
�30�43Վ�3q�43$� 4�d]3���3���3�j�3C�3�vF4E�\3��3�͵3i�3UF�3��3���3�EB3�36%4ƴ�3[n3��3W�3L'�3W��3��S3e��2�h84��H3(4�3���3�3�ʟ3b�4���3��3_r	4�j�3\0F3ڎ�35��3q]T3�3��3p�4��p3�i3{%�3�\�3}R�3���3�On3$��31�r3�w�3Q�D3��3��3#_-4�n�3vbi3���3Uf�3e~�3Z��3��3�G^34�Y3?��3g�3I>3Kڏ3g4Z֘3;�43��3��-3�5�3���3���3���3�#�3��t3 ]4�3��3}Gw3iԱ3*/�3E��3�~�3��3��x3��4��3ן3|�3	��3~ܒ3c�3Lo�3��h3���3�I�3b�4�H�3�ī3�3��4e�U3�-�3��3]N3�V�3�+�3W��3=I~3���3���3[4(v�3(O}3���3`ў3ދO3Tص3��<3Q�3)�3FP�39zr3�Q�3���3��C4�G�3a��3@�3U��3��3��o3�Y�3̱)3�C�3��44��3r/4;e}3���3��4S�3�T�3��3K 4���3�lA4�b�3��03�BP3s�4��3{ �3���3�,4X˄3�;�3�3|D�3&�3���3�s�3�E�3ŉ3���3I%�3%�/3���3��L3~�~3#m�3�4�3?X�3��}3�,3�|�3��%3:�Z3ե.3*?3�3R�3���3D�3��B3��3��u3e<�3��^3Q��3�7!3UM%3�5*3�Ji3���3�U3m=�38�3]S93��3m��3-i3̍13�_3)�O3�+G3M��3�Ŷ3�[3��3S��3n�3��3�
3�&�3EZ�3Y�'3Ui(3�83-�3� I3`��3KH3Ҕ�3�]d3ς�3 OU3�d3N�3+TZ3� �3n�C3�(�3���2�,s3&j�3�m�3��3䏕2���3�Hx3I73��H3mL3�{�3�?3�B�3�+3��3Z�c3�m.4f'334�F3Ή�3�/�3b�n3d��2��o3���2�v�3�E�3�W�31!G3c�3��H3F8�3Nn�2�fm3D�F3Sː3p��2��3�403y=D3l�3�ߨ3$9�3+��2�2d3�3۬83S�3<�y3`3��[3]}�3kT`3	qo3�o 3�aK3>�3�d�2�S�3��J3_�W3�3!�3 �Z3��36}3�$4ޘ13�/<3!��3�t030Lt3�=�3�ѧ3�j�2ͥ�3�A�32�3�kO3�ە3�|�3?�3|U3]��3H�Q31�3�qq3��3(?3�a3��3�(64&|�2�Zn3���2Ҵ43��]3 �H3�?s3�3 x�3��3��3n�!3u3:�3�Y3��#3�o�3���2E�f3��l3,��3���2�r:3��[3��3�b3ߢu3��93�B�2�/j3S}3��#3t�53�xm3h�3�0�3|mm3���2?�3LM�3p�"3���3.'3�<�3��3��x3�!3�W3�g3���3���32�13�<q3��e3�d13��31R�3Y�&33x�3��4`|�3���3y�J3؆3<j�3bh3�U}3��2d�3�K3*�3��j3�3�%3bt!4p�@3S?�3��3��y3E�3ٱ]3�t�3�D3k��3�>�3�5�3^�3���2:�3-��3�w3�5F3#73cP�3J��3���3��3���3�n3��3h�3F}@3\�3M�3;}R3#��3a��3��2��)3�|�3F�3��x3R�F3wŪ3k)83�K3�3�_-3��u3�d�3�"�3�d3�ׂ3YƊ3c�3R1k3�ź3l�3�hs3��3�O�3���3���3\Jf3�~ 4+��3P+y3H��3O��3�K�3i��3U��32��3�ȴ3��%3ߊ�3�;=3�4��3�4�d3��3Ad�3-ń3c'73B�N3�n�3}�R3ߎn3V:4�/�3	�?3L�<39��3�b�3�/S3�'�3�F3eEi3���3�k"4?�T3�h�3��#3���3Z�3�>33ڂ3�,3G�>3��36X�3�Z'3F��3�43;�3�$I3S@3b	�3_��3�!i3�@V3	�E3�%�3v*r31^�3�(T3:��3˞3@��3��3xyr3��3�H�32�3���3�[�3�713-'�3�#4��35:3)�i3�{�3�2�3*�!31l�3x�3���3��3���3ݿL3�o�3	
3���3�&S3?�3M�)3��3�]P3U��3�3m137�33��3��3?�P3a(3b��3��3��x3_4N�^3�`3vW3���3�}3�j�3D��3#e84IY�3汛3��+3Vk�3 L3�σ3!N�3S��3�-�3�N�3dl�3t�q3;[3"X�3
5�3�CU3���3`��2Q�S4Â�3���3��3Xח3�83IW4�d�3���3��3K��3�.`3�p�3iy�3)XG3���3KF�3�2H3G�4���3+��3���3�z@3�[�3�c3���3Z�`39	�3e�33!og3�#D3��U4xQX3��3���3�A3���3��3)�3A�s3�v�3��3P�3��<3$�K3��u3�@3�)3��3IB3� �3�5R3�1b3,ı3Mke3�,o3��B4�v3���3\(i3��M3�o^3��3 �h3�tJ3	�3�X4�#�3Caz3m:3���3��Y3�t43��3X�3bά3ۋ3xu�3��3��2�ݎ2���2D�2�h�2��3��93CТ2o��2Ġ�2=��2]�2�	�2��3Ƃ�2:R3'%3�q3��"2���2N��2���25��2�B�2B��2�P�2�=�2�v3�ݫ2J��2��y2�6�2�3��83�q�2q�2�]3�Q)373�2,Ѽ2H�2ك
3�s�2)޹2*��2aP�2_X3���2>[3�3�2�X3��2��&3��2� 3;�2��+3d��2A,3P+3[�V2u�r2*Ҏ3�� 3�њ2�7�2�]�2\�3�ù2�@�2֩�2{3x#�2v�63;��26��2A��2K�V3�{2,`�2S�21�2!]�2A(�2�'�2�n�2s�2��?3:�03��2�C2���2��2�Z�2x2%3�X2�>3!iq2��3�_�2�@�2䯥2�uo3�e2h��2�73;�i2���2;�2},�2�(q2�'3��	3�P3f��2��z27�2��P3o��2���25q�2#:�2���2$�)35��25��2zC3*>|3��29�3֨�2�'3 ?�2�t�2�2I�2���2Xz53=~3��3�u2���2I@�3�t�2\O�2w�v2@��2��26��2</�2�2�m�2�ޜ3���2Q!�24�2*r�2v+u2�H�2 ��2��~2}D�2�I:3�36f27 j2�L 3ι2"�2ǻ�2'�2�
3p�Y2�.3W�2̭�2*1�2��3,I�2C^�2p��2�73{]�2��27�2���2V�25N�3���2�_2���2�w�2�G�29e�2��2d��2��2�-�2oA3c��2�+�22U�2�q3�e�2_��2���2�S�2�=�2tB�2A�'3A�2�B3,�*3���2�3ik2/��2F�2O��2�Ѝ28~2��(3]��2W3,(3�N�2'��2?<#3dU3�&3�9�2�J3�e�2,��2-r3�7�2y03"�R33���2]E|2k��2 I3�N�2^3���2L�3B�{2|
�2ٯ�2	Ț3��2h�34X�3�p�3�R3���3�8o3^��3�
q3�"73cO53���3�A�3�$�3es53D��3d��3�13r:�3 �I3wB3m�3��3h�3�Z3_�I3[��3p	�3���3n�P371X3x*=3X_�3�3���3��3��]3�4�3V�d3�sz3��t3���3��*3�g3���3�A�2�"3��3�33��38�3Z}�33O�3�_�3=��349�3�LJ3��2C�3��3ӡ93��3f2�3��U3�f�2;p�3��3�<3$Y�3z:I3�X�3�q3F_�3��3��y3�3�!�3�z3��*3��3�^;3��K3,+}3^�13:�b3�̭3�#4in�3��=3�#�2tڟ3@�/3�@3�w3��3�`93�$37gm3��L3�>3C�3(�
4t�3 �3���3/�3�OI3/U�3��3*�53�v�3{Q�3��3Zه3��P3Ě�3T��3�.�3��3��3�e3�R3Pܭ3�a3�5�3���3j674p32�l3 ՙ393z_3���3Ԓ�3��3��y3�4��3U��3<�33���3�*z3�[d3ā�3��"3�]�3�z3�Ӕ3 OP3Q8l3(�3	Z�3�S�3;�3(
\3���3�v3��;3V%�3uk3�3��3��3q�3)s63���37�X3�i3%qh3)�3���3hͭ3K{�3��3�3r3,�r3<e�3�Y3�5p3��?3�Mg3�43�Q3���3�]J3�j�3��3">�3;Ӂ3�u@3*)�3�<e3�aU3���3U��2�-j3�s;3��3��-3��3ǀ�3�4Q
R398j3d-�3��G3Γ�3���3�1�3�3�4}3fb�3$��3e��3�&J3+ȍ3�Bx3��X3U]f3�U3%��3T[a3E��3�c3|�%3}f'3�x�3���3��R3`k�3;.3��v36�>3J�4�2-3��3�3I��3� �3xN�27s�3���3�TZ3a� 3�83��3�V3瑉3���3W?3�̉3?��3݄3a�x3�B3s�3ف�2��03x�3��	3��23{T3'��3��U3��3I�13�S3Ad�2%}�27G3�:3=�3O+<3Ӝ3�mh3��3��3�w�2]�3A3F^83c�2�C53�!3��2y�43mK3�H36)3�t$30>�3���2�!3',3�I	3� \3�2K�3@�3��Q3Z��3�Y3�8 3�3��3�j3�^3.593=�q3_��28V3[k�3a.�3�nc3���2 3ѓ�3��2�^83u(�2c3�B3C^3�0]3ES3���2ܖ�3��f3�3pPG3 g.3	a�2���2� N3���2�3(;v3,35�3fR�2GO3<�_3��2�j3%G3p�3;'3�|D3J�d3pO3wmY3��3�3�3�0@3��2�g3��$3���2��2 �A3.Ҍ3�rt3@�:3F4�2�o3hl|3ƿ3�[W3�3��)38f3��l3�P73V3�u�2g��3��3� 3lO�2�n3r��2�S>3yP3�!3�(3\L3��u3Ί�3Ť�2:=3=Ŏ3q83�<3j�23t�J3}3� 3y��2?�)3�:�2���3�7�2�7'3g�V3�V43$ "3_�C3�'`3��3��3f۩3CVb3�3��2<�x3���2��3wgB33��3��t3 %3�"�2�m3�3ef�3%�3O�i3i#3;x[3c��2�L�2{�3�ȫ2�L3��3��3���3�3 �2��S3'�2TRS3��3��V3k��2%�3"6%3�)�2kڻ2���32-�2��2�se3<�3��2\D3�B3�R	3��<3���3M6-3��3,3��(3T�X3��3݇X33�3��3��2�/�3t��2v�22��4;3��Q3��3~53�^�2�Z~3��$3Y3M�3���3'��3ɯQ3XU�2�(J3��^3_�33ds#3[!=3p��3���2~�3<8Q3k��3���3F��3�i3,�3��2��w3�|�2�Î3�	3�*�2�3��3b�3X3N63��S3��23װ�2�G3V�L3��Y3��3>e3�Hr3�[}3d]73s\�3+b63]��2=
E3i�3��3ρ`3o�M3"�2�D�3��3���3Fh�3��A3ד�3��C3:�2�e3 "3Ӛ�3��'3]04J\3��3'3"N�3�D33�g3�3:��3;�~2Nc3��L34Q3��H3�{p3��3�ð2�R 3� 3.93}U�2B3I3�G3��2&ϥ3���3�E3�m3q��3�Q3�%3#�2���3;�2h^3���3��3�g32b�3��z3�83�2�a30�O3��W2[�,3Á3��C3�wE3w�4��Q3�	3�$3~&4�@3��3ىU3833�C3��3F?�3`$�2fL<3M3�3�f3YN3#3�
~33�}3��2�;3zO'3Cs3� Q3h��3Aa_3e&>3���2dM�3A3�^:3;�3�+�3��=3��E3��3|I3�mE3�u�3���3�{�3l�2�g�3�m�3�Ǚ2��3a�3k9I3�g�2քZ3`<3Vn3�'3�C�3ID#3j�63�p�2�rR3J�3G(�3}��2ŪR3&�3h��3�Ju3�23Z3�Wa3ъ,3Q��2-�_3�gH3�J3�3���3 B#3:�)3��3��3�>3]c�2X/P3,53og3�
�3���3��73 3lM�3ۢo3�G@3Z~�2d�3d%�3�O3b�u3��3g��3=
3I�X3v�=3��H3 9m3܅63�e�2�!k3��3��3�wV3��Y3;ha3�P{38�n3ܸ�3��3x��3��;3Q�3xg3h~�3AL�30�23Muh3m#a3"�3bR3��2/k�2T�4s�3�N�3G��3Kۑ3o�3|G�2q4%3�T3��3I@�3�N�3Ž�3h��2��3^�3/r;3�OQ3���2�E3��3�m�3"O3k�Q3�s335�3uv3�6�3�!�3`2�3�623��3��x3�b3e$H3=�3,�3@ܞ3��)3�ב3f�3�	3!03�D03��13�[G3�ny3�h	4�&�3v{U3H��3D��3�Ҧ3��X3eB3��U3�N�3
V�3aqX3^�F3S{�3$-�3�ī3��C3�E3�"�3V3��c3�؆3'��3C.!3�*�3[�u3V�3�T3q��3��3��3E	33��(38�'3�:P3�Td3]a	3�=�3�8%4z�3%�t3V�3��|3�sO3��3��3�M<3,��3S,�3���3��3&�f3��~3��4�!23k:b3�u3>]3F��3��3X�3o�3��3|��3V��3�K^3�f3�.�3�^�3u#E3#�3�<i3&0Y3{_83��3}	�3�M�2u0�3��(4D�G3�h�3�@�3��^3��3�\y3\M�3>i3�إ3L��3���3�{�3sf
3Ɉ3 |�3XTv3��!3
P�3��3��R3ͱ�3��{3e"N3�3�4b�3�8G3�Y3�ԇ3�h�3��=3u�3[�93^�33��3���3�^3L��3�O3+�3�3
��3� >3�T�3�ɑ3�i�3��-3�U3B�-3�	4���3��3�D3s�3�"�3ܝc3�f3�x3 ��3X�|47إ3�03�3� �3���3�R�3Ғ3�f3�/�3I�R3��$44�b3س�3�і3��64��3��3�E!3�^3mr3:��3^�`3e.�3?��3�Z#4 8�3�O�3�u3���3�)�3��3���3v~�3 ��3��Q3��4� �3��3uB3>�31l�3X3��3$��3��L3�83�*<3�Hd3=L�3���3�^�3%��3��3J�D3>)�3H�q3��z37at3CU"4~I3�y�3��3��,3Ʒ�2�E�3%3L�s3�&v3�*:3��2�ߡ3���3Y��2pg|3�4�2p3�>�3�Q3�ٸ3�[3��Z3���35{ 3y�}3�3A��3�D+3�X)3��2�BX3=23b�2-4�2Dfs3���2*O3�403ys[2���2�&r3�^%3e�'3��2�/3��3�v�2I`�2_]N3n
.3ٌ�2�{.3\�3�M3�<R3*�3�$3.R3z�;3��+3j@�2�L3m]?3-Y
3��*3��M3�#z34�z3�Y�2��3���2W3$U3�@�2[�83�E|3�$93�3��3pq�2B�3�	�2G��2S��2M43X�w2��?3�gh36�3�ǧ2M�:3şX39��2��2��#3���2Wî2��.3�V�2e)3��2HdS3=B�28��2��
3xU3I}3���2l+�26��2��3Lr�2m�F3ke�2��3\�3Ɗ3�`�2ҧl2} 3D{39��2��2��25{3���2�33��2K3-
�2ۢ3��3��3�{�2Cj�2���2�d<3�b73�s2b��2�c3�[I3��3�܄2۷=3R .3�f�2�:�2_��2�!37�x2Zʌ3SS�2||�2��s3��$3�O53��*3��:3��3��3/�2�E�2���2�I3�$�3��H3�<3!¢2�%�2Q<3g�3�S=3��[2��U3fC�2�T&3�h3K@�2�c�2���3��2��3_*�2O}�2�s�2&�2��3�2�25�)36�3�83��3fX2	3ǐ�2D��2��/3n�Y2N�83���2�X3�	3�l3ڥ�2��3�2���2�3ɵ3���2�K3�0-3���2pX%3;|`3���2�5 3ސ2�*3y%�2 Ǘ2�39�2
j�2���223���2��2�}�2�\�3-3�3]9X3�� 3N5�2���2�2vig2�s37�3��73^Xb39��2 J�2
y/3��2�c�2��2>�63���2�N3�S�20y2�Ś2T�3)�2��2���2!t3�I�2�	�2�u3�=�2�,3��03���3��	3���2^{
3Z3�x�2m�2d9�2ߛ�2|��2��?3{�3RF�3�y�3�4]��3�M�3cb�3x}�3��P3���3Q��3W��3�s�3��&4�x�3���3��M3�c<4�Y4�b)3��w3�3o�3?qS3�=t4Sx�30s�3)3��4��3T��3/e�3R3�Z�3�v�3a��3��o3�!�3:�4{4�4��73��3�o3�>c3U�3Н�3<kk3׭a3�U�3 �3xw�3��3�&b4z):3NZ�3�f�3�9�3*�3y߆3M�3�3D�3V4ա�3��3Thn3Fn�3Z�4�73PZk3-G]3�ő3P �3:��3ɲ�3lV�3��3j4�J�3���3�ԛ3r�3#!Y3�Y�3���3"n3�G�3Q241��3�"�3��^3��3<��3a�3���3�)Z3�C�3y�e3i��3�l�3�F3&�83��%4D��3��3�'�3���3�z3`��3%:�3q=3�h3��3�4kr�3�e�3�j�3Ϲ�3g@�3L��3��U3>�54O�r3�4��3i��3�0�3�=4,��3[i~3B��3t��3S�3
��3�ĳ3�m3�3�a.4��3���3ؗ�3��3͗�3���3�#�3��3��S3Z�53�G�3��3H+�3��p3��>4� �3N�3��3��*3GZ}3wƑ3f�4?$�3Ӧ4��4�-4{��3Ùd3��3��3��3}��3���3�3��3�V�3Iֱ3I�3:��3oL{4~\p3Z��35x�3.>G3q=3)��34��3�{#3��3��?4���3T��3u3� �3F��3�;3��3J�h3�£3P�[3�$(4LV�3�J3��3�
4~֝3]��3R�3�8�3={�3i��3-�3�H�3qd�3p��3���3�]�3,^3"N4���3��3��3VӮ3HH3X�3�	�3�B�3���3�a93�4�}3w�3rf{3j.�3Y�3�ot3|I4;S:3��3�w)4?0�35ԇ3$No32�3��3[v3){�3�)73�J�3��30�3��34��3�3���3�g3�(p3��N3�6^3G��2~�p3�>�3GR3�UD3�P�33�3 GR30n=3H)�3U_�3I.3��,3�S?3j��3��534��3g��3jv�3�6�3u�3��03��L3�3N30�03ԦH3��Y3#ރ3�ce3ZTY32�3[�3�L}3���2B��3���33�33�EI3��2�3kg3n(�3[	�3�3���3�o�3�{73	�T3��3TѨ3p+3�؅3y�3�|E3"Ao34�4(�3��23�,3j��3��\34�3xQ.3lM3>W3��3���3�Z3�Y�3�Bk3)�3Fe3���3IJa3�>3�{�3���3?��3*3�l3�6�3�i�3s�"3�3撅3���3���3�i�35�3��3]C33x҉3vU3c3*�3	$4!�3�B,3�_]3�@�2�@3-E[3�T�3��<3AU�3�7�3;�4�3�38�3\٫3��>3�o�3j�	3��j3�8%3���3#�3��93��E3�1�3)3UG�3��o313�=I3m�3 �3�d 32��3���36O�3r��3�eP3m|53J�3���3f��3ֺ3��3+_�2X^3�X�3�&�3��3='"4��$38n~3�yP3B�23-3?3���3n;�3��3ڋ23Ⱦ3Mӈ3V�3z\�3Y��3>�e3�T�3��3&�13#I�3�_23s��3N3�L�3e�3S�3%k3� q3��r3i��3��$3>L�3�.�3��"3[�m3T��3ĳ}3!&�3��03"��3cG�3�673b�3���2��3�`,3{��3-Q$3Z��3��P3�w�3��}3d�f3���3{��3r.f3`PZ3��g3�93�M�3��3��3�s�3�Y�3�e�3^T3�@3��3kH83cl^3st�2i~�3j53^V�2V�3�:45�_3훆3ι�3o�?3���3t�3s=93[�	3��b3`Ֆ3U��3�Y�3�!3��3}��3
\C3���3�=�2A�3o�3�Q�3�T3���3-�3�H�3��3q��3��3�4�s3��N3���3"�3 �&3��#4H��3���3�Á3!��3%�3�n=3�s3���3�3�I%3&��3��3z��3��d3���3�;73ž�3��3P1�3��3[�3�LO3�Fk3��3|Ը3O
4_��3$�2��3=�3��,3��3g��2,��3;<�39��3[��3��y3/��3#�4r3y�S3��J3�3٢�3��]3��3՟�2%��3�s�3dޑ3�g3O�3�B3�`�3�y30ũ3�[�3���3��O3N�s3S3���3/^63h)�3�h�3f�3*UG3_�>3��`3sop3<6�3G�03"{�3*d4���3��|3+�23Q�73gif3"_�2*8L3*h3���3zP�3�G�3L*M3t�g3K�C3��!4�3�3Z%i3Gs_3|K(3UO�3��3��3��63��3>$	4�$�3(�-3��$3��3�p�3�b3(4!S3�Mk3G3���3qm_38��3�}�3���3��23��w3�F�3�_�3�3��v3��m3���3��3n�4�{4w�k3��3Ź3!��3��3���3XR3Ĳ3h�B3|��3�b�3y�=3��:3�^4��3:,�3�VW3���3�C3��W3�Ѯ39�&3Ā�3X\�3���3t�d3�(3�v�3� Z3�e:3`4�3Y�A3\l�3�Ç3�c�33�3���3�.�2ri�3|�+3�hi38/_3���3�-3�d�3�+�3�� 3 �3n��3���3�,,3��x3�N�3�8B3/�3�O4>��2tV�3�%�3>a�3�\3��35)13�D>4RWK33�+4��t3�v/3��3��^33�2���3�<�3���3���3hj�3`z�2���3;��3]za3�< 3��3�j43Y�$3��3�.3���2�44��13�>f3�7+3��3F}v3c"_30�34:�3��j3m{g3$S�3�N�3>�3�"�3C�]3IA"3f�y3YX3��N3�Nw3���3%��3 J3	3��o3}��2��Z3#�3��3�Z3eP33/�&3Kj�2�!�2P��3�13n�2�z�2N|K3~`3Η�2�?�2�r3vt3i) 3z�53��B3�E3��B3#�y3჏2�њ2>��2�3U��2~y#3�;+3��2:S3yb3�Bg3'��2bZ�24�*3&3�3�8�2��2�?3��3v�Q3�2�G3���2�C�3�U3ݏ3�<3W3��3R%�2h�3p�3.33�Zq35�43��2	�2�q+3��3�]�2h�!3r��2Y�#3�#�2E*?3}�3��83SH�2���3q��21�73�3Z^�2�(�2�G3�2+3u43#��2}�3�&33rN3�Pu2�3��3���2�A�2]n	3t8W3���2Ȧk3v�3e�#3�2�Ǔ3��S3Ez�2��23��3�43�qP3k�
3�k�2�3�q[3uk3��3Y��2�/P3�W3�	3��'3��2�VI3ܿB3բ�2�#�2���2C�3�3���2��3�3�C�3h,'3�d3H��2v32��2w%%3<bb3�@�2�+�2:K63�J�2r23��34y�2Ԭ3��3Q'3ϟ�2S�3ߥ�2���3,6�2��&3��2B�3
X�2�{�2 3 �2}�3�ߊ3�U3	�34p3��2Y��2��2�OL3iuK2�Y:33�2RO]3���2���2���2T�3p7�2N�3�3	��2�"�2#P�2b�3�݈2��>3�	3;�30S)3@O�2�qV3���2.��2�o33�y�2�AJ3�Ƿ2E�N3�ߦ2S��3Ķ"3�[�3�3虴2x��2�!�2��2��'3�c3���2}M3�q�3�e�2 (�2Z� 3�t3��3���2y��2���2#g$3�;�2O�3,
�2+C�2�2F�3��2=� 3��3��93���2��=3��3���2"k�2��G3o�U3Ȗ93��M2S�13��3 C�2׼�3���2�c3��2bR3�Ͽ2X�M3=$3��3 ��2Ü030,3��3�v3�zf3��;3�b35�3��4i�p35�u3e�3�G�3.�@3�?�2<3G�33�/�3��3��z3l�3i�3�[3X$�3�S3.|@3M�i3��3^�3.�3��3�
3��}3-��3Z�3�o�3^]�2��3R3���2.�P3�C@381w3�p3��R3S��3��<3��U3W��3��63s�3Λ&3%��3H"P3���3H�3K}353>��3e�a3LBz3Jn�2���3���3~$3�OC3��2�ˑ3?��2(C�3��Z3�T�3ol3�3	3�܃3�	M3s�93�H3H�v3ܮ�3�x�2�s37�3��3��_3Ӓ�2%��3�~3�:+3bn�3Z#3q��3q�h3�)�3hR3L��2Nk3��4�tO3�Y3��m3�L�2��$3e�03��3|�03��J3u�3�Ѓ3�v13p3A�p3�P�2��2��E3OL3�qv3/\ 3��3G��3k�Z3�E3��4;`F3S��3�3���3��2~�E3���3�F3Qpz3ȘP3�Q3 �:3	3�2�7�3�8�3�~3��o3^13�`3ͺf3T��3yQ3^
F3�MO3N�4N�43�ۗ3 �B3U�3JB�3*�3�3]�3��w3!��3df�3�-u3�%�2&!`3`3q3ԅj3t�3���3p3�0[3��53e�\3��3r��3��63ܽ93�P�3�:3�,03mm/3Ȕ3x��2�Ol3S�h3���3��.3�
3�j3]ǋ3���2h0�3a��2�vY3��33�3��3�r3U��3��3�?�3�/�3�Ae33)��3�vU3�f�2\ 63�83%��3O��3^Nb3��3�p3D6�3�zG3�q�3���2��m3�n/3��3s�:3��#3�31��3�K3�)3�Dw3�j13u�3O�b3��3S_:3���3���3W�3l�<3��	3��I3Y�N3�/3q�(3��3a+=3o�N3���3vð3/y�3���3�� 4��3M��3�eh3�[�3��43Y.�3?e3;�37g�3N\4���3�M�3�J�3�'�3���3��3�׍3���3���3��E3 n�3/�3꽰3ą3���3k�3�L�3���3o��30|Y3Gn�3}
�3�p3���31�4��4�ߑ3ֻ;3�\�3[+�3�rj3آ�3P� 3��4Y243k4qg�3�æ3̵43�!'4��3M�3d'	3F��3���2�p�3~2{3~�3���3ED"4:��3[�M3-�]3̞�3���3T��3�ʜ3��3�-�3��3��4�:S39��31�;3���3J�C35��3�B�3�[�3fNw3��3�3#l3�f�3�4�?�34�i3b�W3�V�3��3��3`%�3�N3	k3��y3M�3��3lQg3u3d`4沔3��y3�,_3�,�3���3��3*��3w`�3*�3�4��3���3��Q3�t�3�w�3Ul�3�3\�3k<�3�,�3Wb�3�a�3Ǚ3��3��3S��3���3��3߄�3L�3l�4�]|3:�K3-��3>	�3'�3��H3��3YЬ3�d�39��3�}a3�n3yY4�"3���3���3�X_3�1f3g4��Z3�5t3��$3���3�Ճ3�3��3{��3��3�C�32��3��y3�r3kV�3�׏3?�/3��4�vP3���3�H>3]Q�3k4�3�Б3���37Y4>�3!�q3ϸ?3P0�3=�3���3�j 4�&3fU�3���3�G�3���3@�P3�k�3u6D3��e3��3S�b3�5�3���3��3� �3�P3p�K3��{4��d3Y��3u��3��3I1�35]C3#��3C-3�j�3$p4Z��3��3!�O3hc�3���3/�_3�ڎ3�{3q��3��%3�$�3q�3u*3mC�3��4���2�o�3�Ñ3)�3ȲN3hw�3�.c3Xz3��3x��3���3 A�33�3���3��3� �3�B3w��3Bc3���3�+�3�Fq3�Y�2mq�3�[}3��'3V�3�p 3�J3N^3z�93��2�� 3���3]�f3՛�3���2�`3/�$3-
3���2�� 3;ZA3f{�2Ț�3ni�3g�3�(3R��3)�#3�m_3�.3�6�3�9036�l3��`3�!�2] j3�I�3W3��.3�L�2��E3PR3f/3n=O3K;�2$�<3�!�2���3��3X�Z3��3��4X#�2�� 3�\�2L��2K�3�	39�Z3*E�2}�}3��z3j*a3;�2���2>c3JV3r��2�83բ3"��3��2GV3-/3js3b��2���3�C3)v�2�w:3Q�F3�!3���3\5s3'c3��<3��3 IT3q3M�2�M3cO�3���2$r�3��2xY3��3�+�3��A3X�3j�w3F�K3w33��23��(3 �g3��,3^�V31E3[P�2w3�!�3r�_3�m�2��23��{3^3*3vd�3�Q3`�3��3{&�3��2�z+3e 3V�3��93��S3H|3鶅3ǧ3�B�3��o3�3�`?3���3��3�{3��3Q��30f3\9
3�F^3_TA3��3��Q3N�F3�](3�P(3��3���3-Q3�"3��e3�=f3;(3�]3K,.33�53�e3́�3�A3Ԗ-3J��2
�3$3�a�2F�3�R�2��3J�E3�xo3�"J3EK13��3ӿ3��3��3��2}�3�� 3Sr-3�;W3� �2�d13L��3��g3w�2��3"L3�wr3a�3��k3u�#3�v|32�22�3���2X�I3^�D3�3��3V{
3ʫ13Dw�2�&3��?37z|3MU�2�vO3K8�3�x�3DT3�e�2q�3�t3�3�3r�3s��33���3p�P3�W�2;н2(�3&W3Vx3��>3�B3E˺2��3��3E�2���3͐g39��3u�N3
�2��\3���3�3��3~& 3!�"3��73��3L�l3@|3ܕ:3��3ܐ3f�c3ʻx3�ɩ3��(3 �3�w>3Ŏ3�h3P�j3ht�3�p�3��3}�3��3[�j3wT�3��3ŗh3t�R3�@�3T�i3��38 4�w4֋3b��3���3���3��~3A�4i��3�Z�3w�b3�Ӗ3�`4���3J�28�3e��3�l{3��Q3�q�3l��3�J�3��3���3lW@3/�W3�!4稪3*�3��3\�23��|3��r3%�l3�8�3�Ѵ3E�4��34ńd3��2��p3Ά�31�M3ͣ3��-3�9�3+��3�z4۟�3�=�3d�3��3��3䞍3�0a3K�z3z=Y3�B�3�w�33�I3�F�3M�4P�|3U�3�3z�3�x�31X3?�3��2�i3 /�3���32��3���3��P3si4�P3ԛd3�~�3+��3�4�3��3\u4�}3��3�$g4��3&�3�c\3By�3"%�3@��3�Sq3�3H3�o&3�)M3���3�w3C�H3_�X3.�4(�U3C�3bZZ3Vv3��E3e��3~�63ld�2.b�3H��3���3�?�3]3w�}3���3�BO3C|3&�:3Ʀ3��F3�L�3��*3�*~3�X3�`4#\�3yҭ3�uL3g��3�b=3M!�3y^�3�Bm3)�L3�Y4���3�pc3t ?3	��3�d3�ܧ3�3�Vw3ᵠ36y3�$\3�3�r�3H8o3��L4��03��p3��3z8<3�l3��32b�3!53�y?3�b4�6�3}'�3S�u3?1�3�Q,3��3��3`�3^e�3��?3P'4�>x3J�3�nE3ln4Is3�j�3$�3y��3~/�3hM�3y9�3��r3&{03��4���3�7�3J]T3㟫3��R3}��3���3�g63��3�S�31پ3�͍3�D3��3~�4kw3��3�ߓ3�ȍ3TRg3�|>3?-�3��z3)m�3�3x -4��3D73ȳ�3�nx3��k3E?�3^--3�K�3�D3�K�3��3H4N��3	�44nY3 �C3�׏36�4?t3��3KL�3��t3�A�3�K46��3��T3O
V3ϴ�3,�3�U3�y3�F�3��3M;"3�3y �3AΈ32Y�31*4n6|3���3�}�3�2�3��3�Kc3��3��h3 �3x/4$O�3�s�3(*&3J��3���3�3B�3w:3(�3�˜3o�	4ɕ3��3c�83R��3k@�3���3�t�3d�Y3��33us�3a��3V�3媞3SS'4�"�3�KU30�p3��3�ɗ3N .3O �36��3쏒3��V3n��3�ښ3�3ݹ3�x	4730 �3��w3N�3��3P4`��3��K3Z6�3.A�3���3��3c�3Պ�3���3���3$C�3��z3��3C��3���3�3�ؤ3�x3�ʺ3`��3]�]3�H13�f3p��3꘰3�3	��3;:�304A�3��3�13���3m��3>{3���3�i�3*��3��32��3Ec*3��3  W3Q 4��3�#�3�o�3��3m�O3�o�3�%�3�\3�)�3g;4��3�#�3�J3 S4aú3Rc3�l�3�3E?4�U�3	�3��3^:�3�3b3{�4�e`3���3�Ȓ3��3��3��E3�j�33S�38<�3�S@4�J�3�3�~�3��4pQm3@�E3`��3Z/m3���3-��3K'.4�x�3c�M3-� 3���3�}�3,`s3B�`3NA�3\�h3�9�3P��3<��2L֓3���3���3�qA3��3�5�3)ʐ3��73T��3�s3F�Z3�l�3Y4w�3��3�ʤ3���3���3l�~3&x�3lm93kɋ3��x3�$�3�H�3�N�3M�4	��3�ʑ3��@3�3���3b|�3r�3��3��3��3b|�3$?�3~@w3�jE3��4J^3T�3ئ�3Иe3F�3���3|��3A�3}|�3;|�3�m�3�S�3씕3�ՠ3�N3�g3e9�333��3�J3�h�3���3+�3��3� �3�p�3���3���3g��3L��3Q�3��3�jz3���3�{4���3Ʈ=4��3�j�3�#�36�63�F�3�$�3���32L3��4Ռ�3_?�3{�l3x4&4t�3��w3��3�e�3��I3�2�3���3:q�3�{	4��38h�3b�4�3���3�u�3[�n3'��3��^3F��3&�o3Z0&40��3�6�3��P3���3y0�3@��3�K�3���3n8�3�3>ݹ3�{�3}��3�W�3Z�84�3�D`3���3�A�3��038%�3�}83��3J(�3�s�33�3Og�3�]3��A4�Ξ3���3_s�3��3Ͳ�3��3��3��!3��4��@4�%4���3P�/38,�3���3��3�r�3�3�8�3�Ê3F�4���3��3���3�8$4��3-�3�-�3��3�3�2�3c�37�`3�8�3�R�3F��3!��3�3- |3�ב3�Ų3R��3�Pj3���3:�U3�M�341s3���3{�3���4���3:`�3m�3�;�3'!�3@	�3J,�3dX*3ޡ�3Q�4�^4PE 4��3o�3��3�-l3�9�3~�3$�3�C3x�3;d�3�ŝ3�T�3F4�7�3���3*��3 ��3���3�1�3�h�3���3�b�3���3*��3M3Fy}3�f�3N��3	�3�I�3HƉ3|e�34o�3W[&4 ��3��3b��3.b4�Eq3ͱ�32۷3���3>(�3���3Q.�3�Er3���3��4�Q4�l�3?�@3�d�3}��3�Ê3�V	43��3�e3p�3�j�3`KS3�	�3���4\!h3��3��3�ْ3�݌3��3ɕ�3�`�3�M49�3}�4�Y�3�_�3��3���3l�:3�u�38�3'�31��3�`4b��3'Q�3J�g3$wI4�!�3��4��4�3���3��30��3�"3	��3I��3Z4��3B��3�8�3�b�3�d�3JB�3#x:3��^4�_�3$��3���3�!�37�N3ǩz3���35K3��)3Ǣb3�B3�[3⿜3qrs3�s23��3���3M^�3wQ.3���3��3Ic;3-�L3Yy3w�I3`3��3&}3��s3z?�3AG�3i��3O�r3U�3�Κ3VK3^3�A�3���3��3���3�ʊ3cS!3T6$3���3�^�3���3�3�3��k3B^3,3�%�3�OL3�&�3t�^3�ݞ3��03�[�3<�3�;13=x.3��l3�~/3�u3雪3*�3��3�b3���2`3'N3��23�F�3;5P3��3	=/3ݹ�3�vJ3o�+3Lo3<|�3Rw3���35k�3���3c$30e�3��3�.,3�ج35��3���3\1�3;/3B+�3���33O3�h\3�9�3`ѭ3�C�3�Ň3	�C3��3�Bl3���3�LY3�0D3OO 3��V3ʢR3*�3p8�3P�/3�P�3��3om�36I�3�3ח�3Ck�3�N3�e�3E@3U��3�,d3�f�3;1j3ȭ�3~#�3lC�3��3�3f�p3oQ�3�38�I3��3��3���3cR�3+��3vo3�43j��3`3"kS3�2m3��@3e�3�03�J�3�?�3Vw/3B�2��3���3N΁3]�U3��c3�m53l�V3�L3��@3"~3M�3��3��g3�	�24�3-ǡ3��+3WP�3Y-3��d3  33�>�3H�x3-t4�8�3H44�\l3M�4Oڜ3*\@3�G3Nd�3n[�3vt�3o�g3KM�3��3%=k4l:3��o3�t�3�{X3�=�3��3.T�3so23^|�3��3U:3�:3�%�4]��33�_�3��2�*03��A3hYs3�E3|i�3Ag�3���3���3=�!3��d3�$�3�d�3R�q3x�3jԤ3#03�q�3��3�!�2�ǫ2L��3m�3F'3�f3�k�3�%3�@w3�2l3�ZM3eV3���3���3��O3�>�2�5�3^c�3�a�2Eo3�r�2�#n3�3fq�3�#3�� 4}��3���3�Ya3�[�3�L~3k�3��<39�3yV4��}3��3n��3�J�3���3��3�ܛ32`]3��\3m��3t��3Q�3vnG3�e�3W��34^�3#-�3h�74-3��3�1s3J[�3]�U3�ֳ3�X�3�U3��v3��-4���3��;3m
3|\�3��13�F31��3FX3k�3GE�3�l�3�ʅ30�3�"p3^s4[�\3i��3���3�I�3l�93՝�3� 4@X3�.�3�{
4���3�Ɖ3|�x3�,X36�3��3e�3ŏs3�2�3C,�3K�3Gl3��3z�V3W�41�o3`ܓ3�ݠ3뻔3�L[3Wd4d�3��3��{3�iY4���3`36at3�9f3��3Gb�2�c�3�!
3��4�T830�D42�83��3Ns3��#4p�g3��3�3N2�3]�3��o3��3q�d3q��3���3G�3 Є3�W439&�3���3�
�3
��3-��3��3C.3K �3B݌3�	K3�Y3�4Jט3���3���3T�3��W3��3j�>3+\[3�W3��3.�u3��3��3�4�4��3��O3�;�3E�3�D�3S�3?k]3G�3��3r+4��X3c�?3���3X��3���3���3c^�3�f�3�O�3V4���3�7�3�m�3�'4���3=��3y$4��3�1�3鵱3�A�3�o�3��F3%v�33N4�l3�Ÿ3i�v3-އ32�y3E�4͞�3���3���3��.4�$�3vۊ3i63��34�l31O3T'�3��3���3UN_3�4uaZ3C*�3���3M�#4���3�ޫ3��3��3�(�3#��3�_�3��83U��3��3���3�R�3%�@3�3�N�3��3���3ڽ�3\a 4d��3-}�3�ݨ3���3Y�3��?4�gP3m��3p��3��K3>G?3ʽ�3�;�3~�k35�3�d4��3{�4��o3$��3�ê3�ę3��3u�$3��4\f�33{�30�3��3���3B��33}3��3���3�03O�l3�lo3��|3W�3W�3靰3�k_3�t3�r�3�3�]3z�%3�ț3�x3y�39��3v
�3���3@�M3�3�32�\3���3Rv3B��3iM53g�t3Ԃ�3��3��3R74l��3�X�3x��2�I�3��3�j3��3 !�3��3��m3�˾3��3���3�d39��3�B�3.E3z�3��P3NxF31K3~��3nd3=�p3�4ӯ�3=�u3�$�2�8�3{�3�r'3S��3j�3}7�3�[D3���3�ډ3Lƍ3�3z�_49 v3U�3�k31R�3�4l3M�13���3�n�3,C�3��3=j�3�r_3�.�2�~}3`�3��O3��3B�^3�3�PM3`8�3�M3�d!3D�3��b4��3n�3Z\�3&r�30]A3V�a3*�d3E.$3��3��3oz�3�L�3N�2��3nN:3_4%30��3T�>3j�3��33lU�3�I<3TԪ37�73z��3���3�|3[^�3r��3eS3"9�3�g�3��2�%F3��3�;�3䊏3�.�3I��3�ɂ3^ �3���3�ZH3^��3`�p3�҃3�]V3�w3��3���3��p3ϯ�3Cl>3<oE3��S3﷮3�3�3�3�'{3�׹3���3TE�3i3��4�et33)3Q�a3n�b3>{�3C;E3��3u*3w`3F0�3��4 3���3Bh3�I{3Lx3K�e3�q�3DW�3�>�37�4��3IX3ŀ23�a�3�3��3Ϊ�3�5+3�93�ŉ3���3E��3�T�3sx#3��B4�ڀ3]b�38��3Zד3��3�	3}�3��N3�ő3�04b�3� l3&:K3�l3+^�3�_3��3�a3Cx�3�T]3�K�3~,a3͎h3G�P3%�B4���3g��3�g}3h�3M�C3 U�3�|3j	3��3r��3��3���3�y�2�9�3-j_3�973�G[3�; 3�"�3�h34�*4H�n3^V�3�pX3ө�3��3�i�3��83�ɜ3�lK3sԖ3��3��3�R3V��3A-�3%p�37
3�}3��j3PG3�r#3W�3��3b��2�[3�:3v:�3Ԝ�3��3H�J3���3�-a3)x}35E384e3�ځ3CVD3���3���3%��3�p:3GG3b�13�QP3�HU3X��3�&3�]�3�3֚�3�c�3M�3Ȍ 3���3%Q3��3S#�3�)�34�53�
3��J3�G34n`3Hk4�\�3�Hf3�o*3,�v3�&�3��2)fq3?L3aBz3J�H3�e3<��3��3G�25�4�,3k�3��3�0L3|f!3'HH3^�3��.3,�30��33ǡ�3	�3w��3��3TJ3��M3xnK3G��3N3���3��3�cE3(��3�n�3��833��3�,E3�!H3�Ԥ3W�>3|��2xC3]U4Q3�3G��3 p]3UŔ3}&3��.3��3�� 3�&13zk3m��3�,3�13k�3}8�3v�3ZD3~�i3��&3��3Ů�3K'�3 �2ǜw3Gw�3BU�3��Y3Q�)3^��3m�3u��2�K93�A^3�<�3�\�2,��3T9r3�u!3��3m�3�3ϭS3��3!+�3�>3ԅh3o�I3+eh3e��3�/�3�3
Fl3�L�2�ȃ3Pl�3���2n�T3j��2��3�A3�ܟ3�t73]za3t�53o9�3�S3�,3a83�Bc3n�3�@3o�G3ʍ73b�M3�U�3�A\3	mQ3B��2l#�3�
�3��W3N^�3#�:3��3�a3Ndz3��b3��=3;O/34@Y13��C3��U3�O3�13~r=3��73]_�2@܌3�!�3f�3�=3KN53�1431Ӄ3�3!3��33�� 3�u�3�{3�'�3�Gw3u\ 3v�3�\-4S3&
`3�
P3��#3dh3*L�2�l-3w��2�H3p�3']36P63|�3v�a3&y3�O30�K3�|�2�h3U3ꈡ3��V3�Ǹ3{3E�4��3���2��3-^�3�7B3�3 BM3��E33k�3(sm35�F3{�3�F3oD:3�P�2	�3%��3?3ʪ�2���3�>3,K$3{_t3�2u3�|83Tj�2��A3i!D3��U3G�v3,�3�'�2��J3R��3@�,3;�A3�� 3X!e3�23�q�2QW3��T3�k�2��J3��30Fo3��o3*�3y��3?�3��D3�D�2���3кm2Dm3�I�3�i3g
3��4�#v3��3��2F�3��G3���2v��3�(?3�B3���2��?3�53� 3�WD36�3�T3b;3�M3x3��3-,@3��/3`�2�,3Yݥ3R�3z�37I�2�-�3�;;3�>43�P35i3���3{�'33U�3�\3� 3��T3�M�3Xq�3��3$�(3��3��E3�T3�&�3v53"�3�5�3!<�3˯a3e��2�L�3J3�3�C3�53Ω�2c3�p}3[l3;�D3]t�2ળ3�3+�E3}��3�03s3*�p3�N43,�2#-43��3�n3ƻv3u�2��{3�)y3903Z[=3��>3d3���2z��3��3�WD3A(M3)4��+3��3��.3cPK3� 3�׈3�/�3��3Sc3_z�3�kp32�3LJ�2�S�3�qa3��2�G3;�2y�<39�3fnX3ٮ+3� W3��k3�Ǣ3H63l+43і13�n(3?C3a$�3d�b3��3{*�2&�3!�3&]Q3�73��3�;3���2G�3'#3�3��3|`�3��'3�x3OQ�2���3J1h3��%3�G3u�3�3<3ԝ�2A<3�733K�3]4�š3�m3�3Ʋ�3�kR3��<3_�!3�Ϻ2�#3L�2FQ�31�33�!,3Uԓ2���3�QJ3�ڛ3<��3�B�3�R23��,3�a3�3�Ȕ3{a3'ǘ3�˝3���2-�u3
�63�*23�=�3b'�2n�3�w 3��3�|�2 �3PP�3M�3���3�U3�
�2�t3���2C^�3�3Y!3D�T3�}�3�n3zP3G=3��3�R3x�03i��3��#3�F3��3�/�37&3j3gb(3�xn3^�q3�63^3�33{)3��432:3�j�2�p03�O�3\|�3;�%3�±2:4�3?c3M�3��"3"�F39Y*3{�3���3�t"30�B3U�r3��3��'3OcK3�N`3[Ɗ3���2QM?3�.O3��83g�3�l�3�K3JjW3�G�2��v3)�3`E3��C3�"3�S3�3��3�043I}�3ñ�2Y�3P�2�k3�Ȗ3`W3�3H*q3�G�3���24�b3���3Kf�3UV
3磻2BB�3��:3p*03�,�3�22��3y�E3���37�3���2�N3��@4s�	3F�93�Q�3��3qtD3k�3�b3l�[3�3��3���3��3n<3���3(L3��g3W�o3Gt3eG3�83�%�3�A&3�Q�3u|3e�4k��3̰�3��<3 pj3��f3t݃3�83h��2�w83J �33���3��H3� 3d�3��3	%�3()3s��3%�U3�o�34�3��3w�2�j�3�R�3��;3��38�2Uܕ3�q)3�z�3�O�3�*�3~'�3=͞3�Gf3�f3'�3��c3��3<��3�F3!�c3��[3-�g3u�m3�%l3���2k��3�G3s<=3C�n3��,3�t�2ۄ�3;L�3�.833��3y��30D�3�[�3�T3zV�3��3�#3��3�k3� �3�<3uq�3�
E3�y
3�3G��38�3��3-�3��y34�S3S�3fe�3/3xuY3�r�3ˍ�3�K+3>b3�453�I�3��r3X��3��%3��|3��C3N��3���3��3��<34"&4lG(3k��3��x3@ˠ3#�83�ƙ3��P33mO3�ٜ3}�3��93A�3[u�2�3��V3^Z�2A�3���2�Mw3t�I3K%�3.3b�3N�#31,3.ݵ2u>�2�^�2��3Mv�2W�Z3��73&s3��2cd]3�3���2hV�2TpT3��3^G�2�O3��2��;3�8�2�Z�3���24H#3��>3oZ3Ev�2�` 3F�3Ab�2C�3$��2�3��2��3��$33�73(�2$23Q�20�3�k)3Q��2�3��3�s23�3.�$3S��2�3���2pA�2c��3w�03"Ӱ2�g�2c3��2D`3��3��"3
L�2%e�22J32F3���2�3`ҋ2��3��2�Z3���2�93��2�J�3�i�2��2(~�2a��2�u�2@�2�N3���2`3;��3T�k3 ��2Td�2�G3�8/3}�2�3c@�2���2�b�2�d3���2�`�2.82�p3�%�2/�"3�3k��2��3 �35I3f�2�+�2	L3�w33t��2�hx2��)3E�3�Ԝ2�933^�2ǇH3eS�2�R�21��2yc�2}U�2��D3++�2)�28n83��3)r3p8�2���2NS�2B�3�b43��2g��2r��2p�3}��2a��2��E3f�2�K=3Z�2�43T��2��24�2�ɧ3���2���2k�33��2@�3�3d\�2���2-�2#�3��83�3	3#�2�n3<@3��2u��2��2nQ3��2��3Pw�29�2_�3�3���2ZZ�2݁3��39"�2tr�2(.3ጻ2���2A�3��S3�~3ˎX2�@Q35� 3Ĭ�2/3�l�2�73˝�2wb3�3���2�X�2pz�3��2�3i�3�:	3Ll276�2̌�2�U�2��2�#i3�Kl3"�=3)��2!\3D3*3��2���2	_3�)3�F�2��03m�3�V�2��2�ӊ3�گ21��2��2U$�2ך�2�3�	3�ڎ203d�+3[�3ռA3�|C2��I3+3�a�2z��2��2�/�3$��2_�2ݦ%3��3�63!�/4Ǹu3~3�3�"�3q�#3j��3�%�3�5�3�U�3�l�3���3��q3,35l�3��{3k`z3�3�т3�3'k�3��4�6�3
�M3p`3ί
4D�r3.��3�u3W��3�"&3t֛3EMP3I
�3�9x3���3iU�3���3��3:��3��d3?#�3y�X3�#3R6�3��d3kn�3Ƥ�3}�39�D3'��3�%3��3�4�3|M�3"!�2�׆3S�3�!O3� <3�ѫ35�j3R3W�v34�3���3�_53{�3�.3�9�3Y��3J#w31�3_Ő3^&�3��4A�B3�T3�U3,[3�{K3��32�373���3���3�:�3��S3+ X3�Y�3KJ?3�53�-�3�?�3i�3�&z3԰�3?d�3jN3c-3��4�X�3^��3~ұ3��,3�Fw3QH�3S��3��3�T�3J�3�J�3�v�3���2m{�3;X�3�43x`�3~Cd3�|3�b83A�h3���3|ރ3r�53_E4%ED3���3%��3�"�3��63���3�`�3҉3���3�1�3G6�3�I3�Ԇ3Y4�/~3��T3�p3<cR3?J�3j#S3�O�3�9i3Oh�3�N13p��3�R�3H��3yV~3R�`3B�3w�3IC�3��3�S3�	�3�8�3$-3Sn�3~��3��q3�(g3�3�32_3��36�U3��3�ڛ3�	�3�i�3L�4�L*3��3<�A3�3g3&g3[��33�3�݉3��3�
Y3��3�,n3(�3�r�3�A�34.3�Ӯ3B�3��3�/s3�W4�`3�1�3GZ�3�@849d3ь4�L�3aj;3~.3�M�3���3U�3bU3�F�3�Hp3X(�3�N3�3�$�3a&�3�{3�.�3M��3�3\��3��3V�S3�3�7�3�nA31s3V_O3�g�3�,<3�243�-�3QN3�ڻ3���3�4��3h�O3��3Cګ3��]3��3�ה3U�4S��3n1�3�3�`3�3���3�+m3���34BT3#��2u�F3eu�3��/32AQ3pa3~�R3�X�3)Ro3283Q�3�73�3]x;3�x3�y\3w@3R��3�/3�b�3�3n�3S`^3^� 3\%3N3���21�3
<�3�"3rR�3��3�Ƌ3l	z3���26�3�-3FX3��h3�3$��3�i73�*�3?]�3�3o3A�.3Tv�3Sw3�Y3��31�3��3���3���3��@3X��3.\�3��3Ť�3S��2���3~3�"�2$d^3�%�2��V3�bS3���3��3��L3���3Uٰ3��)32�k3x]�363
��2�D�3,��3W�V35��3���3�3�e}3g�28�3fO�3u�$3	Y#3�� 3X��3��03 P�3��3;3�43uD�3U�(3�ia3�)Q3�6]3�
A3��l3���3�H3ؒv3�n�3*H�3<�]3�/ 3L�K3o��3,_3w�c3�33�53|�23��3�,3ѹS3t�3`�4Up3W��3�y3ު3� 3�׳3mG�3�H+3C@3�#}3��3��3�b�2sđ3O�k3��3j�3�L3;�3� k3T
Q3]Q3f'3��2Ro�3��D3=�,3��q3Dw�3�63RDG3�Y(3Nd;3=�]3��4�Pn3pz3!J�2�K�3��3CqX3{�3V�$3��Z3Cm3�,�3}v-39l3�3E�3���3��3��328u3�.�3W($3���3�ބ3�ԃ3"��3��d3:�a3��33S�N3\�Y3��2iZ3
)3��n3��Q3���3�~[39�:3\�b3W#�3&�3�i39C+3�-3�W�3�3���3=(3m�Z3{	�3�B�3|�^3��)3-�93D��3(f�3���3��3�\�3-�3��B3��p34#�2�B3��n3`�3A��3�H3"�X3��3�3w��3"T3>�3ԛ�3"��3>p�3�|�2{=3�s�3#Io3>uF3`�3�uY3��3`0�3MO3�(3C~3��3X�>3c(u3���3��&3��3 '�3df?3��3ï3��3b<+3|}3��@3��k3u�v3��3M�M3��'3f�i3;3�]3�ii3��?3�$K3<�3��g3�ݢ3dVZ3)�k3�)p3� @3�3��13���3vƊ3G�3�!3���2	�_3�P3��2��p3��z3>�V33�G�3�e3�k3�� 3���3ms3	�*3ח�3��3ws	3�3..53���2�3���3N�h3�-3���2+_f3Xh3���2�Á3j`3o3��3�>3HNJ3�a,3��>3���3ޞP3e�3�wA3�w<3�-3ՄP3�r3�<3`3��I3�k�3Q�z3?��24K�3%/�3L� 3E3��23�nV3]� 3'	X32173�h3���2��d3l��2~�F3�oD3V3}�24�S3 �3�m�2��_3��3"8i3�_C3Ƿ3���3M �2�3c�3G3�)31�3�y�3?3�23�j23��3�3�3��;3X$�3�#3��[3AĀ3x� 3���3�ҩ3��Q31-W3��
3�gb3b)y3��/3Ɵ�37�3ɢv3�3���3Ԏq3[pB3�!3@t�3���2L�3��3� 3+�=3K�m3Q�93�1�2�؃3�T�3Z�<3S�<3(<�2(�=3f>k3G�3:3��3�b�3�O)3Q�{3A&73+�E3\3[��3'�3ȋP3]Z3@�3�m/3E	3tx3kg�2�%73�"�3�T3>*f3"f�2�3�H,3{h�2:��3bD�2U�{3/N3H�n3<�
3���2�k3(&4
3b�3q93B�	3@�3�Z+3�C30��2��13V�u3
3YF3"C�2ƀ�2�x3�N�2�Y�2���2���3�h�253NU3\��2��2A��3���2X`93�3�.�2ܝ2��3|�~3���2��:39�3��`3�*3`�2�Q[3C�!3�s*3��:3�>�2��H3���2��3˘3�1A3�2粒3^�3�3M[�2	K�2�R�2�A3�Bc3�8@3i&3�λ3�$�39AT3��.3�]�3�[b3y�2��3�!3m�B3���2\�z3�f3��83�x3R��3c}�3d��3L3C9,3�}35w�3�9?3ʺ!3A�!3O�3�.�3$c�37��2)v3��F3��3b�m3#�3
��3�#�2葅3�c_3���3H�G3�U�3W��3ƧC3�l@3i�}3�n3:�Y3Xl�3@	,3�mM3q�3r\3�@3�5�2� 3��73LW34?3��33w3���2;%�3G�p3��J3�_53�4`On3�E/3�ʗ3+r�3=-/3%�3�qX3�ζ2v63�3��3g:�2 ��2:Z�3>�h3��2�G3�FV3�3��n3�3�3W13�P31w�3�
D3ݽ�3�`3k�*3�΄3DH|3Żd3S�23��3�-�36�s3:QN3�3�<p3��d3��2��3Z�,3J�-3l�`3-��3$�!3�n33�3�4��3��3<�3G�?3�zi3-}n3 ��30x3�w3�38{n31�s3BJ3C��3��P3p�2LST3-8W3=2�3�[
3z�3�q93cZ
3.��2N"�3�Cj3��h3�e]3g;3��3�oF3��U3�63d�#3���3�3�83��3;B3�X53l�3\|m3X�2a�y35�L3s{G3�vD3]sd33�<3@?�3�?"3T�*3	3z�35J3�A3lm�3�e3��`32�3��3�?3�63��3�2?l3h\j3)�(3v�Q3A�34�3�r�2<��2�*�21W�3��3��3>s3���3�B3b	
3n�_3.9�2��g3R��3a�z3�_�3�l�2Ql3��3��3@j?3��33NOQ3U��2�l3��I3"w�2�_3�Ω3��2�=:3�6W3��F3:��2"�Y3>U[3��2�OK3s3]l�3��3���2��83�{3^33�H�3���2��3 #3Bwh3��#3���3��3���3\P�3+�3w�w353�s3'd�3Gh�3fB3<�3og3"�B32��3EO3D��3�S�3�y3S:p3?ay3 �3Ѝ�2��4E��3� �3R�3��4<�Y3�Y�3�X23�Ւ3ϗq3���3�3�3Xr�3��*4i��32�
4��3��3���3�H3Ɏ�3�VT3�d�3d�Y3!��3A�g3t��3�c�3�	4i�3���3^8�3/�3��3��P3���3��m3K��3���3�4aQm3�3M]�3~Տ3!`3m33�pS3��3AD43!��3�RL3�d3EKm3�+4#�3��3�׆3�E�3��438s�3G'�3m�U3��^3@�3��3\�<3]�3���3��3(x3�"�3|�G3�3��\3!r�3X�J3n0:3,��3%>$4c�3`U_3"3%U�38f93�l�3ڂ�3L�*3��|3��3�r�3�en3�i3��3�X3�,3�[j3�~$3���3��3��3�l�3��~3C�03݋34FW3��_3�z3�}j3S��39>h3Ĭ�3V�
3n�b3[4�O�3`}�3#_G3Nő3;ڡ3m/q3U�U3m�3��3 ��2/G�3re3#d.3��]3Q�04�}3Lj3=[S3�D3 ">3���3u�3߱3cT�3��3�3�6e3CR 3�]3�Cg3|�;3�y�3D23s��3�ӣ3.ب3��3y��3��t3���3�.43j�r3>��3��r3Ǽ?3g
�3��4�93�w3���3D<�3�R�3��-3���3,$O3��3���30s,3h��3(�3���3��v3�V3X93�: 4��3���3Y��3�Ò3�_�3	(X3��x3Tp�2pI�31*�3=��3{*�3mg3~��3�3��}3���3A�2ﰤ3.(3sX�3.��3��3ѥ;3.fO4�/36�t3���3�)p3�)3�(a3��3�w03=��3��3���3L܈3N�3�;�3�8�3�Z3}ԍ3�U3�3RTJ3�"�3:�3���3�h3,�3;��3?{T3팋3�4OYT3���3�D�3�%i3f,}3i`�3.�3!��3���3�#�3\��3|�k3�ם3#H�3%9�3��3���3�#�33�	�3Wa�3n��3g,�3�;v3{Y�3��T3�`�3|�3��V3"��3K��31��3O�p3JX3��~3&O3s�i3V�l3�d3]ģ3{�3g 4�kO3�s3�3R3��]46� 3@=t3(��3��3���2��}3:�3�b3|p�3��4<Y�3n�a3ѿ�3�+h3���3�S3�D3���31��3�g�3=*�3�/3�;3Zt�3��4k�l3oD�3�+�3��c3K�:3F	�3���3PD3ډ�3�֊3r��3 �q3���243|��3��3��q3�>U3��3�	33��3�\�3�r�3׊@3��.4ʩX3�CD3�+�3!h�3�e38zR3�ۯ3�4p3�q|3}��3���3�V3W�2��3|1�3�S�3�P�3V�3���3�	736i�3�83%Zt3;z3� �3})3�3K�$3q53�E3WoN3�x~3��3r�T3q#�3Bc�3-�:3.�*3<�3�%�3�'$3���3��h34�d3I�3L��3b][3(��3��/3���3���3i�(3��G3xa3_n3�׬3$�3���2Wl�3�x�3�ҏ3�L�3�;Q3<t�3�w�3�3b/�3h1�2L�A3�@3r0�3j�Z3���3k�3"��3�rU3��3v��3��/3(��3��3�d3n^3��j3dȝ3-�3���3K83tg~3kf�3%R3+�g35�G3R�A3��#3ӵ�3"[34�Z3줠3���3��$3�z�3D�~3�lu3��M3�#F3Ș3�Y 3�߆3Y�3���3{<�3��I3�3?3ܯq3s3n�35�3Ih�3���3 �r3�;|3�\+32�S3�n4?,3iZ3[�3K�3>�3��E3�{3�I3=ޠ3u�u3`8�3-��3�c;3�[�3߄4��f3�H3Dc�2U�3�_�2���3�dp3�3H3��!4OI3�q.3�ԍ3Ae3SM3�<p3��>3�jz3�(�3i��3IČ3��3��?3�b�3��3f�2�3V�E3O��3X3��3�?p3���3T��3��3��3s�o3�l�3��3�sA3u��3��4 ��3�4�3���3�7�3�(�3=��3�3�1D3�Uu3��3�2%3���3'D3vͽ3�p3��3,2?3��3�c<3��X3��3
�3�
'3�y�3I�3��3�N63��4!�3۽C3*i]30$�3]m3�G3 w�3���3�޶3���3�4�x�3���3���3!�"4�1�3-�^3Ή�3Å3.Tc3t�i3���3��f3p3��3��3��"3��3B"�3��3�713��3��_36@�3��3'<�3/Bi3|�N3g��2(\�31�P3:RJ3 ?�35��32�3�R3ԍ�3j3���3pw�3��3'��3)3f�353ru3�3W.O3EY3: r39I�3j�3N�=3��<3ۧ�3��@3�|�3��+3��3ϊ�3&k3��3��2Tċ3xB4�ΐ3���3���3��3�3Fv3�Y3��	3`g�3��3��n3�3q�}3��93�4e�3��36�3 vL3�3qI^3�3��;3��3�[�3���3.��3Na[3.�3�B32�3�H�3���2�]3vb3?��3�&�3.�3p�r3�|4¯X3�T�3�Q,3�H3��3��3~�3�
k3h)w3O�3��350�3p�/3�	�3਑3{93�q�3��&3���3VW=3�{�3�x3���2��3��4d3%'�3�a3��3yXT3Q��3�v�3�`[3@ņ3sɲ3��335J3�d3&>�3�{�3f�e3���3i39f3O3I_�3��*3��)3c"<39��3��t3�ܪ3��3AGk3Z]�3���3�ܢ3% 3R�3��4
�42��3��2���3C��3��&3���3��63HF�3Ŵk3��3�V�3ᔈ3���3\��3]213ܪ�3���3Ӝ�3	�3��a3��3���3�3�.4�3%'h38�-3�,�3���3v��2�e3wf�3Xt3#6V3���3b[3�>44��3�F4���3��3nW�3R�v3�w3U,�3��3tA�3���3k��3��3`ͯ3pqi3_��3�[�3;t�3`��3Wrp3���3k��3�;4��3�<|3ɾ�3I�3�.3Lf3�ڣ3*ت3 �i3,��3��3�X3���3�
4M�+4E��3B��2�t�3[H�3I�"3���3��r3�[�3�g23^��3�bp3R?�3N4��54kx3��3��3��|3�0�3RF!3�%�3~53��P3�A 4�8�3)�3'LY3���3�?�3���3���3|�3��3�3�3���3�{3~9L3Y�u3���3	JW3;�3�a3 w�3�q�3�@�3� �3��3:��3��4'�4ɨ�3F�3��3���3�P�3�7�3_�37�3!�3�Q4<Լ3�#37)�3
�g44��3�Ʈ3h�3���3a�q3D��3^�i3q6�3���3Յ3d�4$P�3-x�3lL�34�,3�3UP�3��3�r�3�m�3� �3�}3 �3B��4&��3PC�3�+3�p3�h3!��3�Ɯ3�u`3I��3�Wb4��3v�l3��539��3�2k3*F�3���3��V3��3E&K3(Q4p_�3�%3k$�3��-4��,3�0�3H-Z3k%�2F\G3�;3fq�3u�3I��3 _4���3X)�3�6Z3�=�3�;�3�*�3�4�/03B�3�A3~41cD37�Q3`/�3T��3��3���3� �3]_�3J�3�+�3�3>,3#��3��4���3���3���2n;�3�+�3i��3��3�Dd3���3>y3��4��|3�uj3�'3#�&4�2_3�Uu3:�3�m3�Y37}P3��3�D3|h^3c��3���3�E3�'3���3�U3�J3��3��U3��K3��+3���3�63�M�3��R3M4���34�3���3~�3��3-��34o�3���3��^3�,�3%�3��24�,�3$��3��W3�493 g�3j@s3��3L̙3��3�p�3��3c;g3]�3�6/3��3X��3S��3"�s3�3�]�3O��3I�b3f��3��3w�3�^3'�4�K�33��3��3���3p�3�ɋ3�24��3D.�3*�[3M�'4��3�~�3��3B��3`K�3N��3�l�3���3�ֱ3��3}�3�ʾ3@�4)��3���3�D3k�3�z�3j4d�3�4�-�3�X$3��l3��4�`s3��3W�3#��3\+�3��3H��3�r�3�^�3�4eP4��3�sP3��31��3�c\3�ӌ3J,�3ץ�3ۤ3�)	4���3���3@i3\4J��3@$�3x��3�3�-�3��3Fk�3sK3`~u3�4aO47�3�W3f,�3���3�uB3�>4#@3��3��g3
)�3�&<3��3:;\3ت
4eK3B�y3/�3k�l3O��3�Q�3�4�3g3���3���3��3�Pk3t�S3P��3ʶ�3�I53+>�3�~�3��3g�3��3-�r3_��3U�L3bX#4�$53�K�3��3��Y3+��3�S�3�ʠ3�)X3ZH�3�794,��3�-�3CJ3}@�3���3� S3��3��[3�r�3���3���3���3L�3��3�46��3���3��f3�!�3TL�31Z�3v��3��X30�3�s�3�I�3�s�3��V3K� 4!S�3�
N3*��3��s3L �3�~3��3�s�3���3g��38=�3�b�3�3��4>�3��3�p�3 ��38�^3���3K��3��3��3��3�#�3d')4_|q3�ð33h�3�4H�{3���3B*�3!s3���2�G4��]3�3D[3��g3�T|3��y3F��3#73�f�3b�3���3�O�3	mR3�@4)'�3N+U3�Wn3��;3��3�\!3�u(48˶3WY�3#�;38�3�-W3y�>38�?3��13�~)3��g3NC^32�(3�"3�Z�3��a3�n3�-3��y3D�H3�tU3���213��'3=�3yͭ3��H3֑�3�\z3���3		X3ƅ3��53\�M3�GZ3�3�3H63]R3?=3
[�3!ʣ3Jl�3<C�2x�?3IC<3/�j3�I3���2W}F3`�2�^�3�`�2M�3��,3�3�`83Z�2���3V3�Y�24�?3��3jH�2�4O3!,�3�Z-3s�"3䷣2��'3�J3��2�f~3%r�2�cr35�>3;y�3M9R3#8h3���2���3K{3X�03K�3*�#3�z]3�S3i']3��33Hk�3a��3�?�3�_#3-@3T�-3~�T3?�`33B�3~��3��&3�dK3��3A�]3齮2�-4�)3R�Z3�223:�3.�!3z��3��E30��2��A3>3�36Os3�&3�v 3}
+3}&g3G��2Ht�3�4'3&Ş3�/3�ҍ3-{n3�N3��!3��3�Ն3��M3�U,3ҧ"3�2�2�<3�n3w�2�3���3=a83W�E3���2�<Q3=�31s�2g�3�3��l3���2.��3^/3u}�3�o�2��4��`3�UI3�;3��?3�g03p�K3�+�3�&3OY#3��%47�o3IS23�3�/�3?mF3��S3ھX3@v3�iO3v:3 Ҕ3�63j+3M�3�|�3#�3��
3�q3�q3��.3�h3�>)3�O3�$;3}K�3�p�3�o3Б�2�
]3��g3IvK3#��3�2��m3S��2R%3�(P3�?.3J�3lQ�3Iv13��32��3�Fm3�Q03f�3��3�'3}�z3&��3A5�3C��3Z�2D�j3���3�Հ3|�3�4+3��?3Eq 3���3�,3��b3�1*3a��3�
�2;?Z3�T3��P3���2��J3�b3�'�2�M03���3ˁu3�P�3E��2O23\�3¡�2z1*30?3Rs�3���2c̈́33$��3[�X3[j�3�-S3z�G3�S3��13��03~/y3���3�3�et3��3I��3fk=3>
r3�ԉ3���3�ee3��3V3ǅ3�p3�l3,��3p�3}�o3,5�37+�3���3�;#3ѽ(3g�73`��3��c3�;3,OG3CJ�3'�3��C3켾2�~3���3�37I�33�d3��3f}3���3wH43��U3�93��3�!3��n3�D3���3^�n3��+3��3��B3VQ�3��4+خ3S�3EQ#35�i3Aa3D�2ߍy33%3fG3!�=3O�3�@3t|3���3�o�3Y�]3E͒3h;�3���3 _33�3 ]�3�\}3��3ju�3Aҁ3�$73��2b�l3ڥ�3��M3�p�3�9&3���3*!,3��3M�;3�3�:3 ��3*�*3i�2K�T3G53���2�f�3�]�3��3h��3_M4f' 4�>3��3Г�3>�\3�)Z3 �u3�oO3�q�3t�3u!�3�%53>�q3J%�2�E4V�w3�\�3�M�3?'�3�3~3��03)�g3@�3Б�3�N�3J��3/G35(3|�W3J��3�U�2 a3V3�3o?13� M3�=93�B�3��3/z
4K��2���3E�3��3o�d3��3P��3��\3%zO3(��3m�3��)3v�U3�a3�X3	�L3Q=G3?�*3�A3�@L3Zܭ3��3��3�. 3���3B0N3��W3�t3ii�3��63�c3=��3��	3��3)�4य़3k�R3�W�2���3	�3l��2�h�3���2���3�_3���3���3��Q3J�K3��14X	3Z�3O�E3YG3-n�3��|3�33�~*3�d3E&�3#�3�)�3t�2OMn3��Q3�݋3��_3���2ԃ�3_�837�3�3]�3�*3�
"4��Y3��A3ic3�MV3�>3��	3g3�,3�Θ3Mͭ3YD�3/�3�k�24��3R�q3��z3'�3�fs3�S�3|J�2��3�3=�3w43��\3M��2�M�2�D3A�H3�ۤ2��93!+(3�3�3��K3�3޶H3�š27*3{n 3�<�2�3��3�H!3R�2�3;�'3e�&3��*3�+V3��3`��2iQX3�+�2;%3[3y,3ƪ�2u�3MC3�"*3�Փ3��3q�B3���2�2�4�2�H3��2|�?3�c/3��2 73bp�2�Ǥ3��3��I36�2k�93�|�2Ll3>�-3��2��2K�3��3�ȴ2���2�H)3%x�2�ڵ2�3���2��3+��2bS�2KC�2��3��3��v3J_72wF�2��33�?3�2'��2��13\�2S3���3]�B3wJ,3'"�2�5!3��Z3���2��!3�$�2�� 3�I3��$3�y�2�3Qǽ2��m3�n�2p��2�+=3���2c�3�D'3�V3Z 3`
03��3�(�3���2"`�2�53z�13��Z3�63C/�2��3{2'm[3�0�2��2�2���3�3�k�23˦39c�2��2'�3�E�2:--3�]3C3T3�Ř2�`�2A6k3�3f�^2���2D�3I`�2��2�}3{3��3,ޫ2���3��2e3�~�2�E3�3yJ23d�<3��2��3P�3]��2#�3�C�2C�m3Q��2���2ٶ 3��2�#3�T,3�;3�J;3k��2�]�2���3Y��2Al83���2#3͢�2��-3��53�0�23�c/3Jb,3�]3�*�2�>3��2���2eL35Լ2W+3�5�2+3��2�#3ˬ�2��3�z3Dh$3��3C��2a!�2e��2>zd3�X�2��O3U��3�w3U��2J��2�Y03���2CZ13p�-3C��2Rߴ3��2�^3�xG3�-�2���2Z�3�3�2̓3B�U3�{�2va3���2W:3�8�2�3�8A3��!3$A;3���2��?3p� 3߯�2�H>3�2��$3���2O�@3M��2���3>�3��3�:C3��X39�53��3t�+3߈3&��3ݜ3�73R�3���3�
_3��Y3��3�]3�143�uH3�Ƞ3��63g+�2��a36t}3�ڐ3���3��4x3���3��p3v�N3�4=3�Fj3Bǫ3�"3�Û3�Ҭ35�_3�~p3�H�2���3ƈ3��/3 .T3��3�p3<$3
�3��a3�x3�3�Y�3-["3R�B3�:3�h3A��3c�3Q�R3�\�2G�|3���3���3ͶU3��2J»3%�3do;3��d3F�p3�U�3�W+3d� 4lZl3�U3��3i�'4��3�Wp36�a3��j37e�27�33eD3���2�/{3w��3�!�3�O�3�A�22�3c�3��3��3�26x_3�'3���3.�3�&3pw23?�4��y3��~3�I�2��032�A3FI�3:��3��T3E��3f�3�3��K3ř 3܋�3��-3�=3��3ȳ�2
i4��/3�i�3ă�3\3_�B3w6�3>mb3�ܣ3U�3l��3�LJ3��]3�z�3Z��2;9�31��3_צ3��Q3�:3��3xv93��@3��3�3-�L3��D3�,�3���3/Z3}q�3�4�e3[3��3�\63QD3R��3u��3E[
3�.�3�n�3�yF3�n3��2~3�3OW3�x3�@3C+3?Y4r�	3�o3d[3��83(��2X?�37�3��L3��3mL,3� n3��i3�l3K�3�3:��3Z~�3�33}�43��3W53�3�ã3,��2V�	3�&*3Hy�3kHM3*�Q3��k3�=�3�OD3�{3���3�M53xx
3��S3�3]3#g]3S)�3�R�3�3F��3��&3�\3;��3(�L3yߐ3��_3ƍY3)��2͓�3�3�3��L3T�B4�:3��3ͷF3L�53��Z3��^3`�3}3ᵏ3M�3mh�3�1y3$�2�\3�Q3'-@3I�R3�j-3���3V �3U߽3�a�3o|�3D3�^�3��(3us3�3�$#3S2)3i�I3�3��3b�b3Z��3�{�3OKM3w�3��3Z(v3-�2"�3)�n3�f3u�2"v4�RN3�n3�3�@ 4*�3pU�3���2JF3�3��Y3}˙3�n3�>�3۾�3K��3)d3K�2X$73mZ�3�%3�rQ3�3.�03��3F��3�E3��?3md3>ذ3,_F3J�}3��2u#�2�RA3�:33��35�;3)i3I�3â�3.�2;�32��3Q�3�c53j�a3g%T3j�3�3��3$3z��38Hb3���3�}�2��g3�u3]�(3 !3\W3\�l3��2�_U3f5�3 C�3�#t3�Z<3��3}�I3�2-3"��3�z)3��3��'3@��3�e�3<{.3���2]��3	^G3RGt33+p3�N�2%83Pjk3�^P3��3�F3��3�9�30zL3�H�2c<�3ۼ�3���2ٱ�3��	3���3�3��y3�'h3z��3���2-3/4��F3�J?3�ZL3�mR3�%3�O3�OQ3L��2@�J3�4�+3c��3�3/3���36�3c=63��]3�L3��3�y�3�O3vt3���2?`.4�3�P3\�/3�3f3�243�W43x�]3��i3���3�:�3v��33�3���3j�@3GT3h`�3&�23��3�sC3M�3o�3!J3�H3��3�p;3�!3��3s�3��3�"�3�ӓ3��3���3R�4cF3�d3��3!3�?3���2�0f38S!3)�3�a73�Q�3�}D3�G3�03�4��3�;�3/�|3���3oE%3�R3P8e3E�2�E�3��3��~3�ד3|y�2S�.3j_U3`�c3�.3d�f3��l3jL3v��3���3u�2.U�2��&4LG)3 �3��H3-^3��63A�e3�Pw3��2�13D�A3W$�3/�E3�3.�b3.]73�<3���3'U3�>T3�3��m3��v34ߦ3:��3�3ž�2��3a��2�j3�* 3�F3A�[3l�C3��3���3��G3bb�3��E3�e3ggD3��	3T��3/�83��H3� 3�7�3�u03�.;3 ��3�w�3�W305a3"|�2�Tk3�� 3�ck3���3���2	��3js�3-��3,v3��3O�3��.3J3h#=3��!3�-Y3r�2�}�3�z�3@T�3�3u��3�73�V3�g39-3FD"3�;n3��s3��3�G(3#F�3�p�30_/3=��2�X>3ɺ"3�-3G�3���2�Yw3��2��q3�=3�a�3�!\3d��3�g 3��r3��2%E3�33,3��}3`2�2�%3�j�3�.X3��K3�0�2M�3��k3T+�2�q�3<3�2j�@3�I3��}3W�Q3�u3NI 3���3�a�2�f�3�rV3��[3�8�2�P3��f3�,3m�3ɰ"4�Zo3+�B3�
�2�H�3YL$3���2�8h3�+3�ރ3�+3A�3QIk3�x�3�>F3e�3|�P3Hiu3f��3�	d3%��2R3�m13�N�2)g`3oM�3\��3�U3@��2}I�3��36U3-��3�3�]�3Wu3��]3�E3��3�3̸�3Z�;3x3�c�2���3`�33l�|3��3t�3��N3:��3R�i3�.3+��2�*�3�_3��#3�H>3�"3��C3�U3���3�nQ3�:V3'�3���3{؅3�X37�-3K&|3Bo3|�e3c�e3/Z3?Y:3��3�|3���3*�3]�:3Ka�3�>3U��3��s3��T3|;3�(�3��Y3�P 3�>q3�^�37L3��13Z[X3�l3�T3in3��D3h�2 m3	T�3���3�s3|R*3H�3��3�
3x�3��3�~�3�I3_��3ΐ3#��2V�3���3��38F,3�d�3��z37U�2#�s3|�3��3�=E3���3ܶ�3�w3�3쐒3�O?3��3!�^3�3V3q�b34�2��343�$�3��3��%4GL3��3⼋3��>3��3gE�3��3�֖3.u�3�k4��3l@�3~r^3Jy93p�U3��K3��D34�y3�d�3�j63-ƿ3��3,ȱ3?O�3�<"4��z3�Š3.�3�-�3�Հ3�Ԗ3p��3��23�#`3��4 �3K�4ގ3\�3߫�3��3[w�3}�Z3��3,r3<P�3�L�3�3��Q3�;�3e�G3��3�{|3i}3��%3���3_f�3�3�ٗ3�B 4�0�3�x_3rX131��3���3Pg93�y�3�4�3R��3��3��3<�x3f�3�W�3y4;ݯ3�v3Eֈ3&l�3}�3:A�3ޱ�34��3zj�3��=4�"4�ջ3E�3)�3P��3t=3���3,g�3��3�D�3���3Y-�3�ƚ3��Q3ʗ�3�o�3Cg]3-�h3c͒3�=�3��3��3��[3Ô�3RY4� 4���3�]n3h��3���3�h3�Ŧ3�`�3j��3
$3&�3;��3�$I3R/�3�/4�r�3��3���3R��3�YQ3K�3��4�]3T�3)�4s�41+i3gT3� �3��3�$q3�F3z��3�S4N�3<��3"��3�^�3��/3=�;4��|3	�h3	�f3,.�3㖂3F3�3RX�3ɉs3,\�3�N4v��3��3�S'3m��3��{3�r3m��3�@3�m�3|�;3T� 4c+�3��3`��3��34�:�3c�3:��3��4��3��i3��3�	�3[��3��3�u�3���3�h43�!4	��3V��33��3i~3�B�3�L31<4��3t��3�[�3��q4i[�3�30ֶ3�~u3�i3L;u3���3��A3���3��64(K�3,�3Um03w��3R�3���35C�3�g\3��3�/3��4=��3���3|��3�I47��3<v�3f0�3Y��3��p3�1�3㠝33�"3��4�4�24R 4l'3Z�3_��32n�3��3��3�$4�^�3T�3�{4�Cs30��3�8�3h�-3֘�3V�x3�3��T3���3��3P�J3ɪ3�8�3�V`3"��3N13I�3-�3�1?3#�A3sd�3��3��3�$�3\��3<�h3��93EV�3Ğ{3���3}�A3���3�(G3�>�3���3��b3CKp3���3T�z3�ʧ3}�'3��B3ԅ�3��h3��3��3��3��3���3�8�3�߅3��}3M�3�f|3��-3��3cF�3�W3Y��3���3ޣ'3��e3�i�39ǎ3��J3�AH3�3�3t�3�
B3늠3'�"3<�3$0�3�9�3�=3���3�03���3-*3��f3� 3b��3(M3�(Z3�"�3V��2$v3�3]��3ц3,��2�)3N�:3�#O3E��3j3���3�|#3��3)��2y6A3�73=)�3�+a3'�Q3�WX3¡3	�o3�q�3q+�3]�2:�i3Y��35?�3m�3��H3k�3M�c3��2��A3^�x3.�93,3P:�3K��2}fa3��3b#�3�?�3EU�3\�3�qU36�63�/�3�1[3��Y3F3>݊3F�3i��3�}3��3!ٚ35@3W63�3��P3ԚI3Qܪ3�X3��W3OiJ3��4���3��3�13ۯ�3�{3�_3�T�3��3��#3���3	��3]�%3�s33^�3]3�)q3�4d`%3��y3zd�3Mh�3�3��\3�M\3���3_�[3T3�"m3K"�2��>3��)3Ξh3QJ'3�r3��3�x�3�Im3�R3�<�3��R3a��2��3_�B3�3363�K�3��30JD3H3�4�S3��{3��x3LQK3��b3�P3�3�TG3��3Z��3YR�3\�3��3砇3g9�3��o3ZΘ363�I�3�� 3'$)3���38lm3r�*3gJ 4^>3� �3#�V3�ve3�}&3��3�>�3�3Ș�3�_]3�5�3}�3��3M'c33��3��A3�L�3P�43���3��3�H�3�P�3�3�}31}�3�c3 r73j�	3�S3�3Bk$34�:3��=38V]3؃�36��2I� 3��V34�I3�]S3U�3Q�03�2~3��a34>�2و�3�K3�kM3�ng3:Ղ3d!3�M{3}[3tsw3��2��H3��L3��2�63��3"I3@�D3�Dh2S�93�!3�6r3@p3[�3�ZV3p
3��_3و3��)31c3�0�3�E93� 3�^p3�mu3˦3�3��J3�FP3c�L3w��3t�h3��53F��29�3nMs3F3�VB3��3�.S3��!3h�G3�643g��2�]�2�$M3އ3��2��h3��h3QZ�2l��2	_3�W3YC$3�Zx3M1V3I_3~�2o�13bFc3��3��Q36��2Mi3c�3յ3-�3$3	�%3���3�	�2��!3�BZ3�E3C�-3�^3r�u3[8�2�_j3��:3])-3�m3���2�P3��_3ĥ3,�B3t�2���3}W�25�T3��B3xC3�F%32>p3y;*3�d03��3\B�3�$G3���3
��3��2y>3.�s3�g3�o3�33��3dz;3��2]~q3ˌ3�if3�3 3��3�p3kӂ2��2���3h�3��"3k�2��=3M\3S̜3f3�83yyu3N�n3˃3U==3�V�222�3~�:3�e33��A3Z�03��13�q�2��43X��2��W3&�A3�ǯ3��3צv3��3��&3983$��3��x3Za3i�:3S��3���3��n3��2�`3e�%3)*z3��D39d�2�6;3xy3L�3��43_��2N�3��3w�3'13��13��w3��3��93�xv32i13cQk3Jb�3k/3�|E3�x�2��V3b�3&�3��j31�#3�ɘ3>��2:��3�Q3zv?3���2t&�3�5&3�R�3�3��B3�\3X3B�P3�{�2��W39�3Bk3���3���2�03��	3��3p\$3�@3{>�3�B3B��3�-3X�K3ШA3E��3`�-3�a3R�43��n3 \3{3/�M3�G3�2k�B3c]
3yT3�*3LY3�+3��3��3�.j3_�3���2}�F3���2��!3�U3>.y3��3h3��3�|13��2h�E3�3�3zGU3�kt3>)@3��3w��2J��3K�3F3��33�Q�2)�2�+�2!��3@G33>(�2EV	3��J3��3��33;�3y�>3��33���3���2Lm�2��3���3F��3�UB3ح2��c3D~�2�<�2֘]3[H�2m�3�}�3bJ3��3�ZB3�Ӆ3h��3�r3ƭ53�.43�n3�q23�
3�L3��2��\3#ru3Df�2��73'�2�Re313Q3�\i3Z�3$�63;��2��x3�>)3 �2*�33�~n3W��2�$3^�3bV3P�&3��;3�E3���2<�X3o�$3��3��63��2n�)3��3_"�2�Kx3_3J�O3��3��E3�3Ȭ�2���2��3^j3�43�*:3iK�2@ �2��3I�P3Mh39P<3r�b3f#�3�3�l�2��3�`@3�E�2fm3��2�<�3q6�2-w~3�1*3Kd'3�28;�3��T3D��2pO3�V83�	3[�23eh=3��2�[73�+�3�b3���2fM�2z �3�� 3o�2Ze3��2�3+3F��2�Qd3�333�M�2 ��3\��2Z�2F\3Y�&3P�2���2�/3Y3N~p3��3�:�3/�D3Ȃ�2j33��2JJ3%�_3���2�w3���2Բ�3��3c�H3$��2�3�3��l3y3�C23�O�2��2�[3*�?3U-3%5j3z��3+�\3�'3���2`3tv�3��03=-�2�P3�Lr31)�24k�3Rk
32:�26ǈ23�F3���2�!S3q-376�2s��2��3D3jv�2�)3���3^�03	133o��2/KF3�b3�%3�l'3���2քO3d&�2�l�3��3�Ed3��93߃�3� 3�G3�
�2�i;3��2�Va31g�2�"�2_V3-��3T�?3�ď3��:3G3T3��:3�'�2(̰2W�a3�3X�2��3��O3d��3N��3��;4Fvu3+Mg3�U�3՗3�$3�"�3�G�3��O3�3�30��3kZ�3A�t3ƅ�2��370�3���3�́3t\N3�A�3�GR3ź�3��3qCO3*o32�3ٯ�2ig%3�z3�9P3��83��,3E΢3�`30��3U�3ͶA3w�3��2���3\633�3�A�3'&3�ɕ3U43]�p3��3φ�3�Kz38�3�Um3��3b6b3h�E3�U'3�3p�3�M 3Q3�3j��35Ma3��U3�-3�5�3[�B35.Z3�s3m�83�F�3��C3Z��3�6~3��3��23�̭3#@3�M'3=-�3e�3��@3�Wz3�X3(h3%u�3�@�3�~�3ZF~3�q2^44D�Z36Q&3h>�3&^`3��3�I�2��3P�43�s33�E�3�w�3��R3�Vc3��k3;/�3�#03� 3�s3� 3]eG3&4-E�3�(3;Y�2/�3 u�3#�3��43�F3�L�3XY�3oU3Z?3�|93�+3[��3��E3��}3�bP36�h3Xtm3�?�3x�3/Z�2���3���3X�3�I3�� 3�63�I3� 3)ۡ33��3�+3�(i31�Q3�-F3F3/�4�{3���3s��2`xL3��B3�e30�!3��33^3�#�3y�&3}�W3�2�n3&�3DJ3%�Z3{3�$�3���2�m�3^�c3��3�AQ3*w�3.3v3s�3c,�3�73X��3-s3V�q3�ot36>�3:2�3��3Ʃ�3?��2��;3K6Z3N��3_sw3� �2�+Q3:;�3@>�3�۔3ܗ=38�&3�[4NC;3���3��3;b3�H3�WZ3�ӱ3��;3�Y�3\a~3j-�3�"{3K��2\�3@an3H�3��3"P.3l�3LeD35A3c�35\�2_�2%3�"3��73��3��2�73�	3I�2z��23�83��x3�L3a&�2�`3�?�3c	~3���2In3�2R3�D23�Q�2��3�,3;�43�!�2z�v3�֤2k�3W��2ɮ43��"3�y�2�3"|�2Q{,3�1�3��3W=
3i��2�30��2�|2�K>3M�2���2ß�2�p3�$33:��2�t3�3�y+3Q�38�3��2�~�2�s3ꍋ2�3��A3B�93��3��2Y�36�2� 3}J�2��2F�H3��3��93�[3�m3�R�2,6�3H3�"3�z�2Cw�2�.3�})3-S3�;�2���2@X�3���2:��2?5�2L�3�:3J�2�(3�3��3^��2�aN3��23��2�i�3��-3��3x��22��2��63�qA3�3-3钼2\Q3�ͯ3/;;3-��2�e�27�(3{�f3}c�2ah�2S#34B3p�*3�$�3�u&3�D�2��U3��~3��2rq�3ecE3��3	k>3�E3��R3�C�2�Z3q<3�c�34�C3�=�2�M3vׄ3)a�2823�?�2i��2��2�$O3й)3a9�2�i�23�3�63�F3D�G3�K�28�26�2m�3ZO"3j�K3�b?3^3�3c5�2��:3o�93��"3Դ3z��2B�`3��2,�3/O
3V�3e'Q3fv�3:�73��3A��2	)$3T<�2i/83���2���2,A%3)Ŧ3o>�3��3��2l3ֶ3�:$3��)3P�2���2�)�2�|�3¬3�#�2&>�2�Y�3`��2�d�2���2,J3���2�3x�3CĻ2o[3�83
_3���2�ҋ2�2���2ܞ�2ҷ;3.h}2
�j3���2�^63۶�2��2�޳2�i�3���2Z�/3p�)3vk�2��2��(3���2�G�2��k3��03���3���2M|�2oq3^`i3଺2�K3٦�2	KF3�N�2�HW3�u3�p�2{^A3�s3W�l3�
�2��=3���2���26�F3G�2���2J��2�<=3�w�3�e(3���2��H3i3s��2fS�2�3�O3k��2uPe3)?J3��{3�39f3��3R�;3Ev�3\H3��2��:3e�g3��2�73;s3�x63��S3l�2&d3ބ93(^�2o��2��2i3�3"`u38J13%�>3��3$��36
�2-=	3�e3l�3O#3��23�'3׎3'��2X��3W!?3��3i��2`FM3��3ݶ2%�b3!�L3�!3��3��q3{�%3�(398�2�3|q93�#3��3�3A��2��3|:_3��33��V3��r3�3���2�Q3|3z�R3"�3�%3ge3�}�2�H3z_3,�V3���2%S\3-33
�:3_�=3��=3fY3�SR3t:3cY�2��J3���3G�3�@)3](�2a;>3Q*3˹�2��3�
3�t�3|��2���3�r�2�^3��V3^%�3~+3e%R3��3i��2^
3O,R3	&3�2�>�3��*3Il 40V3���2H��3�3�&�2�eW3]3�2LQA3�~l3��S3<p37L3�w3�\�3=3��(3��2$��2Q)�26Q3��o387-3���3�@36��3W��2a��2��P3�� 3���2�zP3ƈ�2Y�c3�>�2(��3#��2���2,y�2fê3D��2Q'3Z�3qE
37l�2��2F?3�%�2��Y3.&�3��Y3�23Lr2rwD3�3�2���2��3�p�2@Yn3@c�2-ӣ3˭3>�2r3�K�3TJG3�Z53�U3z��3��D3��135�?3&t3|
"3�a3�m!3�23�s�2=3n�3[�3qF;3l?3��`3�U33*J3w�V3Mȵ2[�2�״3��03��93�; 3I�2P�3Tp3r=3��3��3�@�3�3�2�Y?3%�2+3�h%3��3Ӡ�3��2�3ڎ.3�43�s3l$�3��;3�C�3u�S3�x~3G��3=�I3�,3�?L3�o�3��!3�'G3��3]x�3�Ժ3��2��3��3��(3�/!3C�93�3�3��3O�3Ud�3#'�2�m�3�Z3�'R3�2�A3�9Y3��K3{0&3���3�t]3�2u3�S3J�|3�3 e�3�N3n3a3��430�B3��;38n�35a3�@D3OP3�"�3 K3-�3}�33���3B��2a&c3�ޙ38�537�<3e��3a�3��}3t��2���3J�3��3�I3�n%39x�3���2��3?�S3�3�L}3q�3�D37M3hk43�?F3�e3N�I3>ѓ3��3DW�3�)�3;��3�G3B�2]��3|3��3��"3�)o3N�3lC43��39<3��3���2g�3I&3�p3TD3|h*3�'38Ъ3�:f3h3/[�3{Ǔ38U�3y�;3EA23�n�3�W~3��=3�S�3Uh3��)3[3��3]5�2Ff%3�y23��3��-3TK3K��3�Po3��,3R3UW{3y��2l?3���3of�3WZ"3v�3��T3ץ53�3&,@3�&$3��E3>)3�y�3_|�3�Y03�:3���3$�32o�3�13�\p3`�;36�Y3*�v3��(3��3���3�SN3k$33/n3g�33m�x3tj<3�z3)p3)�83���3D 3l+�3���2�4�3�z3��3��3>�33!�3��73x�3�3�gx3:��3&�13"�r3�M�2��3�-3D�+3�y~3ְ2J��2P��2���3k3��3��3���3]�A3Z��3Y
<3��C3� �3C�3�o3Ox3��3X�3�A�3P�j3��W3Ori3�y38*d3��`3���2�W�3�K3B~�3@nA3<] 3�03+��3�>3�j3�153�?>3x3NF3��x3u��2�$�3a��3��3��e3�F�2�V3��3�3�2;�f3�-3n]�3��2�>4��s3k�4�{�3���3��3�?�3���3�<�3�M3���3�_3��,3F��3��04���3��A4b$o39�3��3��n3���3�S4�B�3ٌ�3��3���37�3kv3��<4��C3��3���3|�34��3��3|��3$�	4�\�3�2�3@7�3�<�38�@3 ��3 �3�mP3J)}3k�3�M�3�3N3:�4�ɐ3&h+4�1�3O�44 �4d�3q49��3��3�v�3u,4߁�3��3B!4���3�e�3���3Uv	4���3�-43���3G�3�%�3���3k�4��3Y�3���3h�c4�+�3zK�3�w�3�4b7�3���3�x�3�lF3X�4�l4]�4�X	4!��3�^�3&`�3'�3�ˊ3�2�3���3���3�6Z4=a�3�i�3��3[�4Z4�Ђ3�+�3Դ3���3��3�{�3/R�3�#4&�4O 4���3B�3���3
ˁ3U~�3��3ο43Zq�3�	4��54�3�ܱ3�`�3�4�?4 ��3��3�y�3.3|�3�4��+3k�3t�4K��3p�3B׊3²E4��4;4�2�3f�3DZ4�3�94��4�3��3�&�493�3��3;.�3I��3��t3n�I3.4|��3U�3��@4.5�3-��3z��3��3:��3ʭ�3(�4!�3&�37�3��
4��3]\4�B�3y�p4W�%3Mb�3��3�Ɲ3�'�3K�4�Z74^�3���3N�B4P��3�{?3�K^3Xm45�3��n3LW�36�a3�4��3	��3",�3е�3�A�3�b�4�ޝ3�i�3�R�3;��3���3���37_�3�3^4$��3�4�@�3�X03���3=�4i�?3Dҭ3�p3J��3��3�l4OJR3��3�fZ3�-s4b}3��$4�t4���3�Ư3H��3�e4v�3��3v84%B4�-�3FU�3i��3���32י3���3r�3�X!4�O�3c4eJ�3���3h�S3�u�3���3��3N�n3���3Hߘ3�[�3$�T3(@x3]�[3h�3�i�3ZÒ3F3H3ڙ�3�{3���3N�\3�!3D3!ƺ3��3*{*3
�3�@�3J�?3���3cBa3Ϣ�33mt3N�{3J�3{�3:7U3�ʲ3|d�3�3}!�3�4���3Z�3.n3;��3���31�3��3�@3�{q3�b|3h��3���3Te�3�g3��,3ɰ3L��3��4{��3�8�3D!�3`Y�3[�+3I�Q3,i�3Π�3�E03�|i3�2B3�3�3]c�3���3��-3��63F,4�v]3ɀ\3�K3���3��c3��J3o�P3c��2�Er3���3E;�3}̎3Zz�2���3W�q3>�(3|:�3�i�2~�V4�3��3%�n3�z�3��+3.�H4�~3�|3���3Uk�3I3�^i3�zP3�/'3�?�3�M�3X��34��2�Q3i^�2�m�3"�}3�Vq3�d3�3&�!3��3
e83��3�Au3D�3��3f̨31�3�93�q3�Uw3$J�3N�3�mI3?a4#M�3:�r3'e3���3�W�3�zW3kX�3P�3��J3�E3_��31�B3`N(3,%B3��4R?\3x�3�m3>"K3�߁3��H34�3�{3B��3U��37�3�X�3E03i�32e�3ی�3��3��53��
3�(3,��3�l73k^^3�&O3NZ4�n)3�a3�>3��`3�03��3z{�3�%3b�.3��3o�3�Ɛ3FK3��3��3�03�3=*�3�C�3,3r�u3��63�9�3S23��4ܘ�3��3۲3���3�"3��)30�3zs�3s=4��4�@�3���3�k_3/�3��3h�3e��3�3��b3j�,3�ۚ3��B3�3��2���3��q3��@3���2��f3<P3@X�3��3E�3��<3N�3�_�3�U�3�w3$T�3p&}3�
3�3�3���2 ]�3}}03^��3��O3{��3ɮ�38��3J@3��T3�@N3���3B'3���3{�b3�53m�a3���3;��3�4�3��3���3-�w3�3i��3��3��3a3lj4��g3���3�L4yU�3�'3�ڿ3�3g�4	��39Ra3j�3R��3Wx3\�3\��3c\�37_&3[ˇ3��3�q3o�g3.3�Ў3n-{3�յ3�a�3l٦3�]w3`W�3�\3�bJ3�E3�ɣ34723~�3���3U��3)��3�a4Ư�3�hQ3=�3���3�-H3:�3�ϯ3M�:3�N�3F6�3�
�3�^�3q�3�5f3��4��{3�_�3�Y`3�X3��31�N3���3ՀL34aZ3?��3�%�3/�/3�H3P>Y3���3�7�3��3�Y�3Y��3}�33�  45�>3Wnq3b�3$>A4y�x3��T3��3�R3]�M3���3P��39�X3�T73U��3݀�3��3s�3s7�3eTC3Q3|�3�V(3`�d3�v73iɜ3C3qa3��H3��4��3��3!3W�M3���2��3���3t�2�!3���3_6�3�3\��2]��3n�3jq}3˞3��i3�ͪ3���3�0n3���3��3�*3�&47�3 X3�V$3g�3���3K�]3��3��93��n3�S]4f�46 3��+3=��3�>�3�}3���3�m(3V�3*��3�E4��n3�xn3��2�n	4�AP3�w3�A3)�3�sn3�ƙ3e�3�/3�3�V
4�*t3���3T(36xg3�`�3��r3��q3E�,3r7�3o63]��3g�3SP`33r.3FB4�)~3l�3-��3�Q�3Ic3��`3�/{3qm3ZX3���3��3��3\2.3C�3��3�_�3.0�3N)3��3��37U�3#�V3��O3��37�34E�$3�֑3�e�3��3��93�p3��3ˇ.3�g�3��3{ޕ3�nx3:)3�/"37�3��3	�r3��932�39�3�w�3��3���3b4�3��3Z�y3��3�eo3� 3�(3�!�3T��3a��3�z�3Y�p36��3(X�3��]3���3)s�3��*3X�i3�d�3|�3��w3�45��3�?y3���3H��3��3�Wn3bgk3�3��3<�3�2�3��'3.��3���3�D�3�t�3LT23s3L>3�f53�y3~:i3���3	z�3
ļ3�؆3�	�3_��3=�Y4�x�3�<3���3Ϻ�3�K3�43��3[7|3Q��3֗�3Q��3~��3D�F3y�3�v3)c�2���3�N�3�n�3�Je3h�3I�L3��3�5)3"B4�|a3���3��o3�F�3��U3��i3ݚ�3L243H�3Ͷ�3���3d�3τ@3i��2�ڨ3K��3*��3(;;3���3G3��3�^h3�mY3��93�}�3�Bl3�*3-�&3E�:3�?S3[H�34��3��U3"��3���34��3�l3��3-�3�_f318�3bs3(�@3]ȑ3��C3<�3�ې3�<�3	�30]4��\3db�3w��3���3�V3B�3��o3��_3`�|3K�3�
�3�م3�J36��3T��3}C�3C��3&�D3VW�3є03r6�3��c3��L3�B�3 4g�-3?l�3�u�3E�3�e3��3�`T3��#3ϯ�3���3i��3?F�3E0p3Fק3$�{3۶�3�wa3�3{�3���3��3>��3�o�3���3��4��M3��3�=�3���3�XQ3C�3k��3�/33č3"�14o�l3�є3U�B3`��3z]3���3Q��30@33S��37��3֊4銉3��"3Ҭ3-��4=��384�3�3��3���31j�3��q3��3"г3���3s �3pҷ3V��2�k3�ú3�e�3E��3�ڂ3�4��3c483�3�[93�5�2#j4��3��3�=j3�Rl3�-B3��.3���3dTj3A8�3���3��3gh�3F%3G�f3
:o3�13�ʎ3oJ3�/�3E`3���3�i�3��3��f3���3�CB3�|p3�N3߫�3<53}.3w�3�N3��3s��3*}z3]�!3��J3s��3Eb3̴3�3[�3�3���2q�3�L�3���3�#'3� �3�d3I53e�~3�n�2	�3�=3�Ms3�2q~%3r��3o:�26F53p��2��Q3�[+3�s3��I3�K�2u3�/�2<L�3�I3i�2@��2A��3륆3��3h}�3�W�3[�[3D=H3"�D3E�3��/30�3���33j.3�,�2O�*3��)3e��2DJ:3;�'3w�3�c�2^A3Y�^3�DL3,��3c�3h�2��D3�a3�;3�j3�t3[�3��3�23�.�3��3��93�<#3K��3��~3�F32�#3X�2H(Y3,��3�a<3�33�;3��2! 4?��2��/3�39�63A�i38%�3�JH3H%3��\3Z��3��3�N3m 3�pm3�?3�2�`U3���2���3��O3�x�3��2 V3
73#��3=f�2)x3��N3�]B3�OF3��3B6J3�O3&�)34R�3�G�3��p3�63`�A3(3G�o3�'>3�3S3	$�3xpE3AJ�3bDW3Ô@3�[h3�U]4�ig3g�3�9H3��3��3/Ł3�?Q3{&�2��-3Ii�3�/�3eP3�3zb3;�3zE3w�+3�n3�^l3-@'3{1A3�CV3�P3X��2��04�73>��2*�2۪�2�r3/^3΄3�3��M3�ˉ3�mN3�};3���2��K3w�b3�2Fe3��'3��X3J�H31��3�vE3��3�J3V"4� /3J��3��_3��"3�y3,nd3��#3�*�2|�/3%Z�3܆�38T�3@�2��2 ��3�B3�3�#3Q��3���2�Yk3�Ld3�>3��3�;�3r>a3P�3��)3�'W3���2Y3�'�3� �2��3�I�3��3��]3�U3!��3aZ�3RC,3q�S3��,3��3��<3߼�3� /3��3�{3@��3f�=3�h�3e�3�{u3�3���34q�3�Eu3�3X�4�k�3w��3.cb3Hn�3��3K�w3Th3��3�_3�X36��3��3mU3{*v3G�3g�3\:�3�6-3��3�E�3Z��3��3w�o3p��3U��3n�m3h7�3\93���3���3��3p�3Xت3
�3�&3�W�3�zD3l��3��3�4�aP3t��3�:33�[�3�O3��w3�}3�NE3̾L3Mޅ3�r�3�/Q30�2��3��3�-&3�Џ3��K3��Z3�jP3�@�3��l3U�x3��3��4
E3*Oi3�~"3���3��F3��d3_�3F�?38%73#��3�?�3~ �3E��2k̤3�A�3�	H3a�3�`E3�C�3�(U3΢�3fd�2�9Y3&�J3�S�3c}�3u�q3y3:3\Y3ʽ�3�t�3�V�3hb43>�a31�3��R3�IB3��C3�o�3��a3�33~�3ͥ3�j�3M�3u2�3�@]3p�k3���3���3���3�F�3��3x_e3�2�3;_h3���3��c3N�34=Ā3{��3�~3�Q4)��3|B43.��3#��3 ّ3�E�3�X�3zk�3#]x3�r�3']�3�O93�`#3�օ3��z3#3�013b��3��3��3�"�3���3b�P30a�2�$�3��3�X&3_�k33��2#�73OdG3�\3��j3 3�3�W�3���3�F3�t3��>3��l3�(83J0o3zՍ3�t73'Ր3���3]�3f*3�$A3� �3��|3�*a3iC�3X3�ǒ3��35Ɛ3y3 ,63�03(04j�3	Vv3|3��y3�.33�"3��3']�2 f�3ɮ�3x��3�ш3��2���3P��3�x83┝33h�3X��3��3��	4>��3�ta3>o3r�Q4��*3E\e3�9�3N�h3�z3�{3�3x3�p3"��3�m�3�{3��2��3�o3#N*3"w�3a�2��v3��&3�2�3{UD3�v�3���3��3tNT3�YU3DH�3�!�3 ^3}��3.V|3�E3��h3���3��3��/4��3���3�1�3d�3�R-3�bg3��$3��b3���3��d3��K3�!�3�A�3R0B3u��3* �3b9�3���3iҀ3�`3��@3|S�3�u�3��3��3
S3���3�93n�3Ӭ3��+3N=n3��u3�;�3�q�39��3W�3�[�3u��3�$3�^3��32�,3�G�3�$�3��37T3+�3�jG3�F3�E,3�2=3�ry3�1�2��N3׿3+w3u�.3Z��3�A�3�k|3���3��40M'3�Hp3[$d3�x{3r[d3�r35פ3Z1.3�x�3�H�3t"4$(d3ʓ 3���3�oR3�>3�}�3G�3��3�<j3���3Ν^33�y3��H3'�3��3!��3k`Z3Y�m3�r3q#�3�O�3̩&3��L3�*�3�g�3p��3�g*3n�3y�3�zs3	ҕ3(��2���3k�3;��3�QQ3	]�3�_�3f��3ٜ3L��3_��3�Ud3�63�bF3#D�3!�3��3���3�e�3Z3 33�h3�Dt3��O3=3�3�]3`��3J�S3�֟3��2ѿq3B��21�\4��Z3�~�3�=Z3�7f38`f3kw3���3��3$�n3�ͤ3��3��)3}�e3s�3X�37�3hX`3�j3Iw�3boc3z%�3�k'3(�3��2�+�3 b3O��2�2p3�Qd3��2Ɠh34�3x&93�!`3_��3���3@�>3��2G<�3�gG3(73�{&3v�#3���3�g�2b8�3V*3�l3�S3� �3E8�3��3�ۉ3� ~3|� 3	�@3X��3��o3�s3s.�3��3~�G3��!3�	(3�+\3�l�3���3��33'�~3�<3��3ag3��=3
+Q3X�3U�3?j3���3f�G3VN3�DJ3�3�d3�ٰ3�3o�3�y3]��2��3���3��P3ʢ3�234�{3��&3"��3�L3�3�3\��33`�q3�-H3��3�e�2A8638�3�36�K3�ˉ3���2=�s3)3��03�Q3�/�29��2��B3j�	3|t�2֮�3��93#3ý3 0�3v��2�=]3��3��F3J�2���3��K3c�2�< 3�Zv39c3�3��2��3�H23�>�24 3b�2j�C3k��2�c�3�`Z3[�S3E��2Wj�3"�J3�j�2�v3�3>3j�3���2���2r�%3�z3j%~3�W3u�2Z�3��O3Ο�2S3q��2K��3���2��b3���2�T3�g3
@�3���2��e3\U�3H$:3΂93g�3�13�m3�3ӫ�3�t3>&3��2�?E31��3�E3s�O3_�:3p�_3��93S�2�_3|W�2��2t[�3HV 3	3x.3N�03�3d�B3z�S3�Q3bU3��3yo�3�{?3�A�2���3��Z34��2�:J3��3�F�3�,3\�P3�3�J�3�I3L��3,�3z��3vU�3�3�$T3u$3e�3���2��J3�݃3)�3a�`3_b3��3j�3���2�P3��2_�_3��3sĄ383�@3u8�24���2|gZ3|M3o�3��3$�3zTk3�3>Bq3cV�3?�?3ɷ3�!3�&3M��20�27X3�3�3(SP3�]3�!�2��39V3��3�P�2���2I�#3�mo3�535\�3av3��2sz.3��M3n{�3��3H��2UT3�3�2��3&x43.4�2�VM3��3��3�*33��3F��3�A3��2�7�3�@|3C3Ʒ�2��Q3���2�3��O3��G3,��2ߋ3V��2L'3QRd3C`
3���2�J3���21!3�33��2�8k3���3}7�2��3�3!"73�o�2)3�`3�]�2��:3g+�3�x36��2K 38�R3@�B3N��2G�;37Z3���2X�J3�^�3�3��3!3�v3Ұ3�ZT3r L3/),3{2���3�7>33535�{3C�3y�Y3�E�3��3�3״i3 7�2�l 3a�j3�4]3S�2��3��R3[Ԁ3_�13�p�3"�3�h3�c=33"�3˹n3\�3337W3��3뼲3v�3��3e1�3�3q�3@�35
83�Ü3��3�k3N�L3S�=3!�%3��4�3��83��3h�W3]B3N$-3��3ر)3���3ց�3	˝3S�3G¬2wH3��53��2��U3�2�|33*e�3�I83���3��3���3�o83 q 3���3���3��+3��'3��3��3z�D3,p4�lt3+F3�83k�3�8�3�|3V�K3���2s�3���2mC�3�w3��2̮�20	�3AX3�!'3G�,3)P�3?3�%3e�'3��2'�?3��3�E3-�_3���2:dH3k��3���2wt�3&�q3p�63c�2-�X3)}_3���3���2�
�3�+R3šE3��V3j03ܣG3U�c3��n3{��2��3�X�3	�3�g3R,3-�3�t3 N$3+7Z3��33��3��3;��3�>3��D3. 3���3~�3tNa3�_43���3��2��V3��J3�.3�^3l�3��a3"��3�f3[G�3��"3u�&3-8e3l�53X;3	�3��3U�M3c��3�V3
4��*3B�R3��D3��2��$3(lh3�\�3s$�2��3F��3�y3Z<3%3��3���3���2��3�13!3Ex3�(�3�w[3
3�!@3~_4p��3�39�2��3e3�\�2Y 3���2���3��3��3�z3�3N�3���3��2233k�q3�"C3C�2��4��#3��3�C3 ��3.�3� =3M+3��M3�Qy3��j3ax3��2)�3(�3O#�3'?	3�z�23�A3�3Q�3rBw3{�2u]?3��l3.g�3`
3&˾3!�`3MR�3�@�3�3��W3E�34�m3��3$Q3�7�3�cq3�%!4�>3�E�3��$3�u35�3��&3�Gl3@*s3`�3ܸ-3 �3\�3�w�3�{3��3��^3рZ3�c3��3T^D3x�3;W3~��3�ݸ3���3�g^3��{3���2�H�3��C3�)3��3�L3mP�3��_3c�3��2I�_3g�)3��54z�_31a3�_�3�/}3L��3?k�3�X�3��3�o�3�[4�^�3�Rb3#33�C�3�vl3��Z3���3�z33hm3T��3�н3��y3Il3�3ױ�3gn3��3cE~3�D3r�B3T��3�J�3c$3���3�F144��3�4h3��?3+˯3#W�3z��3�v3�3r��3���2[�3H�_3Q��2A�3cd4� �3�FO3���3��F3�)N32�A3��4�73\��3���3�V�3'�3�,3�Z�3�f�3[j3$��3�h�3�֪3
��3)&�3;|�3�#93/�3�3�~�3$��3���3ڬ�3��~3�ˢ3���3��3`�a3��3<=�3��G3��3��4S;4��;3�[�3}{;3ɽ�3�J:3��3��3�n�3мd3�!4�#R3wl�3�f�3H1J3)D"3�բ3|а3��3ab3�@4�/�3�J3}3���3Տ3�C3�Z�3�A3���3��,3��4{Z3݄;3�V3��34FR^3�8�3�o3��3��3��t3QN�3���34��3�n�3Q_�3DL3mf@3ghs3AF3#�?3?N�3�O3,%�3 ��3v��3�g�3٢�3�K3}{�30�q3�H�3�%�3:�03�O�3�>H3��3C�3�U�3�.4��3�ӗ3чk3m��3'Ȧ3n�t3��(3��@3i� 4e�d3[��3W�3��03a30L4�Y3�Ҹ3�5l3��O3�M33��3l��3R��2�!�3��3yݞ3��C3E�#3s�Z3rUL3�kG3�Ov3�Y3Q�c3�ǐ3͒�3y�k3;��3�/3啅3;;�2P�3`G�2��3�%�2�`3M�!3��&3���2Z��3��+3��3خ2K�V3��3��3���2��2^lF3�=�2�-3�> 3�GH3]��2��3�M3!��2���20�3ź24:3�3A�2��2P��3z�2��3t��2�d%3ڙ)3;0�2��3�!03�B3[��2�F3�w�2�*�2�f3�gd3+3��T3���2�~f3��13��d3U�b3�+3��2|3��[3��3�83��"3��`3ZRZ3�Dp3%!3�PV3w<'3��f3r�,3�!A3p3Hp�3N3A�2� :3�o39�2�%J3n1H3���2��%3���343t�
3���2� P3t�2_�#3._�3��2=�43T��2�[k3k��2�13��-3�~v3�Q�2'2�3�?F3�T-3>� 3�;3��3��2� 3%�x3y�]3s�2U��2@W[3m�:35X*3~�3i�3PA3n'*3{63wB3'�k3%w�2�`�36[	3P3��?3n�&3��
3Њ3h4J3=<|2�p�2*�3^g3��93�;3�pT3z�a3��~2�2lm�28��2�V�2�S=3�93�/33�3�ƺ3
3�J3�M3�Oi3��3��D3�O3���2 �/3Ś3yOf3�C�2�a�2V�3�3L�F3��63�#.3�3�K3ʘi3�,3�L3��2E�3��>2�38�!36�2X�=3�3,�Q3�F3�q3�ҋ3�P�3�!3)�3�83;��2l�2�&3Oҁ2�iF3�NI3�٬3\�63L��2w	�2#Q�3�3��3� 3@j	3`�3,�3MiT3��3�}$3&��3�{]3v@23�{�27��2��3Z��2�3	��2"ɢ3{	
3W�c3�#3F]#3{3���37�3�+�2��3�.�2'?
3!>3��43?s3��l3��Z3���3��.3�M�2��
3��(3!3��V3Rf3mȋ3?I3멌3�8%3�E�3��k3e�3�H�3�173zc�2j��3
{3[�T3��z3��3E�
3b��3�а3&�O3L�)3�1j3��k3�>3��2�E33D&36�2j��3��f34~ 3��3���3DS3�d�3�oO3ٍ3��3e�v36�o3T�3~b3KN$3�I3)��3�`�2頉3*�31[�2A�G3)��2�!U3�83���3��83�|3rMH3ҡ#403R�N3�=13հX3��3��%3�u�3��K30�3�6�3�z3BO$3�$3fC(3�D3��
3�]P3���2z?�3WG3	�3w�?3�D3���2��!4Â*3n13��	3Yt3���2��^3��3���2�`�3�q�37��3m�2���2�.3�o3��\34�>3���2A�3T3ON�3.{3��3|-3��3~Ll3�I3��3�33�A03F <3n_3��2�3�λ3���3�A43]�43�h"3,,P3{3��:3�̹2� S3��+3��3t3��.3�\3j��3�(3�ӈ3Xޥ3v�O3p:Q3@�3-�M3V��2�.3��&4D#�3$�o3J37�3��w3SO�3�k�3�31��3�v43�L%3�t3^H>3��3�D�3۽N3 
3�K3u$R3AG3�p3��3�)=3�b3���3(N�3��3��3���3\}3
1w3Z�m3+�2_:3\r)3���3�Q3���2�+3Pۥ3&c�2L�b3�߅383�G?3-�b3�CL3�.3�"b3��b3#v�3��3���2�,3/��3Fb�2�zz3�{3N�r3%f3�Pc3�0A3�G3r�3k~3�m?3��O3���3�3ئ 3_;3h�z3���2��43X�3{f�3��3J%3�3��[3K3�3Ư�2�N�33(��3N�33(3��2��3313�Qa3u�a3�c3(�X3��$3�z�2�>/3�Ά3�I3X�3E<�2�=34�53�^�2�ۉ3O/�2�ܗ3Hp�3Ñ�3�f&3��4�\3���3)��3�;�3��A3���3!eM3�Û3���3�~�3��93;o4�\�3RD�3�%q3���3L��3��B3՜^3v|�3Um�3*�	3wX�3�|�3�d�3�~+3֑�3�o>3�\�3|��3/)�3��m3�4�3�b�3�zW3�<�3Cv�3R��3���3X3�X�3f��3��
3�/�3�5c3^��3ryN3�3�~�3x�i3�ʋ3��3�=a3��3(_�3�Q�3�35rU3m��3� 3�-�3^<$4�	4Ӯ3a3�Q�3���3'�03�̧3��Q3���3�|3���3�DH3n�]3%_b3��j4�}3�G�3�e�3ɻ�3,��3���3RJ4d�A3;<4�y+4�1�3�1�3�5!3>�3Eۜ3��$3o�o3I�=3UW�3�Q53R�3z��3k�~3:vw3sJ#4���3�9�3��S3���3_tB3�A^3��3�Ƣ3oҪ3#�P4�]4 ��3ԙQ3-U�3�C�3:33�b�3v��3�S3�3��3�Z|3/��3ݳh3�	4Gv3�3�64�J�3��{3Y8�3�30�3���3 Z�3�{4_ũ3���3��3�3Q��3E��3+�3�2�3���3���3��3��3>�3�"<4(d]3���3��3d]�38˱3yo3��3BR>3-�3�d4��3�d�3f©36E�3��V3�(�3�I�3Z%B3���3��:3hP�3���3��3���3�b�3"�"3�u�3�w�3⎄35��3َM3���3��Y3�T�39�	4%�4M��3�U,3���3���3�{J3h�3��3��e3�+�3TW4JJ�3�m~3��S3q� 4�:�3�2z3��J3Z��3{DM3�f3�Sq3Ga@3���3�O�3���3�Ë3Q
�3�)]3v�M3|�3p��3Z3q5�3`]I38��3/�m3΃;3L�U3�84:v�3��3lR�3�4k3�r�3�f{3�d�3�tL3���3�~ 4�3�(3j�{34�3>�3�3iۃ3�\)3�ґ3���33�3
��3v�%3!��2��V3b&3>t3�P$3��23��2�&�2*|�23��2��T3E��3�3+k3J�3�(3�5�2�wj2ԉ3�3��3�3KQ,3V�3�C63�%"3��\3�I�2�$3�>3k�}3Z$3�z3� 3j:�28�I3�o3���3�Ǖ33�2v$43	�,3��2׻}3�2�i34�2�h3�3��3�3�A�3�e�2��03*ŵ2��3[S3�Z 3�(3� �2�$3�32�3���2�W�2�3\�28�2Y
3q�2d��2��2x�3<Y-3}�e3���2��h3 �3 �3��3�k39�2��U3��)3�0�2��G3}�^3�A3c��2�@�2�c3��3.3�3��2q x3�*�2d?�33.��2��03t�3��
3}w3�'A3h+�2�c13��`3�j3ˡ�2j\[3r�j3��k3HO"3���2��-3<wK3U�2��D3F73r]37W3�O�3�<�2t�3T^3q3#3�(-3@�!3Fy03R�3�	-3y3;3�2�3��3�\�3��M3t3*H3�3CI�21<3U<�2F13���2W�g3ʁ�2���2��3�Y�3 �3�3��3\K�2̳�2	h.3)�R3z�
3F�/38s3 c3(�3�1�2m3U��2d/$3&_*3��3�113fH3>�y3�.�2�i�2�2^��3Q�3�b3w� 3��"3lҭ2�3�� 3Tʞ2���2U�3.�B3a�3���2*03@��2�2<�"3l�2�p�3�3�.l3<�3�3�l/3ˍ�3�u�2l��2��2�|3з�2�E�2�A3R�3873ڡv3D�53)�3tN�2.H<3|i�2\uR3��2��2d�o3�3�2OS#3��2��3��3��J3�L�2S��2Y�33ҭ,3���2>�R3eK63�ך2�3�fz3�%	3��T3B�2�2	3F�03��2z Q3�3��*3l�2��h3NY73R��3�8�3��3 �3�@�35h3UA`3�
<3��3N#�3;��3,)3��3��4�۝3l�E3DW�3z>C3� [3��3���3�1�3�H3�x�3��3%��3e��3�լ3�vI3g~�3�3���3mǔ35�^3���3pp�3@{z3,j�3<�3.u3��I3�W4׫�3 �i3��3���3���3�]�3!��30y3\��3[[�3��%4A�3&.�3��c3;s�3��3�D�38��3*�3�)�3��4>��3���3QE3;k�3���3S="3]d�3d/k3��3M��3l��3?oi3̗�3�Bl3��R4r9�3ܦm3���3��3�\L3ү�3�"�3D�/3<t�3�#4Κ3�)�3`V3���3`��3�G3�̆3ؓ�3�|�30��3�&4j��3щ3��3�\G44a�3��3dY�3<�=3��3�M�3���3�
3���3 W�3ǐ�3�U�3�]3�}W3#-�3��O3���3�=3���3Y�3T��3J]3}�3ۦ3�k4�;�3�L�3Q�3>��3ZEB3��3���3T�,3�v�3�x#4�3��y3�b3WJ�3 q�3���3�i33L=^3y��3e<3uO�3���3��13BrW3iU4��3v��3��3"��3��3׵3d}�3(5k3 t�3���3�P�3!�E3�53K܋3�K�35�E3�o�3�3��3��}3d'�3v3��3|�3`!4�v�3~�3{�s3n��3k��3W��3��o3�z3�}13F�	4��3�h�3��R3��y3��U3�P^3׿�3�3���3���3�C�3{o�3���3�~4��I4�3�3�0�3��3�X3vE?3{��3A��3��3WLn3b�-4`��3t�3�$Q3+9�3#Xo3M� 4t�$31X3]I�3/Q�2/��3�3i�H3� 3r^4-�p3Uh�3���3莤3��3�o�3�Ռ3fw39>�3TS�3L�3/��3]z3�y�3̑�3�ա3G��3v3!3!��3�Ɔ3���3��3��3J�3J �3a�3��3��3���3�c3�:3B��3hS3]�;3!F�3��3�O�3L�:3���3
�3��3;�A3k_�3�Q�3%T3Ⱦ�33�3|�3=��3r
	4�Ĕ3VV3�[3A.b3�3��[3�J<3��3e�Q3���3�ذ33J�3��"3�:�3�ݙ35 �3Y�3K{�3��e3�3�v�3�I3��h3�CM3䚃3���2��L3^3�Z93iKA3e�36)�3c�83�8�32<�3��3��3�23e��3M�C3x�2c��3�W�3Q�73�6i3��3NT?3��3���3܀a4��3LȄ3�us3<�3w7G3���3^��3��3q�3(H 4܀�3u39�	3uٕ3�143�8K3���3� �3Z��3�C3j��3�Ҋ3r�?3qq$3@��3�(�3�^3=�@3���3��3G�4B(�3��?3��k3�n4%�3,��3#�?3GŽ3��35��3>3�3#N3|�3
�:3�f�3�t3{�A3�ӯ3���3�j�3�~63W�3]X�3VW3�W3���3���2a03�4K��3�ŋ3	xm3���3�.�3�f	3��03�2A3rx�3� 3uݒ39�h3��N3�h3�Y�3�{@3�3j3�e3���3�ğ3ʇ�3��M3�Ƌ3�U3���36�3�{3ȿ;3P�l34��3
Gn32�3��l3eu3uqM3]h�3^x3��g3*�53�q4t�v3�k43b�M3X:3�3mt�3��3$�32��3���3�+�3�\Y3�y236ޱ3mv�3R�3���3��3
�q3>Q@3d�4՝d3���3iq�3�F�3�н3)8�35��3'�3�ך3��K3�sy3�G3
͞3��4}�4!��33+3�b�3W�3� �3���3��#3�Х3�V�3�@�3�V�3m�}3�E;3��4{834�K3�}+3L�3:�K3�K�3�f�3��03m�3N�3�~�3soQ3+
/3K��3�QQ3��#3��3\Y73�`�3�u3	��3�>l3���3TX�3[C�3�{3ߌ�3�z3� 3w�53�0�3�g�3��3��#3L�4Q��3�P�3|"�3�4;�3SwP3��<3���3�i�3E W3���3���3�S43��~3K��3吃3ʠ�3�m83ߗ�3ZB�3���3؝�3G3��S3���3��37W3+f3>�3R�#3,�3<pv3{�3��3lC�34z8�3A��3,І3C:4�/�3�?3U�y3�#�3N,.37�3��3?�3��s3��=4���3�]�3��3�U�3sm�3�sI3���3	�A3�N�3��G3�M�3X �3��3�D�3���3QZ�3ő�3���3�i�3�1�3��-3�ȳ3F7�3g"�3	�4�d�3��n3W{�3��3���3��3��3=ň3:�3���3�>�3�ޢ3�~�3<�Q3gF=4�C�32��3@	3	x�3k�83��3��3��T3��3�4P}�3F�h3��E3`Ʃ3��3rPh3j�3I�V3�G�3�5E3���3]�3�o�3�5n30�45�3�S�3�m38��32�a3���3�2�37g3\_�32�34�04�3�� 3��3�\�3��2�!�3��\3o�3�>3���3�Ń3籁3�yf334�t3:��3~��3H��3�o�3�=�3���3��d3ꪍ3}��3�5�38DY3�M�3�3n�z3�mc37��39�b3��4�0H3���3��+3�U13gR�2�-�3�[�3�3��I3FB�36�D3�,�3E�3Oj�2�O3�1�3!�3�bF3c�333%�3� 3���3��2<��3�`�3��4>�P3�!V3��3�)4��y3�<#3��3�h}3�Z3O�h3�@�3��/3j��3�"�3�&�3I_�3[<:3�0�3j�y3��3x��35�73Տ3��\3Y/�3[Ls3��L3�3���3T43W��32��3?3�3�mn3�ʁ3r��3�r3��3�v�3]C�3b�3j�03/Љ3g3�]�3DjN3}�3���3H� 3��3�٣3j	3�a�2��3�3�aO3�r3LN+3��3�T3I�*3�'�2��2�3�]3�Æ3��u3�*�3]d3W��2߿h3}�03o^�3���2�m�3�!3փ3��3�M�3w�Q3$#p3D�3��[3�a230B3�)�3�3R�31��3��}3"l�3�3/o@3�(o3bM�2��3g@3S�U3��2|(�3߀3$du3[�2�T@3�W3)n}3�13cL*34�31G_3��63�0+3�v3���3�!33�C3���2��63��i3Ҕ�2.N73�`�2��<3e�3y�d3#�3��g3�x�3F�3�,.3��P3j[3��"3D�=3�C]3p� 3�+3�3�g�39��3�3�;.3��@3�,\3��:3��@3�
$3���3�`3>/$3�34�3wQ�2
�3��H3aȀ3���2 :3@e�3~D?34oJ3�z 3�$S3�i�3��L3zj3� �2y*g3�.�3">O3?ip3<�2Q�3$y3'�f303��3��3�.�3��3��B3��3s2E3��h3Tc�3<��3�� 3�P&3�n�3�đ3�33iH33�3��3�l3Qǃ3��3���3=T�3�3w��2���2��3a�4'�!3��N3��&3�V3^�3)E-3��3��)3+�<3"��3���3_�3��2��u3��3���2>Q3^��2�Ux3La�3�:S3���3�,F3ԉ�2�3yt
3{�D3�$3�-3K�356�2&�?3S��24/3�[�3<3�&C3�2e�93"3�+3�d:3[��2�(3��2x|3�$N3%�3#e3��3&�A3u"3s�3c�2n"�2I�G3�K31K�2�L_3�&�3㠟3��o35��2Pg3U%�3"�/3�/�2+i3�,�3e�3[�4�d{3L�3��2%�3�*3�`f3:��3ئ,3m�2�s�2RK3�P3~X�3�3�Hf3�	s3�A�2��(3ˊ�3��29̓3p)3 *w3�.3P�3f��21^�2~{�2�?�3��3��+3�#37aN3��P2k�2��2�q3N��2R�)3,�T3Nr%3ē�2�R�2a^3�_2�Ѫ2���2-�?3݂�2��L3!3�d53	��2�R3� �2��2���2���2��2�*3 �23g�2JY�2��3�c�2��3N�2���2�ĺ2���2�3r��2�3��3�{�2\�2�I�2g��2�zq3˛�2�23	�2d"3~Z3~D�2i��2{3Wը2�Y�3�X3�7�2�M2�8W34@�2ڽ2�#3�#r2�y�2AE3`B3�#3�783��3�,�3ڻ2m+�2o��2b�2�P�2O�+3(�93p��2�]�2�3���2��2�ue23�3tD�2?7�2���2��2�;N3�&�2B�3[N�2���2L��2_7e3P��2!*3:'�2��2hʣ2���2x\L3���2]3��|3[$�2pf$3ѣ�2���2��3}{�2��3G�
3b�$3ٖ�2*�@3q�2O��2SP3�;3:��2 ��2�?	3�t&3*}�2O��2[��2r�n2�$�2��@3�_#3e��2�j2�4<3A?3���2@3�8�2�_�2�f�2��-39��2G��2Iб2��3ֈ�2$:�2�t�2���2Bx�2.̰2�M�2���2l'3�K#3FCg3��"3��^2O�3���2��2���2f�2 32�2�V3	B�2VZ�2g�2�f�3d:�2e��2� 3St�2�`�2xD�2�3$�2Ǯ3mH30F�2��2
q2��3�h3v�2�R�2�o�2g�436�2�3��3$��2̥2u��3��$3���2N��2���2���2L�2� 3�B2I 3�V3�� 353@�Q2$��2��+3�,�2���2�$ 3N6�3(�k2��"3e�3�e�2���2
y+3�*�21Q:3��3�/�2��2�1�2�3d��2F�3�
#3}�213$F�2��3(��2���2�3�Ѩ2��26�2,�3$|�2��3F��3Qy�3��g3�(�3�qt3�E�3���2�41ak33(3�i�3i��3�v�3�U�3�3
33�3�O�3Fe3wߌ3��3۷3P�2��4;ĕ3��h3yn3u��3���3�E�3N��3&U�3��3~��3�K�3k�3oL�3xiq30�3H�3)��2��3Mj}3ŝ�3��3��3}��3g|63
A�3! �3�b3�M�3pu#4�/�3��{3�AJ3���3�Q\3V93���34�3�S�3f�,4?��3���3?M3wR�3��3	�G3O��3��3��3P��3Cb
4�`30�3j��2?�4m3nS3AŅ3�3	�3>}W3;p�3+*3���3���3���3�_�3t�&3�3q*�3~GP3��^3n�!3*�4���3��u3DZ3L�q36Q�3� 4�}3b��3xt�3�rw3�t3~��3p5H3�P3�3rI4��3ĵW3��L3�3��3��_3��u3sO3��3�)53+��3��=3��p3iƂ3��4T܃3��3���3ߡ�3z~�3��3���3�%3k�3k�3x]d3믋3.T�36�47��3�V3Y�3��^3�$�3���3q�31;�3P�'3�@3�aH4RQg3w3>^|3b {3��X3�uq3Fp�3���3�a�3US�3g��3B�u3I��2�r�3�g�3��3���3'\�3�|3iV�3��4��93��j3���3%`24bR_3@,�3%F�3!�+3U4'3�E�3��3�483n��3 �4'p4�3`�|3��4�u�3�h3n�3�?3���3��[3K��3"M�3^4�3�uH3�=4h�3r��3�3i��3��M3�a3UM�3�C30��3�U�31��3z˿3f(3q��3���3Ev3h}s3�`3�b�3_V83�T3�=�3��3|��3��4��-3�&�3=�
4&�3��33��3�W�3�j3�3+��3h�3���3�C3�z3�]�35:N3�g3���2���3��b3$d�3��3�&�3��v3� 4�Z)3�43�!3
c3��3+��3��^3�"3tw3䡨3��3�a�3�3�3+1]3mL�24��3��3��o3���2�cs3�f3C,@3�Y3��3�'3�j�3Dmg38�83�L#3���3��3�nY3�6^3���3� �3я3��M3�?�3��T3��g3@�h3u63�E3��.3�q}3z3�%f3n'934�@3��Q3�3�<U3q 3:;3�R�3M�%3�	3%��3���3#�"3��C3+�A3dր3ES�2m]3�QF3�|3�Kk3�y�3s=3(�3�3��(4b��2�|c32>3��3fld32�93�3	�2Ϊ3Z�4�t3�a3_��2�O|3���3K��2���34�
3�9�3�N3�5Q3 ̠3�n3�03��4�lI3���3\3�+�3�3$�3o��3�|X3�'�3C4�3���3 �h3Xڀ3@=�3��}3��3?��3 LL3�F�3�eO3���3�93�q3�2~4J��3��3e��3v�v3R�3۸�3�3��3TX`3���3�Ҵ3�6J3>�{3ڀ3�k)38V�2�#�3&n�2���3�3�Ď36ɫ3rQp3)�Q3<�$4��=3KI�3�03ԑ�2�W�3cF�3lr3(+3�3P��39o3�.j3K.�2���3�3��3��L3F�2N^�3��c3�`3�,3�B[3;6�3�=4�MW3�,N3,L�3`�3��A3P�3��|3͊3z�23 �3���3S�l3��3ĳ�3w�M33fA�3%3��3`�13��4�P-3��G3��m3���3h=�3K�3a��37�3/�3rl3M}�3l�b3�}�3µ4G��3kS3GB3�'�3o0�3�Λ3N��3��3ǧ�3fb3��3y�3E�2x$3Kv�3[�3�Z3�'�3`��3xR 3|`3�/�3�'3�q3�:�3A��3��p3s"3%�4^a�3�>�2$'u36&3��{39W3��3!�3���3�3�i 4��[3ݫ�3�]3<J�3`3�c�3�ى3DR�3��)3c�3�#�3z��3��&3�F4�uP3q�3|<�3��g3�)�3��3R��3�y�3�	>3V6�3ʋ�3��3ۀ�3�Z
3�*{3?��3gљ3��3�+�3�m�3<�3��3���3h�!3�~�3,��3$o3K�3�i�3g#�3�p�33��3��Q3��93��3/1�3�v�3��3m��3��3��2��L3�-�3֎�3���31~43��3'43��3w9�3\�o3��3	��3�o�3t�<3�>4nk�3P"y3�)�3��4q�-3(_!3{E>3�"3.�3�p�3S��3�3�+[3��4WL�3P73��>3
�3>�$3�3�c3��L3G5�3@ �3�{4ͼ3[=3#�T3��4a��3)��3u�3G��3h�e3�t�3�Z�3�4�3܈3��3^3�d=3�j33��4�4j�z3���3F��3*4�3M�3�F�3�k�3�l3G�M36�3S�O3�Zv3�+[3�d�3�Q3Z�3r��3�1;3GF�3� �3�g�3� �3��+3�Ĝ3M�3��~3q�3Н03���3.�M3�u�3<�3 f3��W3/84��3��4���3�h31�]3��3���3�63d+@3�ߺ3I�k3��3�3e�4}J�3
Q�3��3�,3/n�3�6T3lB�3�ʹ3�"�2e��3�43� 3`'!3J�q3k1�3)a�2[>�3���3y�3�+�3�Z4���3�3�M3��3�6=3v�@3�*�3�483\��3}X�3�k
4�36D3N�^3�.4	�3���39?�3z��3��G3~e�3l�3�Ė3y�3���3�e�3__�3�[.3�e�3k��3���3�3*�R39��3p�2ׯ�3��3�v3�3G��3P53���3�,3�Ad3y�L3b��3Vʯ3A1�3{�3��*4�-�3�aZ3�=Y3�+�3MO3�<3u��3Z3�'3��!3���3I��3��)3��3�o�3�E	3�(3��3v�2oܦ2:g3�f13��3d�3YY3`��35U3mU)3�+3*E�2��2�L3�P$3��M3���2���3�|<333f�R3Jg�2ʸ3*�3�.3���2�/3c~3���2�!�3�۞3��3�{#3�e33X3�>3�3�3[C23���3�#(3��!3ԢU3//B3�"3Gt�3%3�#�2(�3k�d3-��2Mi 3ȷ_3�!3�[13�^3�.3���28è2�LX3+-3�3K��2�I�29}�3Cʾ2D�u3?�L3W{3�3\�I3U�2�03�X�2hC�2��2�C�2Db'3�T�2�NT3���3��33&Tq3�{ 3,�53c�3Qu3��3D8/3u&3�y3�H�3K�3+�3z�/3 �4�"23y3��3�}I3��B3��q3�܁3 j32F3�O83%d3,�3�}�2=�t3�j3�E3��q3�A�2W3�/3;�}3^�23aqL3OL 3���3�6�3B 3�3��S3���2��G3�93�i�2	}53k��3�x73�3��A3jbz3q3F)3��^3�b3D�b3�O3�l3�I3��,3���2���3X{�2͝�2���2S��2�#3�'g3D�T3lO�2Na\3i��3��3�&�2���2���27l�2ȝ�2��>3�83��3#%3��f3�"3Ln3Yy�2�3r��2�T3�s3��?3��2��2�
U3��2��3��3�"<3�[R3([2�g/3��53���2��2%A�2J[i3���2S��3�i�2���2!�2,�4�SZ3���2:�B3k%63j�!3ћ�2|�3��2��-3�*H3��3�@3wo 3��3q�j3���2�%3�3�3F��2�i�3��63���2���2n�4�3��$3�U-3K��2rVF3��d3)J3��2j�J3�>_3�3��s3�$�2}�3'ܵ21�2�G3$�2���3*~"3W�73q�93�O�3c��3]�3��3�x�3l�l3	��3��M33��3���3uDe3�R�3z�4���3�={3�ds3���32vU3&aY3fҟ3�Y�3zt�3�3~�3���3�)�3:J�3=�+4�#�3���38�3ц
4��3�w�3 "�3�P�3V��3f�3���3��3��F3��32�4Y��3��3�63��3i3G��3@l4���3�Y3;!M4EF�3O��3��3��S3���3C4�4��3^G�3ֽX4�4�P�3��w3��3>m�3��"3_�3I��3�d94r��3�D�3A$�32��3a�3+�x4vm3�A�3H�4��n350�3���39�3�M?3���3��C4"�47ֲ3(�]3�S�3Ş�3��3`��3q$�3�&�3<H�3Xw�3K��3"J�3�۬3��!4�s3x�3M��3��b3�zl3�V�3�4CVY3���3�404���3۫3)��3~��3Û�3c��3w�3�zU3���3|/3�4Y�n3�I4.`h3�B4��w3���3H��3�/�3$y4��36�3� m3#N�34�04���4s�3O��3�n�3M�3�K�3dU�3>J�3,x�3g�m3�Y�3��3�C�3�3��42�3��3U33'�3p@�3�]�3׾�3�f�3���38�"4_	4]�3��.3���3l �3h�h3!+�31^}3�m�3���38��3 ��3��{3�P�3Ü+4p��3ю�3�6�3:s�3yR�3ȗ�3��4���3��3�b4��4ة�3�1�33v�3)�3R�3��4��`3��3Br�3uT4���3��3��3;�?4Zs�3�*4�/4Җ�3���3�+�3t�3���3-X4��48�?4�@94+<�3cZ�3q94A��3�k�3ܠ3�j4��3-�4F��3�3�X�3]�y4��3	ۨ3L��3M>3NF�32��3�~�3><�3��/4�9�3�^4<-4Q��3�p�3���3H\�3M��3h�V3~>�3;��3��q4Q��3��24�o�3-Q�3��3a�3��38 �3�;L3l��3�o�3��23���3�(�3�#�3w4�N�3yR�3�Y�3��3"EW3��4�<4��I3��4bV�3�R�3䀎35"4�Q�3���3�,�3�	�3G�3D��3b��3���3�f3/��3"�'4�\�3
z3/+4��31�3�&�3��3��4p��3@�3�¶3�m|3Y�3��U4K��3/��3��3v�y3E>d3Y��3?�3�s�33�3���3�;3צ�3C�	3�)�3���3wd�3�р3 ��3A&4���3�7�3�0 4AGB4]��3x�4m )3AВ3Y��3��3~4�3��3M4ꨘ3Х�3��E4&�#4���3WaV3af4�N�3D�3j��3�$�3K� 4h��3���3�t�3;��3���3��34�3	�4n�3�i�3���3�C4=c	4ѩ�3�B�3,�64��3:�3��w3���3gj�3jn_3��4��3���3H_�3�S�3���36�3xl�3k�4�ּ3�_�3�3��3P��3�s3��3�-<3�_�3�4X64<3
4��?3)<+4���3�0�39�4&ů339�3���3N��3��D3C�e3��_3۟4@jv3���3C��3��14\��3�>�3���3ת33�s�3��.4(t4�<�3#o3FH�3U �3���3N��3�2d3~�4��3�+�3K�f3�Ϛ3#g3|T4�}�3ip3���3 �3�V4Xl�3�!44#�34��3�j 4֖4$�K3E�64��33�3��3��3�R�3:��3���3�Zv3�3R��3�D4x��3'�3�54u��32Ʃ3�N4��3ݧh3/��3�X/4��3��74\�|33(�31LI4p�3F��3c-�3J�"4e�3?�3+��3tEW3�8�3ĝJ4���3E6�3��4�0m3.qW3�j4_�3=3�4�z4�O�3b��3H#C3��^3�n�3g��3�^�3�OY3���3���3���3��4��3 b3t�f3*9M30ּ3�φ3<��3�,36�$3,��3!V3�9
3+_�3	:�3�Sa39�3���3e%3^-23�>X3f��2#��3C�E3R|�3+��3�h3�v 3	�3Ͽ3�3c�3K�/3��=3��r3ք�3��e3��U39��3>Z3���3y*3���3UQ3�u93�`	3���3PM3���2� �3[x�3;�83�y3^�3�3jh�3 ��2�҈3�,�2b�.3�D3p�I3ƙE3�:�3ӭ�3C)C3D43���3Oo�3)�3F�3�k�2���3�W3�k3c�[3$tb3�@3���3��V3���3��3��O3��3)��3�x�3��?3��N3��3�up3R�3"�33�]�3��(3��3Ĕ3V�j3�`�2��3d(�21B�3ɏ3�7�3e�<3�3�r[3,�13`�z3��:3㝅3gv�2�Ia37H�3''�3]J!3�6.3f�3F*3ͷi3�؂3�)3Č�3��I3�/>3!9l3�7L37-73�,�3O��3��n3��W3p ;3�1f3ǌ"3�ŀ3���2l�Y3ރ3x�3��s3�33k��3�O�3�/�2g�b31�3��b3�B3�FH3��^3vo33�k33c�4��3Re83B`3�P3*�3�Ι33�i3�/3�}31Ճ3敭3k��2�@3>5�3+3��3�_"31ji2���3�_3���3~7K3�r3NAJ3DQ�3�!3�t3�X33(ҁ3��53��s3��A3��M3��a3̳�3�h�3�m*3)h�2��L3�=C3��l3�i�3f)3��3�<U3i�3�.�2�c3�޺2�e�3�c�3�cg3��&3C�!3�3H�?3�z3l�3:�l3�-�3��3��_3r�3��w3���3;�h3 �*3�O-3�2�3PJ	3渱3ܸ�3ڧ�2���2��	4ю3��3�.?3=J/3�23	�E3߽)3j��24��3Ĭ�3�3�b3�Q�2��'3���3H�2:U/3�e3?d�3CP 3�r�3�3���3��2��33��2&�3�3�S�38�2,��3�iE3:�3X�E3��3��f3N�j3H��2� x3��J3���2�i3��G3��i3!�2S�3�.3�^B3v`�3��3�b43��-3�ZD3a�N3�9�2�-s3*�L3�e�2��p3֡�3#�3�!�3��3_ܗ34q.3߉L3<�L3��3�2�3��3�Ԥ3��3���3��.3�)3T;?3�:3;qI3&�31�3�&�3k�u33�38,3¦ 4�=3� 3
�2��3��3=*�2ΰ�3N�3X03Mo~35�3l7B3r3�n�2Ȳ�3<�F3E�^3��3:Z%3���2�mc3��3gp-3G�3�V�3��3��T3�H3,sP3�\K3J!33�e3�"3O��3ۙ33_��3��31��2�m�2$��3�/�37�,3v�)3 g3��<3f�;3ZqE3i3-t�3N�t3ͬ�3U|63ڇ�2���3��|3��F3���2]�<3���2��83�5�3�V3��3��33�v4n3B3�M�3�v3��33C38�T3�Xx3x83'93�L�3�q3�*d3h�,3�Mr3�Α3�Q�2D 3S�"3�dO3�+3�W3��83h;23J>@3��3�Kr3s�U3աE3;�E3�3_#P3o�3���2�!n3B�3݂�31�J3O��2j�3�)G3��`3� �33k-3#(3
3[��3>�3�.g3c83}�35.3Z��3J��3CPs3E��2tW3H~3�_3v$X3O;y3���3|��3р3H�Y3�H�3}3�}s3�,3�7�3?x38�3�<�2Z�u3wK34_tX3(}`3�+N3�+&3�9;3��3u��3	�3�Y/3� �3fG�3�N3]p3�SO3�^�3.z*3�>3�u�2뢓3�q�20;3)�53d	�2�3���3��2��M3�+3���2-�13��-3>KN3f�2q$^30��3?�|3L�%3��43ͼ�3Y�D3���2@��3�h�2�Z3Օ�2On�3O�'3��3��*38�3��'3�� 3�4�2.4�3P�3�W-3��3�O�39EJ34��3�
�3k0�2`3���3t3��2D3�c3#3)��2:�T3��'33Y�3�qy3db�3��m3Ӑ3�0�3N��3�w3�r�3PZ3�B�3�q23B�3��3�"�3�-�2��h3�Pc3U�C3m�3��Y3ɽu3�3�JO3�Ƀ3"+z3F�3 ��3 ��2hC�29UZ3Q�63���2-F�2S�]3���2�l3WA�3�Gx3s�2>?�2���3J13%-3R=�3�x!3lO�3��*3拼3�aB3�h3�;3��3�|3��3��-3f�E3�3�383}ω3o�3��g3-�3�M3}�93va�2E�)3�(�3��\3w;3��3���3�S3m�b3"1q3�V3�n�3D%�3��3�S3�߀3�B#3�<�2�Ň3��P3��
3�;3�%4��3g�O3�23t�J3ܛ�3$�3q(�3�%3��3�3Xc�3g��3��J3߅/3%�*4Ǝ-3�3(�D3
�J3�[3��C3�o3��2���3"E�3@H�3/%03b+3��B3)�f3��(3I��3= 3��3���3��E3q�.3��j3�03���3WVX3�},3�n93z^3)233�}"3(ZA3�TW3��%3�6�38�c3��13�T3�م3BT3�/3�33di3��o3���2�L|3�33�ʒ3_�,3���3CP3xvr3�[3	L>3x��2���2�ג3=�2 ��2Q�3-��3.5�3�3 "39I3�O=3��u3��3�\3�83հ�3&B3V�I3�_p3���3�33C�B3���3*kC3�j/3e@�3'_3c�j3�Л3ky�3�4Z3�kV3��~3(�~3Q�*3��3a�3�X03�7d3R�	3�U�3`�H3��#3 �3Mk�3G�2�:3tk3�L�2'\Q3�<'3�VF3V��2��i3���3s�3ΟY3G� 3��3ˆ?3��21�3�s3g3Z3.�83F�3g 3o�3r�2�O3�{�2�H�2��3���2,�2+�2��3&Я2}f�2�=)3;@3�93��x2�+!3nf�2�=2�<�2GG3��2���2�13c�"3۲�2ޤ3�3a�2|m�2f�2b��2}��2�x�2&��2/g2���2$�3�3w�3���2��L3}�22�3l��2�L�2�� 3%�E3���2��3~7�2�Up3��2�T�2��
3��2U
�2+��2ϡJ3?h�2�/ 3zP23I�3d�3.M�2Ƶ-3�3oa�2�}�2��2��3��
3��3jw3cJ�2v��2�!a3�L�2���2���2�f�2y�2U�3z3���2£�2ő3�t�2{g�2m2ϳ2�+�2k�2#u�2O��2p�i3�x�2�_3Bk�2� �2���23D3�,�2��R3��|2�{3���2
W�2�!3:�2�+3��3���2��2ZЙ2�>�2~�2�4�2B$3Z�2}P�2�D�2ȓ13��2T`�2���2|/3��3+��2c�)3QV�2���2�D3]�3D�12���2˼Q3��D3��36�|2zt#3�ZH3�!�2=k!3��2<3/��2�3=��2���2��3�[3ܔ2��2��g3��R3,�2�3��$3��2ag�2�3oct3c��2���2�3q��2T#�2��3��2U�3���2�/3_M3�V�2�r3k?�3,#�2�2��2���2Vk�2W'�2O3Ƶ�2q`3$�3X�3J�2�d�2c�&3v��2� 3��3���2c��2��29�H3��2Mz3E�2��/3L�13&<3��2	�3�3�2���2�C3�A�2��3�ű3��%30�3�"�2m�2���2��2�f3hy3Y��2��w2��3��3\b]2��S2� �3�B�2��2k�|2��3<��2S��2`*�2 2>2��2X33� 3ۊ�2�)w2�D�2|��2��s2'��2:��2��3���2�+3b��2��R3�3�'Y35�L3Lי3/u23=�3k�2<�C3��93�6/3&,�25YT3�D�3���3�lD3;mj3bz3��#3��3
ac3j=�3���2�߫3�t=3(�,3?G<3}�3�<3^�\3�b3���2��3��,3���3��53�g3e�x3oi�3f�j3���2ǲp3�z;3�K�3�h]3'��2q$o3H �2��T3W+3�<'3��3��3��!3*
f3by3v>3��3��3�193�3cZ�3-�%3J�36p3�w,3�Z�3��c3d;33`q43x�3���3C3�d3(	3�QB3�a3��3�3*|�3\��3-43�A3��.3��3�(3tUR3�3䖆35�'3���2���3��C3��3�?�3�3k�}3��3���3F*3�G3)n�2��3A3�d3tQ73e�=353,3�Ic3q�R3�>13���3zߔ3�8U3�Q3���2� �3�uJ3)3{��3���2�3�>#3Ρ3}US3j�83�qG3()4�R3�#3�3�q�3h,C3�X3�D3��63Xw�3��3k�3]�G3~o73�\�3:ˀ3���2aJ3�413�V�3c�a3�n�3��u3��3��13��3xnH3��63�gv3�Ct3�q43C��3)7a3�|�3ٸ93��3�P�3���3�3��G3/�3�Z�2�mm3�o3>v3��3�/�3�XA3Jۤ2q�3[?�3��3�Oi3�Q3H�w3��3ͷ#3�S�3w�-3v��3��3ڵ3X
3&��2Vwq3S V3�-#3]T�3P83׿3'3�b3�}83_j
3�Q3��3_n83U�2��Q3ԯ$3g�(3�AD3��A3N��2H�3�EL3�)�3
fZ3�Z�2�?3f�3 d�3��3�2�j�3�J=3y��3)+<3�؏3��/3 R�3`�=39�\3"�{3=jI3��30t43�h3�3Yg*3c:�3��p3O�3��2��T3��G3h~,3�53A�2�!�3�13:�>3�3��C3��354m3�T3k�3>'s3*1~3�{ 3z�q3=73=$3[1P3�4��3I�)3�3�2_3���3zP3��H3��C3��%3߼N3z��3S3��n3F�
3��38L3�DB3t�C33vv3��-3��3�"�3�y�3��;3Xu�3�r�3@=�3�M�2�q�3���3:�73.��3�&�2aUg3�<d3��93v\3t�3>3��e3BZ"3�73B�3�-�3#�3���2u�3je�2w�(3���3L,�3w+S3i�2�R3L�3o�E3Cg/3��-3Tq�3\t3炄3I3�j3�L398<4�)3��3zcr3�H'3��3��V3��u3Q"3�?�3�P�3lE3q�3�2��V3mo3��2x�3�[3�33H��3m�?3��&3���2���3/>03��\34� 3.�g3M�3���3��q3�]"3�	'3�j37T�3���3��)3d�`3��43�6T3�[�3�ˡ2Wh�3��3��F3�?m3�#Z3y\3�&4�3#F3��<3Z53��2?|\3�Xm3Mw33�H3{9�3ui�3�7�3�`333��3� �3]�v3�u$3�p03�i�3�gs3�G3�323��C3�c�2�*4h�F3w*�3'5y3�i3���3�>3��3Uh36Y"3���3-��3�3�>3�G3z�3:�,3�E3%��2�J!3>39��3H@03�~�2:"@3j�3Z��2�H3]�3)`@3���2�;3��3�t�2r��3���30��31�:3�3 3�N�3�D�3��+3�%D3�6*3��[3�3Ն�3>X3J��3*s�3ŕ�3�3=3n
d3��n3�g3n3��3��%3yCQ3.X�3B��3V��3��3�J�2�,.3�a�3Q\3��.3;�3��3��S3a�3�X3�q�2}u3���3��t3��2�c3
X�3�n3��k3P��3��F3"x�3*c�3�M�3r�)3��2���3�~B3�B3�73�3!k�3H3G3�@�3� �3Tc�3`�I3zV�3 �g3ZO�3T�G3
y�3��j3���3��3�Rt3'�3q��3��3���3�393� 41u�3ŉ
3��@3]��3cѳ37�}3�5�3)pu3�r�3s4�j�3�S3�y|3���3h�38�3�Z3D��3�(3|_o33�3�>�38�3r�;3��P3�ū3��3���3��3�/,3r�3���3�-�3��r3�+�3��3���3�f�3��U3�_R3`+�3c�3���3؊�3�5m3�K4d:�3�H3H}&3V��3l�\3��;3Qu�3���3#�3���3ܻ3_��3�^�3�"�3��.4D�&34�3�ԉ3BU�2�5�3�35:Y3,�l3Oh�3eq�3��3��3��2���3t"�3�M�3w�53��3�/�3
�3M��3��Z3�Z3�3M��3.�r3X=3��l3�a�3AM�3˴3� D3��@3�є3�=�3���3fTV3�o3�A�3q�3�8>3F*4Y�3���3��3��3�Ld3��2�2�3��"4�|+3��Y3E��3wʊ3��431��3r��3�a3��3�4A��3�f�3�w�3Ш3'��3�.D3��3f�_3�g�3���3���34�v3h;�3�(43<�#4�P�3%_�3t��3u�3�IY3�n3زr3l*C3�(�3'�4���3��3o>34�h3�σ3�G�3���3]�|3�4Y��3�u�31�3'�3�t�3U:4�N�3.�w3N�3}́3�|/3a��3;ʭ3vh3��3��
4��3n��3�83s�p3�hE3Gb`3~�3��3�Ǐ34��3G��3��3�hR3J�3?�4$C_30۲3��3j��3N��3�Jc3�Z�3�KN3��~3(4���3�e�36�I3Mι3A˯3�P3 u�3��M3�T�3^�3E3�3*0�3�FU3K�L3C�*4�J�3���3��B3|��3_�]3lЁ3,T�3|N3i9�3��3Σ�3W�3F3�3_��3bȣ3�
_3��83s��3�3MZ�39�3k%�3~��3�4���3��R3��3��36:3��3��3�=B3�t3F�4܃3�i3z��3�d	4κ�3�d3�I�3�M�3��N3q�b3�θ3j"o3�Iy3��^3��4;�t3��3��3��[3R3��3���3�w�3
��3�n�3��3K��3�gI3���3���3�^�3�8V3S7J3%P3 �3�u�3�#�3ڣ�3�_3��3`H3pUX3�y�3/=�3�G3�;>3|KY3I213��\3D:�3�3� 3�'3���3O<?3�h3�'�3e�c3��3$�3a,�3G� 3��w3�m3�G	4��3H��3��3ڍ3>g3X��3���3�mF3ĉ�3�U#4}6�3@[<3��s3$��3�\3�q`3?�3��"3�:�3Q03iD4��3�f�3-�Z3�#4��3�;]3E1�3/��3�OW3���3#�3�3b��3FAX4�M�3K+l3w�x3��3cN3�<3μ�3/(13�ۜ3$;l3�J�3��s3[v3SU3JN�3��l3�Ht3�V|3l	4}m�3Kn�3��3;�3���3~n�3�7�3S��3���2�vg3?i4h�"3Q��3R�i33��3~'3T��3��3�W3��B3�24_	�3jeT3B��3[3+B�3��m3ȑ�3�n3#0�3g4��3��{3�53~V*3�`g3n�o3�5�30�q3���3��32�4��k3@iR3��3~u4�%B37��3�k�3�"�3^�b3\�3���3�3�n3�;�3�3	�3ܨ3yx�3}��3�"D3��3r(23�w�3�D3_�3E˂3}l30`%3��4ij�3C;�3W�3�E3@lT3'q�3�I�3���3
��3�j�3��3�Ⱦ3?  3Ƨ�3j,�3���2%�t3,`{3��3V6v3o�3��3��W3��32�S4�5�3���3�G3���3SfN3X�3'�3d�3��g3��3͏�3k�35#�3Vg�33JX03f�3��J3Г�3q3_3Y��3��3%��3m�K3���38�83Ԉ)3�&3��3���2��,3l^�3�b 3�4�2i�v3��`3��A3��@3(*3	�V3��2+�83�0T3%Dn3���2���3��3y:3�ُ3�3m�63t�32![39H3�.3�,�3��E3�rA3*�W3�	�3�*3��-3��3�e#3�N3e��3�=3�^�2��3��3s�b3���3�F3U�S3���3v.$3
:3���2��3��3+ӂ3�?W3�tL3�"f3���3�mZ3�˫2|m3�Kx3IdD33�+3��33Qe3Ϊ43J"�3��23��3�>3�N�3^3�r3��v3�?�2.y33�H3R�v3_�2�433�E4D�~3#M3�21��3^P38�3%1+3yt�2�J333��3��3 ��2?-T3�i�3 }3ڀ<3en�3�kA3���2Z�U3� H3��2''B3׃3C��3�3�	3�0�3K.3[��2r�I3y3�2283]^3��j3S
N3�S$3,53���3�L^3� C3}I3�̀3	p;3Xbp3	�d3�3�=�2���3ճ�3�WT3Zd23��M3�Qz3�_�3!��3��3��3.=%3�g303r^03u��2jн3_XV3�r53:�3ՓJ3r[3��3�9z3�X�3V[�3`��3=3�3% 32��3�
F3V��2ͅ3�/3�ő3X�3!҉3H/23�S�2o�2�i�3��!3�M]3&q3�L93��!3Cx�3G�t3�>�3wϲ3��3�K�3��3>�3r�3ɡ3?�3$�3�]3v��3�t�2�ڼ3���3�Ή3&g�2F4��A3z�P3�fB3�>V3uV3>�H3�o\3�j�2�R3RK�3�%�3P�3��3԰3�҇3�C3�H`3���2���3�2[ܒ3��=3O/53p�435KU4� 3��3��A32h*3�T�21 �3�p�3[H�2l��3��3&�g3�53���2�u�34�3 3�L^3�&�2�'�3��)3��3LTw3�y�3z�~3��3�Ø3ys3Z�3"�3x�c3�P�3�ka3>�F3%P3��!4�r�3khO38��2�3���3�:�2�C3��W3�U�3f�3�W�32]�3�cO3�ey34��3,�39�G3T0a3ײH3�.63h�o3_�3��43.>p3u�3�4�3�c�3��!3yp�3�N~3�}3P�3�R3-�R3ԃ:3��3[IQ3*�O3SpW3�4q03釁39�.3��3>�3Љ3�Q31�^3�zs39-�34p{3�Th3���2zĚ3�
H3��&3�f�3��u3��3kDa3$�3I7&3]�W3��d3ܧ3��03�J3H��3�D`3eT3��3�3��3I^^3e`*4.��3�93}b�2�p�3�x�3lO�3i"�3�j03��3Ԗ;3�C�3��r3l��2��<3b$4}�3�e�2�#A30Z73��s33�[3��l3^73#�r3��3+�3w�_3��3lW�3F�T3 �?3?��3��3&�3��93�3ICp3H�m3k(3�d�3G�n3�|3)vz3��Z3lVQ36�V3�*�3�[30t�3g��3�S�3i�3^.3ٜ30�P3H3��3�33�-�3��%3bM�3���3~�43�3G�3
�239��3@@�3�673��>3���3��3�p]3M�Y3ʳ3C�4�^3�P3�W�3��-3��t3���3J��2l[�3�"W3t�3�*b3�XU3�Y�3�#�3�?x3�
m3BK�3A�3Xe3�1H3}��3�Sd3�!{3�\4�6�3�ev3Jj�2�̵3.;63 -3���3�$3���3���3��3_*X3��43��w3�G�3�h3Ur�3��>3i�%3�#+3y�3t(v3FrN3�}3��3#d�3��3�^�2`�x3Vv�3��3��3H�v3%��3q� 3�E�3\��3N�O3���2�Y94�IJ3#X�3i.3 c3<�)3��3*�O3�M3*�3r+4j%�3D�3��35�P3]}3�3�G3���2�/m38�V3ho�3� �3�3(E�3��3_�M3>�3(�3�J�3�RW3�K�3"io3z�]3-�3�
�3$T�3;�3�L�3IX�3J��3D~g3�:�3]��3ڪ�3�a�3�5�3��3L��3O��3��
4Z�3�!�3��V3`M�3�R3r}�3c��3�p%3��37��3lg�35��3���2Y]=3=��3�i�33��3�%3���3�c3&��3K�a3�i`3׉q3a�3�3�k�3��?3�f�3.,w3?aM3v��3r�&3��3�j�3DT�3�"3/93T��3x3^�3�X�3�!%3\��3��l3
�3��3a�3�]�3��84�>13���3��3�n33���3�f3n4�3�6$3�>p3�s�3���3QU3���2�B�3�3)��3�3�DR3��3��3ƙ�32D%34>�36GV3;��3zeF3e,M3Z�\3��*3J�c3j��3�X�3�p3��[3�n4%�3Ie[3N� 3P�u3�3NU3S¦3�Z$3�&�3��3�ս3��3���3�0�3<��3�9�3
@Z3*ň3d��3Wڏ3Ԥ�3;e63?�,3��Z3�r�3���3583��=3���3���3��3��f3by63j�33���3ZMi3��13� V3�lM4��<3g��3��3�$�3n"�3߈3IC}3��3�3cK4�9�3��q3��Z3v�J3C��3K]3��w3pF3��b3L�33Ȉ3"4.3��3Ϲ#3�f�3��l3�DF3�l35$�3�\�3!N�3Ū 4k 3Ma�3!�3�S�3��3]>,3�W3D�3�!'3f��3༅3���3/�3�p�3�3�F�3'H63B�_4t�;3���3g��3�fc3>d53i�3�˥3 �K3��3��4���3�P�3�Z23O�S3�3��\3@�3~�3�f�3 z3>��3�	�3z
L3��2q��3�3y؂3�?93[�C3X<�3kЊ3n;�3T� 3���3�4 ~4`(�3k�3�3�=�3��k3��3hdM3s�3�m�3�ة35R�3�43t�35�3�<�2�:3U�2�̯2�53�'3�a#3T�3�3�v.3c��3���2�I�2��F3�H�29�2�l�2��2��2�M�2�Ax3���2�n3~m�2���3k�
3Kc 3��3{,_3�I�2�+3�r�2�e�2:	V3�F3�~�3A�3���2�Q 3QC�24�3b�2�W�2<D3{	35�U3p��2�X_3+��2^3���2�/�2g�
3��3#�2�[�2qQB3M�"3�$C32�3�h:3�,�2�܈2g�43+3ę�2�K�2�o�2':}3���2u�3<83��35��2��W3���2)O3j�H3Ma:3�3�!3�z3�l�2?��2�\�3�0y3|39��2:�3��3���2 �\3ݑ�2�"3e&3$q3���2��32�3jd�3� 2;
3�3�$'3�f�2�U$37y�2�þ2su3ue[3%�2�3!�2e=3B93���2��$3�J3�=3���2eW3
�3:��2��2%�3�3 �3��2�m�2�d�2$e�2w�#3a��2�8�2�d3�S*3.'�2{��2;03�P3�}3�W�2g 3�D3y��2&X'3i
3K�2��2gD�3Z.3$�3J%3�3x��2��;3��2��2�J3�j3��_3I�H3IY�2~�13��2��
3a53-��2��H3�Ŝ2�@3 W*32�2��2-i�3 �3ȳ�2Ï�2?/�2�'
3�n^3Ōg3^�2�Z`3Bf�3��]3��2$��2�F53��2[)�2Ey3}�2�� 3�k3j�j35H3{�2�L3?�n33v13E�T3
�E3� T3<�83��2��)3!��2<3��j3O�r3�j�2DͰ2eN3L3q�2b36v�2�V*3~7�2^L�3b%3��2��2�?T3~# 3x��2��2?53���2u�3��3g�2SZO3�oC3[�V3�V3v��2d�%3�\&3���2DC3��2ٶ,3a��2.h3z>*3�J�3}�F39a�3�9~3�N�3Ĭ[3���3n�V3o�o3H13}�E3
Ƌ3�&�3/�3�W�3��L3��3�K�3�xh3��Z3\��3�>V3�jC3��3�^_3��b3L*W3V�3� 3Uֲ3\>3B�34)3ǒ3:�b3cu�3WN{3,�3��}3J�k3�93"��3Ҙ�3���3�B3��T3#<�3�b39�3=[{3�<j3�	3^�3^u3�ɛ3��A3e`�3�C3��3��3W�3z��3B��3k��3�2��2A��3�3��
3Z��3U�U3���3�23�>�3�[3q��3*o�34�4��3�*p3�3L3�Ps3ŶU3O��3E�3��73i�3�V�3jDJ3��_3�y3���34(�3�23�3)�H3C/�3��3���3	�83�ݕ3�Č3�4,�I3�Y[3�Y3�c�3��Q3�3la�3��k3��3���3k��3C�U3��K3��3��>3H�2O�3�*Q3��3�p3��3�]3��3��3�w�3u�3��53k:�3�}4�c3�s3��3�V&3�bJ3Ũ�3���3O�a3�3�a�3��3Gx3��l3З�3��3��3�ӫ3UWm3��A3��3�84��_3�d3�[3~�e3:�!3?��3Z:F37�z3�k3�4�SF3Bl3��)3��g38�L3��s3�ү3�K3�}3I�G3�XU3��3�/�3L5(3H��3}J�3���3	`3��3�"3p�_3J��3OQ/3/�3�3�u3���3�u3�Ƹ3s"`3M^b3��p3�;�3jۏ3�L3#�4YU134��2��031P4֢v3�5)3��R3��v3��3��}3�3�*3*̓3]��3<�3�x@3�V3'��3��,3k3�`3�3��3ȫ]3��3
�o3�f3^�'3��4U�63h�k3��Q3>z3�.3�Y3"i3~�+3��3u�3�O�3��3��36�3�W3�F38��3��3tǿ3=_�3��3�&B3t�3��21��3��2�yM380�3�43e7�2 ��2v)3~3Z��3U�R3�F�2n�3 `�2��$3Z�03L�3�+�2qd3��3���2I�u3�� 3�3AG83��X3��3�u�2<�2��l36�2O(3�3�4�2�:@3e�l3x��3]�3�$�2�3��A3���2X�.3�3!5�2��d3�.3`�3��03t�3$�3g�
3��P3�c3�	3���2ڕ3Y�o3 �2?��3qK3<�73!�3Ӊ3A*�2��B3J��2�b3z��2j׆3��P3�gK3'J3{�3���2�3�Պ2ωH3%3f�38��2/�3	�\3�g�2|�3���3��33I��2ˍ�2Z�3Z�*3��2y8�2	�2���3c��2/O)3_z3�h3w��2��3��2�c3u�3��2î�2��3K�3���23^3'�g3Y13+!�2�`�2c�}3@��2���2�3-38T�2xF�2��<3s�3k%53�A�2\n3��2^(�2�M"3	8�2���2�3�3r�2�m:3WM�3c3���2�3�u�3�3Lh�2j ~3��2�'�2&K�2��38�3�73�J�2پ3O.:3��i3�e�2�sm3��3�Mj3'+3�pA3B�;3��35z�3��3C�&3v��3�G�3�� 3 �L3��2��3�}13�9=3׽@3)��2*��2.>?3�2��#3��3�C3��!3]*#3�A)3�V 3/x3�im3��B3�3�2z4*34�2���2�F�2Te�2�t3=��2�.G3G�2�H3�J3�`_3��3a�3��$3^=3\s�2�&3��=3�F�2�@3V�O3׻B3� 3��33b3���29B3v�3��L3�lF3&��2ah3
3�$�2!��2c��3��3tU3�F�2�e�2�l3�{C3���2�R�2�:3B��2�<�3\�&3H�2�"93�3f3��2Q �2�ܥ3N3?3�X33��u3��R3p��2Z)�3�;3�/
3֏3U�J3�|�2W�3���2��2�i�2Jq3�U3r��2��A3c�2:��2݈2�73�c�2#�3P��2�T3�|�2�3ʽ
3@N�3uOF3B:R30�;3+R?3�*�2ͧ3qI`3��3��/3̜�3�NR3��$3B�2��]3�%H3��B3�'3�4�2��'3��2��|3��3��2qX�2�[3
="3h6�2	b�2���2���2�s>3��l3��2(�H3&t�3�u�3�3'�2�v3[�#3�t�2Ā�2=\�2L83Z5�2"�C3]g3V�3%�2���3��2���2=b;3�B'3?�2��3`g33�K�2{X3�xQ3�83��;3�2�3�m3�j�2�2��2~܄3���2/z[3�3��2�-�2=��3��!3+� 3[� 3�Yd3�P3ߓ�3o3��2�.3iB�3qXG3��3Pe3�0P3�X3#$[2�ZY3��2+�P3���2Oy�3Ջj3ȫ33l�2o��3��-3�c�2���2�T_3��B3�83��N3�A�2�`�2��t3�{/3�D�2�B3Ȝ"3sH3���2a��3���2�|�3p 3���3�3h<�2 8
3p>�3�[`3O�3�EE3���2���2ZR3�c3���2�S3->3>[3u38��2t�2�
F3�2��3��3+O�2(J�2��+3�V3^?3�aq3��3ND38�2�)�2��$3B3�Es3�@3Rw�2j3:�3_9(35�?3�j2��M3е�3�3��@3��3�Kp3|
�2�d�3���2T2*3A�3�f�3s��2х�3�G'3���2�	3���2\�b3�|3��o3��93h�3�	,3̞�2�:3�[#3R�3J�23#��2��f3p��27w3PAM3��3r�13��3�2���2p�2���2�`�2Nq3�^G3�ؙ23�*3�,�3�D[3���2��2"=36�,3Č�2� U3u�3�3m�2323��3�ș3E�w3�e�3-�&3)(J3'!r3�M�3|�73��3��\3�eK3#��3b�3��Z3b��3�<43�=�3[��3r�o3�e�2C�O3ލ3�E�2߬3��3�2 3�=r3O�3o�3�(f3nNM3��]3c�3�W�3X7�3s�)3w�3���3"ت3���3�y)3���3,p3Qe3��}3�R"3=��3�-q3rö3L3Ȝ3�p3��4�&3A"~3G�R3��3�UJ3[�3�B�3�3l��33�23Z��3�F_3*�3x�3���3��$3x>�3��3��3��3~��3xP3�غ3^�f3;��3�23u@3]�@3��3��|3M�p3Ӎ�3u3��]3fU.4#�)37�'3M��2�?r3��23�G3��3�!"3|�3IT<3�ο3o�C3]�3z;3z�3d�3�n�3�\73��3)0 3���3Qa�3֝3�É3���3��3T�`3.�3ר�3�z3��3D/>3��
3�g�3�=3U؁3 �E3��%3��Y3��3M�C3}{�3�3�ɝ3�Lh3c�#3�Fk3�f)3`K�3�3X�3�i@3�I3]�3zP�3z3��3�p3�<�323ݮ�3�u�3��>3N�<3���3�y3��f3�̍3�'3F��3ī�3�np3�e�3�w�3M4ψ�3sP\3L"3Aܠ3Z 3�S33�~U3�\,34Ad3�BE3�X�3�U39��3@43�4V	3ÊI3*�39��2�NR3Z3��3��Y3��?3���3Q��3ق�3j.i3%H3�˝36 �2��M3��z3��[3�H03���3}f-33Ϛ�2P��3w�E3vq3�
&3��u3w=3~�t3�I�3I/3��H3�G�3*�]3j�3!3Hz3;d&3LE�3�݀3��D3��A3��2���3\�H3n��2!�28[3��"3�\63��93x5/3
�3�Cr3ĉ|3B3�h3�<�3e�3ڻ�3���2L�3��S3��43���33��a38s
3��3�03�qU3�H3HO=3�3j�Q3~ 3�83A��2W�F3�R3�y13�*3vԜ3M}3CX.3?c�2w�:3��R3&�3c435c�3�Ѓ3�� 3��3�qc3�	3�I3G��3k3�=3�uB3�bL3�a3�33�t3�Oj3!C3X�q3N�l3���3���2�9�3=�!3���2sـ32�!3TSC3DX3�[�3[�D3�K\3UG�2]��3-OV33�2L�T3��;3�2
F3?Rv3���2 �'3��3!j3<{U3�-�2�F3!v}3�_3�93�]�2��)3�E�2]#3}*23o �3�33�-�3[�3%�h3X~/3e�13ZD43߸3}�3���2��2L�3�N3��O3Wv�2��O3��a3���2�$]3�23�W�3��3$={3�S3163^n3��]3�-f3���2$�C3�ww3AZ�3��3�PY3��3ї3�1�3	U3�53&�X3�X?3�]38�3���3�8m3m&(3��2�4s3��_3^�M3�
m3ND�3HB
3j�53���3V�P3㽇3?a3`K3W�23 �3���3W3E3(¢3���2��3W6]3���2X�.3�}3E�q3�;3%�D3D��2ܺ�2���2i�+4��,3��D3GT3�?V3ĵD3���3S�O3�*3�*�3u��3u�R3xd�2}��2��#3y33�k>3�C�3��2�F�3<3/8�3u�3>ay3*9�2�q�3�03�=3�&�2���2<��2�/P3��T3oդ2ayG3?W73��3^�q39z73�M�3�Z 3��'3�43C' 3�K3�2�cl3|��3R�&3�;�2aT4w��27S3r4r3��K3�j%3��53C3V��2���37�s3�L3��3C9�2U�3-X3�	'33�2P�k3ҍ;3v��3��<3	Z,3n��2���3K�2$�3
��2�>3��13�-3^7m3���2��3�U�3�H�3�&�2s�	3���3�W3��3Ӧ�3��83�U3�|3�<�3K)3�T�3�H3-��3��3,~3V��3��33,\3WC{3�.B3���3n�4�v3�p3�83��3ТT3���3�(E3t�32�d3�3c3�:�3��3VZ�3�3�	4�w3�]63`i3���3@E3֜�3���3�Sc3?@3Oݻ3�)~3^k3��)3� s3�c3e#�3g�p3��z3���3�^�2�.�3x��3�L3�6~3Իc3t:�3Y�L3=3���3��j3Ҝr3[�3��3[��2�;�3${g3� a3��N3k�3��l3�3P\�3��!3��3�6�3$ȿ3<B�3��3۔3�j�3;?43k�\3Pu�3U�3��3��c3��x3�3��A3{�3E�3yPR3Ā3Mh�3��33�#3��3�Y3�Ы3�43U�U3!!�3J3�L63K�4�
U3Wg3r2N3qe�3��[3��3���3e(3ڇ3ݗ�3�Ω3�~Z3x3_3��q3iB83�_36�W3a֬3y�3+�3(й3%H,3�VZ3��3�b53d��3���3�3�RN3e��3ɗ�3([�2�3�B�3�Ф3��83t!3s��3o�3LrI36u�3S�3���3�b39�3�33�"�3��)3�g�3�dl3�@~30p3�qr3�b3b�3���3vM3�XQ3��3���3W�w3��2Tڃ3k�3ʖ!3WSO3��z3�K�33'3ƶ�3�V38�d3�23{��3�L`3H!k3��3�ۇ3ma3�O3�U3�b)3v�3�z�3�֧3WST3�>23�J�3��3�53� �3��L3�y3��H3��4��M3�H�3#2`3��Y4	��3���3��3-Rx3�U�3�)53�.�34.3���3�o4��3�|�3�A3�w�3�3˷=3'w3�>;3��3
03W��3�?3��A363;4f�-31K%3
�v31�L3V�3Y3\��3�2u�3�4�}�3��T3�;3-�47a�3�v*3�<�3��n3;3'J(3y��3I��3��3��3ΜF4�cd3yF�3t�3��3�+D3P��3�u�32��3��3��4�@�3ڠ�3!r3r��3�"_3��t3v��3��3L��3�73���3���3Ď�3��3�Y4��3�B�36Q3v -3���3�m�3p��3Ps�3]3�'*4�X�3,3WJ53�M�3x�3�s3��30cL3��3�Y13��3�g�3��3��W3a64��3� �3�&q3/�a3J�3d�h3!v�3S 93��f3vU�3���3a�3!�3l��3�9�3�	e3�"�3��W30�3��30
�3C)�3V��3���3[-648L]3Pˠ3W�f3b�
3�3��3\�3%W3���3�#�4��3X�l3�n'3K�3gPc3�`+3��3�ډ3���3��#3��3�J�3ь3KH�3��K4�<�3�y�3���3Q��3Bl�3��3�R�3��R3�v<3i64c�3X$�3�j]3��3h,�31��3���3$�<3>p�3�:3��3��3�q�38.�3�7%4:.�3�K�3��k3ݯ�3�03F��3��3�,�2H��3���3���3ɢ3!UQ3���3�%�3`X@3�&q3`>3��3��t3J�3��3GiB3.�o3��64�"p3�n�3���3��g3���3��3i`�3��w3�q3�R4�.�3R�c3��3���3D��3�Ż3.ă3+oG3��{3Y�39b�3���3��R3�b�3��*4#�3�"�3
r�3��A3&�3�3��4gr�3x�3��4�	4�Y?3�.93c�3�7�3��3�4�#F3i�3ꢫ3�� 4!�3�:3�L3!.c4���3%�u3}��3�=\3:��3�\o3�}�3�d3���3ۡ�3���3!��3y�'3��3���3�H�3���3��X3Pz�3cY�3x4� �3hZ3��3k44p#(3��3(43(^3l63�Ȗ3}o�3r�;3˾3��3[��3L�3�
3���3Mܐ3���3g�3��M3F��3���3��3v��3m�4f�3�?/4�=�3V��3���3a:�3A��3C_4���3��3��3�]:4�!4֨�3���3���3�L�3��3V��3�$4��3�(�3Za48:	4��3���3��M4	*�3�b�3���3H��3�Ũ3�0�3���3/%�3 ��3�� 4]Z.4��	4׍3Z�&4U?�3���3[� 4O�3��3��4׍ 44 4X34���3�Y4�G�3�#4Q��3j�3�2�3B�3l�/4�P�3 
�3�vH4�(�3�ٗ3VW�3-�!4�v�3�d�3��3�X�3��4Έ�3�V�3���3uɳ3�J�3�9�4�+]3"c�3�Y4B4�3��3�D�3�#�3$f4��4?�4�\�3黃3S�3��4g�x3��4�54%��3���3h�
4�_�3\��3[?�3{q4�.4�,�3k��3IM�3R1�3A�4A�4��X3og�3I�R4v��3�X 4ڷ3G]L4~64o��3���3s:{3UH�3xi�3��4�_+4Y��3��3}�34�/4��3H�3e��3��3j�3��4't3�^�34A%4��3h�)4�P�3I3�3w�44仌3���3G��3#��3qu�3���3��3pM�3��3L�#4�<�3D�	4���3;4=%�3k4�9�3"��32Pn3�o�4�L
4h�4��3���3��3]�3i 4Z04S��3��3�g4��|3�Ǣ3R��3x]G4�՟3��4�e�3�3�Ǆ3���3�d4���3}4�I�4�4�t�3y&�3�*�3�$!4э3�!�3,��3�פ3��3�y�4���3���3q�3,̕4j�4r��3�{T4o�39��3�Ϛ3X�	4I,�3���3�Y4��4��4)�3V6�3��^4j4[q�3�۶3d>4bg�3�H"4,D�3"��3lB3�֘4�ը3l]�3���3�D4K6q3}{�3T� 4B��3vy44��4��3��3�3�74��3�/�3w7�3���34���3$mV4[��3��A3�T�2g�3:�3�K3��3�w3�c�2W:3��&3�:E3C�3��3��_3s�3�s�2eQV3	)A3?��2AC�2.?3�]3S��2�
3��3�j53��3�1�3v�3�(3�3993!��2�o�2��.3|�2E��29��3WH!3�-�2�ߌ2��3A'93773�q73S|�22I3ν3�	3�3�?3�J*3;��3�n#3��73��3�)3w%3R1�2�2Ă�2�a3Fq�3�}`3}�$3��2i�
3�j�2퉹2��03!3^�S3YF)3�53��e39,�3u>3Pz�3cb�2�y�2 Q3� 3_0P3%��2�f3Q��2gG3dh�3�p�3̖�2Qv�2��/3m�J3sM�2��M38��2�@�3���2��3�� 3�3��2�ؖ3�"3N��2�3�S�2WR�2�t"3jr3�43$HB3�F�3�[3��U3�>�2S��2M33L��2�3��3�L3�%�2,F3m�3c�2,��2I��3��2l '38�N3�Q3X�2��3?�O3	ȑ2���2�"z3
�?3Fl83b��2rr=3�!V3��3�}P3�~"39�'33��26,�2(3�$3���2���33���2j�93Տ�2��I3+��2:�3�3C�3���34ig3i��2Ս�2�R3�t3���23-3Lo
3��2C�2@��3�C�2�|�2s-3�U�3d�3�o"3��3��3'��2Ea�2+`�2��2R��2Uߑ3��"3Kq#34�2͟!3�F3���2{30>3�Y�3m'�26c63�83��G3S��2�ߡ3)H3��W3`�T34#3�#3���22�3�T	3FSa3�<�3*�<3&$3��2��*39(36(i3_��2%��2+T3���2�!3"hi3�p�2ݦ�2�B3@'3�9�2�)3T�3*3(y 3�36�2��3��3��V3���2���2-u3�r�2WD�2p&�3���2
N3-��2[r�33@3��3�)3#��3��
3�@�3y	D3��3O\3Z�x3[�&3o�36�_3?��3i?�3i�g3��3��V3�g3i�2��3r�3��d3�W36��3�Е3\�`3�>�3۟�3Y��3f3a~�38W�3��a3'�3��3!2)3	��3R_G3�7p3~�3��j3Pq�3�b>3�@B32u3�l3���3��=3��3~�`3�mN3I�'3.4$8I3�d�3aS:3z�_3��A3&�K3�v�3<z�26�R3. 42U�3 �I3J�:3�]3��3��3��N3�&d3���3Z��25>]3�˶3�Gl3(,j3l	I4<~3e�L3�}�3�dc3RN3�@G3Q��3��3�u=37(�3���3�Nx3t�3ssf3܊�3�r3��N3�GE3��3r�36��3���3��G3��3ý
4�:36�3�;3���3~b3TV�3H�m3�]*3! f3�3��}3��3S\3E�3�\3�~Z3fSx3-9s3�f3׊"3�ߑ3��3�<�3��3���3�ӥ3᰷3�4�3�pk3�3�j3���3m�3x�73K��3���3P�3,3׌3T��3��2���3��-3��m3�z3�W�3h��3oE\3�3
a(45:�3n�3@�S3-G�3>B[3K�l3�ݗ3�m*3|�3�|4L[�3�I3�3�1�3�$�3e�A3B��3��3
z�3!�35�3b��3!m3�E&3���3�_U3:Vw3�f�3W�93���2�R�3c`o3h�3�	�3l��3,L�3x�'3��3E�U3L�K3D�R3�x�3ƢC3 \�3�x�3��3�~73��<3�_73��*4Sg3�P3�8y3qY3>e33"�3�(�30�3���3x�3�ώ3��3�B3�3`�`3J��3U�C3Y��3%��3
83)��3�ě3U�-3�l�2��4��e3+��3\W"3�3i`C3�k�2-��3O73B3�3^��3��3��Q3Cz3:Դ3	��3,�3�im3!-�2f��3T;.3p��3�<]3M��3Ԏ*3%+�3`��2p�33L�A3�B�2���2�ɗ3|�3/�T3�>3@��3�y63���3\{ 306�3/~3x��2���2xgV3	�3>� 3���3J�'3�Js3O�V3�3T��3-ښ3�63�G*3�j3I��3V)s3V3�r3��3���3�Y�3.5�2�q�3c&3Z�2�3J3�/.3��3�[^3� �3l$3^Ld3ڞD3U��3�3��3���3�83�2'3u3jY�3�B�2J��3�k4:O3��F3S38�Y3��13���2D�@3��3�h�3�G�3��3h&D3ʔ(3u�*3U��3(U3KC3�[3��3��+3��n316�3_E3S_3���3�f^3e�-3��"3��3�R3*M�2�+3��3R�3�'3��3kM3�!g3��3��43ge_3
�93�h3��3�>�3y�;3��
3o�g3j�3�$G3���27�)37y3l��2�'�2�&w3"��2�x3��53���3�.B3Ӷ%3<03�q�3,��2xQ3�'3�{3��-3�3K�p3�x3��U3�~�3��3~(i3�3�6d3S�3�)Z3�ws3@�3��)3tU�2��3�hK3 3]^3��30�&3-3�w!30MT3l}I333�!B3�Z3��^3���3q?�3.�/3���2�s�3^\3;3� b3A�M3��+3��2�3E��2L!q3ѹ�2��4�%C3��`3�i3�h{3yJ83��J3���3�3�A3!�3�7�3#��3�33� d38�^3e� 3g��3�"�2� �3�033�w3�j3�*�2G�83�u�3N3�HM33)�36gF3GpW3�
3ʩH3-3̓�3ຩ3̫�3�w3yG�2�Ѐ3�U�3t3�V23��2�zZ3��3q<�3|�135��2�V3���3��Y3Z�Y3c'3�;c3ӆK3߀c3(Ȗ3"!3�3���3�Xd3��x3�8&3�O)3�MY3��3�ױ3�;3�*3�}3N%4��k3�4Gw3Q *4,w�3S4�1�3�s�34 �3g��3�3�q3$�3kZ
4���3 4���3� (4p7�3�4|3G�3L��3�4��?3��4�C�3�`�3���3��m4�n�31`�3�1�3K�3e��3�Y�3�X#4�v3��3AH4Ï�3�k�3���3�I�3��3�t�3mH�3�Tv3ܹ3��35!4��'4�h4���3�4S+�3���3Gs�3���3�e83x�3�4�d(3ћ�3��74L��3�3�CK3�54�.�3�ǿ3i��3nL�3�}$4]�3�4_cl3`��3~?�3/%j4Ō�3���3��3���3ǿ 4���3 �4�x3%�3�8G4���3«�3�xm3oݵ3�г3K��3*��3��3�U.4���3�0�3�2�3�h�3���3��[4R��3"L�3��3v�3��{3�e4Bڧ3�Y�3���3x&-4��3��3�=3 
4��4 AK3^i�3��3xE�3��3 64���3�9�3`�K3��/4�f�3r��3��3aڣ3�4�3qi�3Ǵ�3	�3���3�m�3y�"4�V4i�c34Z&4yZ�3��4��3��04Ō�3d9�32j�32}�3$Q@3�(F4H�4�&�3en�3�O�3�k3���3Я74���3ٷ�3A�D4��4�#�3�Q�3��4`��3O�3�w�30�L3W�3�v3�j�3U��3�Z�37 �32s,4��3@�h3�:�3/��3h5�3��3F��3��3M�4OA4|�3�<�3���3���3?��3m��3Qq�3�;3��38�{3��302 45�I3,f�3�414-o�3��3q�3�h3Ug3��3H�Q3��w3dr4�X4$g�3�2�3<�37��3]n�3�	�3Zc4
BO3�3�X3J�.4�R�3��3���3\.O4���3��3���3��
4�F�3^l�3��3�v3��3_@=4_��3.��3E:&3�I�3,!�3/*3 A�3�h&3���3�c�3A�35�3��3�:�3Y��3>^3�5J3dz^3�ր3���2-�N3_�3P3�T<3k�3�HY3�m�3
.H3�q3b��3c��2(*�2SD3�=3<n�2fT�3۠�2,F3g(.3J:V3�(3��3H&&3�s3�$$3�^{373��	3�`3���3�Ǳ3 3e 3{m*37w;3�&�2�(34��2v%3��3�g�3��&3}a�2	�<3y�3��3�*`3��>33��3�>3�]�3��^3G53T_3�v4�3�r{3���2��L3bP3F{�2��f3�f3��03�W 3\��3��e3�'U3�3w;�3A}E3�X?3֯!3�:V3l33^��2�{v3n�3�}-3��z3��3��3��/3��3濄3�,13��m3u�3}w�3�v!32D�3�tD3�2e63i*�3�*3.>E3\&3$�W3e�M3��3>�43�=3�13���3��j32�]3���2 G3��3�!�3�^3-r�2w�k3�f�2�@y3�d3)(I3͎{3�ޏ3���2q�V3�V3��3L�3s�3/ʂ3��3��3��3��j33�I3��J3D��3�3rQ39*W3�,�2G03�Me3'}3��K3���20��2gI�3��3��3��/3#��2�Wj3�;3�C3WB363_)93�E3ua�2r�?3�%�3WvC3�3[I>3+��2��3?�<3�rk3��3SQ3�%3�Ԩ3�3y�_3�3��3��3�1E3�83�q�2�D�3 S�3H�3�ې3l��2� L3oH3��3��^3�C)3�[b3�w�2e�3�M3��3U��2 #�31w23�?.3a[[3Ď@3lL3X6R3��g3�)�2+V@3:ˎ3�HV3�a�3��3Έ3��3��(3�^>3M�3�S3l��2�х3\��20�2���2�[�3F�3\�3L�"3y� 38�2833��O3��3vx�3?��3�!}3��3��2�3+��2wF�2�|S3`� 3��R3@�2��3x��2���3+>!3���3�13�ߦ3�X3���3���2� _3Cp3o,3��V3&��3o3N�73*r3�L4�NN3�3u�E3_3���3��F3���3�%�3�K�3T3n��3�.3��3�9�3	��3�%3I�:3���3Ƴ�3��3f\�31�3 2�3wP3+4y8t3'+�3��3HB83G��37F3�4U�s3%`�3��3D�4�w!3eN;3�9�3�Ҟ3��2�x3[±3��,3�ʹ3��3"u�3DAB3eZ�2��L3�3��(3�_�3vO3N��3�J3J��3��b3�]b3Z�13��04W�z3���3>Ҫ3�O�3\:3CX�3�3�zG3��3�V�3K��3��3�p3��k3R�3/4%3?ZY3��T3���3=��2Nڞ3-�c3ˉK3�F^3؋ 4�w3
U�3J�h3%	M3�N�3��3���3i
 33��3��3fx�3E3ȣ�3>M3)�l3o<�3��2��3ub3F��3ʛ�3K�3�$T3.��3� �3�SA3�T�3�0�3!�^3���3��3�l>3t�l3�/4"�3䂍3��3�z39��3�33ٽ�3@�w3�6i33�3�ۦ3P&3��3�v3.4i�3S3���3@�(3I�3n�W3Ө?3�E73=�S3���3e
�3��W3�K3�B4��3��z3��3w�3��3��/3U�3�VU3��3�[3p/�3��Z3+�D3�P�3�F38�m3G��3*+�3��363m3[��3���3rx�3��P3�4�3Ʀ�3�c3��3�*/3i3��Z3|�3�EU31�3h�33=4o�3�8�3i3�3��37�l3"J|3}�3�l�3ރ�3lz�3���3�ǈ3Q��3�T53��B3���3��3��3��3��x3�0~3�Č3��2�;3�E4|�3��?3�D�3���3�1=3.�K34;�3�Tp3L	�3�Z4��3��[3�R73%$�3��3)�\3�3��t3�]3äI3��$42	n3#M3�/�24L3畑2��3J҂2���2)�2	13I��2���2Z\�2d�^3 ��2�z�2�Y�2�.3�P�2ȝ�2W��2г�2f3gy�2�513`��2�h�2�	3bJ�3
g39}�2'�3E�)3}U�2��2t}�2nJ�2�2�2��z3(<73�E	3��2D&03s43f~�2g�%3���2H&3�C�2r[\3<<G3i �2�G�2�7P3
��22k�2u�L3V��2A�2��2t�	3.�31tj3J�V3��3 Q�2B#�2C�V3�8�2J�2u�3�s�2�\�2?�t25}83���2d3�?!3Um|3�r3�j�2�b�2>�3���2��3�H�2�w�2r�3�D3��?3�x�2{^�2��2� 3ڵ3K~�2S3�u�2�n3V�<3@h�2���2��3<(�3J �2a|3+]3��2մ3�i
3 _3���2�:3���3"#3 �3�gt2�(�2 e3͙�2{�y3�ߩ2�3� 3��@3CW�2jX�2�{�2lJ3��2�3�+3C��2+��2��X3xq73��2��
3��f3��53�q34�2X�3Usc3E0	3�d3�r�2�? 3��33���2e� 3�3�>�3h��2���2�ر2>>3��2_zV3�3'��2g7W3@��36�3��3{@�2��3?-�2�_�2l�3��2ҟ3�393_��2�a�2���2aP�3�X�2@�2N�3�A�2�43��43��O3�?�2.�3��[36�,3w��2���2�q3��2::�2 �3�}�2G�3��3�]K3a!35a�2���2��3Y'3�*3p�3>��2�&�2��3[3H��2��	3��d3��3kE3|:�2S��2x��3��2u�3§�2}r3���2�x3�Q�2�F�26OR2f̚3�F�2
83)7�2�\�2o3-��2�F3��02 h3�r>3�3Q��2j��2[D�2`��2H�z2p��2�y2y+N3j�2�GV3 �2t��3�k3�7�3Hc|3�P	34~:3jY�3�03�T�3��3��f3�Nk3���3͊�3ko53�M3⯫3�e�3g%23�3�2}3l5�3��3�t�3,�3sr3�=3N��3�/3>l�3~ʍ3��k3�r�3i��3=��3.i+3�3յ�3\��33��3O�3��r3��s3 S23]?3F�3�D�3;�3]g�3��3}�F3
�F3�g�3$ C3�YD323+�j3�=:3~�^3�:3L�3o(�3lM4���3{�M39��2A��3I�}3�A3[��3P�v3N�$3�d"3�R�3�r�3�6�31�3�b4H�_3 �j35��3�X%3��f3p�37L�3�]23�DR3:ҷ3�4m�03I;3O}=3|�j3�z�3�ׅ3+3�!b3�/�3���3�b533�'3�}3�T�3�?3d�]3>�3��3�Q3٩3T�N3;)3
?�3�)�3n4�/E3ʵ33��3�:3}t.3㠂3�#A3��3~�r3�03;��3�\�3��>3��(4r�3��Z3Q�3��y30?3ڠ733��3�3��3�x4V��3r��3X3vc�3}[�3Mn�3��|3��?3wIc3*�93�t�3�`s3i�w3tF�2��3:�3G��3a#b3A/3S�M3�J�3j��3�,,3�ε3A�4F.�3�Ep37��2�o3�)3�MY3 �]3��3���3�9S3|l4�u'3!g93*h3?�4A�L3�]�3�͌3��3��A3/۔3���3a��2�,31�4
�3��3��3&��3���3�93L,!3};�3�A�3͎C3f��3���3��Y3Hț3�p	4�*03�ˁ3��u3�\M3Δm3;)3:��3al3<P�3���3��3"g�3]p�2��3�_p3l1�3"�]3ǋ�29�D3�Z3�r�3�#3�B3LE3�4�MF3���3�zc3h��3y�p37�<3��h3��$3�O�3
��3��4�A�3��3�R3�a4�B3���3!q3�:�3�M3��}3��C3o��3^�P3�į3��;3�k3TBx3�33m�{3��`3��T3��]3k�3p
�3Z��3w�3���3�z3�t�2Q~	3�3Xno3��2ݝ3t��3++�3v�\3��3d�	37\;3�:}3��3[c23[څ39��3��3��N3��3���3`݀3�U3�3I��3ϱa3f3�73��=3�V3+"|3AdX3*13��?34�93�xz3c�\3��G33�3G�D3���3LKW3��V3t�4	P^3��3�3TH83��3��13�qT3��S3��3|�y3�э3f�U3�Y3��3��4�U3�f3��o3"�3�u3X�3"��3(�o3�G�3_4@��3��3��3�q�3�ku37~ 3Q}23��3:m�3�`�2[��3a�$3�3��,3�(4�63hbp3�3_��3�3�{36�3�h+3�M�3�Ә3׶�3�lU3W3G-�3���3'3?2�3yd3���3Y�.3�l3s'/3[\33p�3���3
o3��3�h�2�=�3�Y3��f3�t3��'3�*3�4�3T�3B�3�3,߷3�ri3=53<�3���2�\�3�!�3E3��Z3c!^3��3���3�E3��t3��93��M3]3�>3WR3�f3�yR3p�4X(�3��,3q��2}�o3kF3iA3b�T3�,3��`3��93*ns3��03�
(3�U3��3�,3G��3��H3h�h3�@3Ei3Z׉3��3�?3�s3��3���3��#3ي�3/d3�23̖Q3��(3α�3>�3��3�{3�53��_3�]�3r9V3�f3d�[38�V3}3j�3X;�3E�3M�g3���3-�13I|e3#�3^30b�3�@O3J3Ua�2n��3�;3E@�3R�c3<��2��2ӆ4v�3Bi3��3đA3� 3(f23
�3�T�2�ԣ3�0�3a&�3�Ė3;a3�k�3��3d953ˉ53�)3�Em3�'3���34^�3�[3͇A3S�3�K73>�-34�3�� 3/u#3���3�v3�03��3�[�3�n3�I'3��!3�.�3~{]3��2I�^3 �!3�\z3B�3|*�3XG<3!r3� �2��3��6323Fby3���2ߍ*3��n3�4B33,3�)+3M��3�oC35�.3��2�yp3	mk3s2�2m3�
3���3��!3I�3/X\3A�G3��3�-w3�3�%�2�53�m�2L�33��2��83Xt3�UY3~��3�=�3GT3���2�r�3���2<�2Bq63��;3F][3�3��J3#�33۴l3�J�3�#3��23Z7\3�kR3��[3�U3�#)3�}�2�.3�,�3��K3��2���2�J�3�o)3�3�ܭ3��3��3+��2I\[3�t\3�3���2ܼ�3�\3L�$3F�3:�53gd3�P;3���3n(�2=^Z32B3OM�3+�l3�3M�O3�&3C��2YY3_�2!�Z3Jx3O��3�3cj3Ͼ)3/��3[�3`�>3��o3u�!3�)O3�$3'3�3�?�2!*m3�1�32_�3u-03�M#3��)3P�U3R�G3K33Һ�2ƴp3�Z'3S9O3�T03���2
D�2��4U�30P3}�(3�K3�m�2��13�53�&<3齟3I��3��B3` 39v�2y��2��%3�O)3Me 3$k3���2��2��3�R3	AY3cI3�b�3�QX3k�.3�E�36�L3x�03+�|3"q73 1�2p,3(b�3$|53}�:3y.3�tu3�tK3��2<3�3G�:3���2]�3
Z33�2^H3��3�83��<3�]'3	t3��Y3I,a3x�35��2��D3�cn3�:�3OB�38Ϥ2�OJ3w�3��3	h13�23'5�3�,3"��3��+35�2�m3���3=3>^�3���2��2�13��3Z�C3bO@3�S�3=�3��3v{j3,��2�Iy3�3�|?3�@3&3*C3N\*3i�3z�3{��3��3*�4sǝ3Y�3se`3N�3�8�3��3��[3�d3l�3��3���3]�3)�K3���3|�3�=3��3;<�37/�3��3a-�3�M�3z��3И�3�$4�̣3��3UW�3Ԣ3�yr3/�4��3Z��3���3H��3���3��4-�G3�r47M3�F�3���3sE�3b��3G��3�4
�3��3y2e3��P4*uL3�,�3�m�3�m�35�3�3u��3`7�3!�3�:48��3���3��v3�R�3���3� $3�J3�Ж3���3��~3�^�3A�3u۪3�%�3>~24@��3�k�3�g3{+4`IN3��3^��3��c3Rw�3��4�$�3n"K3w/l33��3t�3g��3N�3Tf�3QL�3���3f��3�f�3R�3Ђ>3͊4��3���3seg3Jr3�m3���3K�3`�L3`��3k� 4sE�3?;�3e�c3\,�3��3�)F3v��3��a3��3�un3�O�3?\�3�{[3P�3s14=%�30�W3��+36�3���3�H�3M�J3��3���34�x3�0�3튕3��A31$4���3<�3�3�?_3�F�3*�3~�3�:c3�|b3Xy�3L�=46W�3w�3��3M�3��3ܞ�3l��3��l3� �3�n�3��3aQ�3�P�3«3뛭3d�~3��3Ot�3U�3�Q3V�3�O�3>-�3�~�3��_4�q�3!�3�x3��3�n�3��3���3�,3�3vl44Ա�3Mb~34�?3��3=:�3(e�3���3j��3A1�3�d�3��3�=x3*ɉ3�S�3���4�r�30w�3��3o��3��3�Ur3�1�3�A{3�X�3w-�3,�4A��3�<U3�7�3��3b��3:��3~c�3�6�3%��2��3� }3�0t3j3���3�W]3Ћ3�O�3�C3�Zh3�N3���3��M3��3�z-4}��3e�3��	3���3{.�3��3O�3|s3��3�'P3�24x̿3�΋3C��2�LS3�3A�t3�f3%v38y3��:3��t3��.3i\3̏�3Uɀ3T A3/�Z3���3y%D3р31�3�i/3掗3�93��3�z3��3��U3%j�38v;3~x<3�/3��!3A3���3��3��3!9q3g�3$��3�(V3��3���34�i3��V3��!3P�2��m33���3�~31X3lP3�w3:�3h֤3��23X�X3�1�2�J3�W3,�3k�u3U�3O/�3�/3���2���3��k3v13�3W3�3J3p 3Ft~3V�.3�C3SA3���3`�39ܸ2��23-�I31GE3(�3�F�3vo%3�83v�3@��3�F%3��2/��3�3��i3��#3m'/3Y3	;o3�c3�%G3y�*3��T3��3g�D3��.3��Y3�c3��3���3I0�3���2��3�f�3c�3m3*n�2�*e3HIL3��J3�V�3��2d�3L�43�O�3[5u3'�53kl�38o	4׃]3z5l3�3*$�3�	31�s3!�K3.��2��Y3��3���3�pY3�S"3>�3��3�� 32Ə3�)�3���3rk}3&o3�h3�Wu3�n3Y��3�M3k��3�U�3M�]3ԩ63�B�3��u3�1 3��63/G�3v �3I�<3�33� �3�i83?x3�k�3I.�2Li�3�l3Ї�3I�D3rBj3 '3"S�3�,53�'�2?�03Wu�3^2;3�j3�`�3*�3-�3�V�3O�V3t�Y3jy�2�J3��]3��)3��R3�+�2��3Mvq3ZΙ3Ǫ3�p3r#3�N"4�(3��=3,V73��I3�,3s��3	�3'��2;��38�3��N3�F�3n��2�R3���3<Op3��|3A_3���3��3�E�3LO'3*.�2� 3��"4sZ3�83� 3z3� 3D`@3��B3>3�Q�3���3��4�6b3�m�2�3���3��13x_�3��2��3]x83��3m��3F�3���3Y��3�Q3:�w3/�3�}46�|3�j36,Y3ðk3!��3��3�٥3��4Ƙc3���3q|`3�MA3��3DII3�u�3-f3X
3p�Q3@��3#��2��:3�3M,X3ទ3!$�3J�2���3�2�3Ȑu3�,�3�Ŭ3�4�3D��3��83��3:A3��}3FT93d(+3�^m3.3c��3�݃3_�E3��G3��M4,�73��3�X3A�|3�^�2�3���3��3;� 3�(�3_n3�_�39C�2:�/3<�3v�2�^�3�=A3Z �3�:G3	��35�3�A�3��W3���3�:3�Cr3f�G3�H3M7�3刄3���3��3H�M3.��3�Ʀ3\��3�3�+�3��_3R&3�d3X�3+�3��t3�.�3G�3;�Q3w 3[HF4|b3#J3z73�'3��^3L�3�w3	=F3�%j3|ws3��O3��3f
3��3"ʏ3;�|3�Ō3�13J�'3.�X3oڗ3Q8-3�w.3�m3`Y�3��3��\3,^\37�3��3Y��3�=Q3�i`3�bA3�b�3tz�3�Yt3� 3�3�}3��R3� �32��2E�3�.3Ѽ�3���3z�j3$43wX�3�'3�o3@]n3`-3��3M��3�ı3�`3�mY3Ҷ3֒�3��C3d�3mG�3`�W3�D3��3��3��\3)G35�3�p!3[L
3�/3�L�3��3cm3��V3G�3��f3,3f~3/s,3���3�S4=�3�W3n��2"v�3Q&�3��l3f�T3��k3���3�PI3f4Χ�3H3i53ߌ�3���2��3܇�3A�n3�$3%I�3��3o�W3�}3 
4K�r3
y\3co3�a3�NG3l�3���3�-3\��3>T03lx�3��3f�(3��2(((4��!3�EC3]�>3~�u3o83\�3��^3�~3�GA3���3*w3W�M35v�2��q3ZlF34�;3��l3��"3��3�3+�3�30��3��3h�84s��3�S=3m�3wC�3�.�3���3�1�3?u�3�r�3т�3�տ3-|�3�h�3�L 4�y3�D3'y�3;��3��3��3�443�3�z�3OU�3d� 4bi3(�3L˒3nʒ3�G{3_��3�3\*h3�]�3��4�j�3<u�3���3��3@,�32��3��3O�3�Y�3��3�C�3���3;��3F`�3X�4��3&��3OK�3�"�3��3���3�^�3�Eq3k=�3^f4�}�3]��3
�3��3�p�3�i3D4�33W\3�1�3�/-3�3��3Ù�3R��3�s4��o3T
�3VZ3��3��3a��3�J�3��23���3�3���3+��39y/3z>�3�|�3%)3&��3þH3���3��w3w�3S�w3�x3Ӣ3��4��3�(S3�.4݂�3y~32r�3#|�3�G3uq�3�G4�4gU[3�1:3��33�s3�`38H#4;Q3���3$Q3*� 4Mͅ3 i�3ܨ�3lF�4��3��3�m3,4��3��3���3e�^3/��3J'4�+4K�39��3�q�3S$�3�{3
V�3(q3P�3�$3L4<��3���3�o.3��B4}��3�M�3:c3��i3���3:y�3N�3�*#3L��3���3��3��3���3k��3UXb3�43ķ�3�3�Q04Ԯ�3�׬3݆�3f`�3>V�3"&4��3³3q�E3H*�3��w3Gی3�{�3Uh3G��3���3+$�3v�38O3���3sk�3�
�3���3�`b3��4/�3��4*<�3l?3`��3�)94�A�3��3�o�3�M�3�{t3���3�3��i3���3��3_�4h��3i��3�3��3�m38��3�1D3��3.f�3�]�3�;~393��3y�44LE3�S�3�)3��X3�\}3+��3�3�3���3�o�3W!4��3w«3�Iy3�3���3�3.̯3��:3�4$n�3�k�3�0�3"p�3�K3*�&41&B3�I�3Aœ3�Bw3��:3�Y�3 �s3��3Ͱ�3�3���3Ⱦ�3:i23O�4Ǖ�3��M3��\3ӧ3���3O�k3��4��3��3�X�3pq349�3��3�D�3�>�3��}3���3�d�3{�34Sm46�3D�	4��b3%ڍ3��3~�n3�S�3�ч33��3i�z3cO�3s��3w3�W 3�;4!֍3�_�3���3��g3���3�j�3=�3�i"3�4�3Y�4$��3�`�3�v/3���3 �3��13�4>�J3��3��3HO�3��3m��3x�3��(4Á3�N3��3!��3���3��3��3˭3r�3B4a?�3��3d*l3W�l3#5t3�T3a�3F3�b4�323��3�2�3�6�3�Q3aq4=B[3G��3�3�Xj3&W34�3o�3B�30�3*d�3�E�3��3Cln3��3�s3�?�3>��3�Ɍ3�XJ3@��3P%�3B��3`�\3�@C3��4{o�3�:�3�6�3Ș�3&��3�p�3C��3.�i3�Z3�!4�j�3��3�ڐ3a4��3爕3�&�3��p3�3n�3��3]x�3�Ȝ3��3�4���3x�3��3�D�3�ѭ3��3c-�3o�V3���3|.4rt�3di�3�lT3��o3@"�38
�3q��31�3:\�3��3�@4_�3�o�3 ��3�d�3��n3�3�3�U�3&��3Y+q3��31;�3mOr3���3~Q�3գ;4<#�3�v83ɐ�3�h�3��D3�,�3�cy3i¦3�{Y3�'4�'3�˘3��3�4��b3 ��3ڠ-3V�U3/;3��3 4�3��t3mA�3�W�3U�4�3�݌3�[�3���3��3C�3��^3�{�3}��3���3���3k?*3fc@38314��g3V�3]�q38 u3�Y3P3�5 4d�3��3M��3RѰ3�K�3e'�2�D�3��|3��u3�_�3�Z(3.t�3��3g�3u��3�<>3k�^3휊3��a3�D3ꀀ3C��3X�3LA�3[�3d<3θ<3�5�3�v{3��3?�#3��+3�?�3-<�2лa3��36��3�3!�d3�?c3�
|3 ̭3͗�3�1P3@�D3�V�3�_�3��q3p��3Y�3�tb3�4Y3|��3���35��3�3�|3�2%3��3�k�3��T3�3��%32V�3CG3Ȋm3v3Y��3Z��3@b3�.b3��&3�;23a�A3|:�3(h3��3�s�3��3 ˂3��E3t�3��3��3�q3��"3�I3�g+3-��3�nb3b�i3s�{3a�3ň3��A3{��3��?3���3Q�_3��3�L3�[3^��3��3`��3�(3�\3�6k3�}P3��+3j��2��X3��>3<1s3j�&3�.o33S�2U�4b�3��y3��43W�<3�`03�3�3�l�3
�%3ɶ�3Q��3���3,ď3c�3jB3Hr�3��35gu3�=3q/�3v�n3��3[ 3O|�3�3<��3?[3&J/3��e3s3}�~3��L3���3��93S�T3�X4���34�3��H3�a�3ɤ3��3�3F�R3;I�3U��2Dj�3t+v33�3�^3��4�-3�G�3�9�3���3��Q3�"�3'�}3}}~3]0�3���36l3�Ӗ3��2�3��3��+3�i32�3i��3��&3� j3��13� �3���2T�4��2�k3�^93Dۼ2?�>3��C3l�3�
3�Y�3�O�3���30pd3��3[&Z3E6X3��2)l3��3	<3��?3%V�3�=,3X�)3���3��
4��q3���3�G�3J�3�Wd3�K3t~C34� 3���3�L�3J��3TV�3.i$3��3+�3w�L3�C83��3z��3T!G3<�3�t�3W��2)�31��3HjK3	@�3�{�3#��2S�3��v3�K�3�Z23�R3:��32�32bH3i��2g�3��H3G,3��}3�0�2��3�3q��3�3:�3��3��3��*3�5�3��y3n@�3�(3�$�3���3��h3e��3�:�3;��3|�3!�3�<�3~�3hy&3T��3')3�ù38S3ϑ�3!ߖ3�x3T��3�D�3g�3H��3�V�3��i341�3;�3к�3�N3���3�o�3]��3���3Ի�2[��3�3:gY3B�3��K3�ث3K��3P7�3��N3�\�3��Y3��$4
L�31��3��3�ۛ3>@/3
Ae30�3�zW3�3ߜ�3���3^E�3�eb3�w3�Uk3�]l3n~�3p�4�S�3���2�8�3�3&��3�np3,}B4�w�3�E�30�>3#tx39��3�$`3�n�3��L3B�l3�!W4P��3��R3]�3���3�v�3�� 3~��3��3��y3TjI3$0q3�A3��"3��3�XT4%�o3=��3.�P3�V3��3���3���3�+3̪3�k�3���3W�C3�K3tޟ3��V3�3bF�3*U3�ݣ3��3ou�3���3�$e3x�d3��4�13Cy3)ۂ3��3�g<3�~�3~�3ݘ63*`�3���3��3@F3�@�3$�3�4xx_3�޹3r4�3!�3��q3��3Ă&3kj�3P�3\H:4�ʳ3��3��03B�%3��3(�}3{s�3/oj3Z�3 ��3kb�3�b3ˎH3Ǯ�3̛�3;8#3&��3Q!3$cF3Y�+3&(�3`�[3q��3/a=3U�3��A3���3�@3(�s3o�&3�&P3,�z3�>3���3��3�A�3Kߘ3~Q�2�\S3㾢3j3d�d3qL?3]��3Xz|3�Ǥ3!��3�[3Z�P3Ȥ4�}u3���3)9�3�`�3\�I3C��3���3&f<3���3kð3d�}3�}�3�?30��3��3^C3苄3TT_3{ʣ3�b�3Ra�3"3� 3u�63P%4�.Y3ȹ�3b�j3�'3?%:3���3�YT3�3��*3�p�3��3p��3sQx3��3�ƒ3�3��3\�\3�Sj3K�"3p�3�Y3l D35W3���3�,�3�3n3uЙ3%�3#�S3HkZ3�R3O�73���3ώ}3E*@3��53�@>3b� 3G2�2�D73V�3~F�34�3�\�3x��3Q0|3a`3a͟3mu3}�v3?�h3��^3� <3r3��34u3�3�>�3.�34�3�E>3x�:3�j=3i2/3�<\3��k3G�u3"�13���3/��3��S3�v�2��37R�2NT63Ayl3!�Q3�*�2�e`3g�(3!@3)iU3�P�3�f�3[�3H*�2-�{3�I;3�3O�F3���2ى3�=K3��3�0b3�'y3k��3E}4�M3V8z3N(,3��k3�7�3Ώ3+�3��"3�9�3���3�_3~Q�2d��2r�&3^�M3��2��3�o13���3��3-D�3�D3�+�2D6-3Y�3�.393�+P33n|3��3�Q3��3T�-3O�3��z3�Ɓ3qx3_��2-܄3츇3��3�\3��c3P,3d%3���3DZ3��3n�A3�֭3�u3�8O3��*3�<�3��3v3�a3D�2���3�w�3�-h3���3��2K�3Qv�3�|s3�wE3�83A�Q3�y3�3��n3^�3��3�W�3��2W�A3b�3uV3W6�3�a�2�"H3��=3��3���3�ء3�j3���2¥�3W�3��2�*332��2��3�t=3�h�3�wP3ӗ93�&83[��3�s3�(3�G�3��3��3#�3Ri3(3��3�4�3�m�3�Jh3;��2ͽc3 � 3��
3���3+\3�3=&�3�v{3��3���2{�2��4�@$3:?3�J�3�@�3ݘ�3GH@3!~H3�� 3�b�3ї�3�FX3�a83��3��n3B��3�~�2FG3��3��3߿�3�ݗ3��13�Z;3IA3E��3�i3�G3R��3��3��/3Tq�2oLc3u��2=w3O��3Q�f3�c�3-)3�X�38�>3��3u�3��3��c3�W3�/�3�3&W�3��2�G�3.N=3 �h3(ٌ3��3��/3͚m3y��3�v3�g3CY�3e�3�A�3�Y93�O�3��3�.3��T3�3���3�1�2���3�3��3`d�3,��3�A3���3�eA3���38_3[�3��3
3���3e�3���3�x3�n#3�>�3�+�3��#3� 53h��3{��3Ո	3Xz�3f��3��3�u3i��3}3��3k^v3�n930�3��73�ʈ3�E3h�33j4nG�3�>3돬2��3t-�3�u3��h3>�2`Ń39�<3��3ƑJ3�ׄ31�F3�:�3͌r3v��3'q�3�93F� 3��<3�a�32�H3��I3gK�3�s�3ve(3�3L�$3+��3�QY3��3 M�2q�f3��3���3��43�~/3��>3x��3w�N3�F�3�n3HXg3��2;ܳ3R�f3�g3��<3/z�36��3�i�3)�3�J�3pEQ3H�+3��d3�W�27/3䵂3��36�3�e�3��G3�(�3�,3hj3Nz�3m��3E$3��93�<T3��2r�r3 S�3� �3͛r3��3\�13X/�3���3b�3Ζ3b�3P�33)��3y�k3���3hH3�r44��,3��3)3��3Ē�3jg�3��(3��A3zΏ3���3�e�3㐆3T�3(��3�Vw3U�<3iz3��2�˜3���2ӿ�3i�X3u<a3�3
N�3J3�K=3�� 3�)�2��2��y3��{3��$3o\23 s�3k?�3!�o3E� 30��3ޮ63k�	3�,�32,�3N�w3��3���3�93_23�=�37�3i�13�;�3S!L3��~3��3�b.3j�3�`"3��%3?��3�.�3
(|3W� 3�
c3�ک32�K3�^l3P�3ӗE3�>:3{�P3�'3��X3��H3k�E4Å�2	�3�X!3�O03ĥU3��S3�ǣ3�V�2 M�3s��3�\�3f8v3���2ӞI3��2�j3��3�t3���3PL33=�3ӅF3��4�5�3�44��3�Ψ3��3�Ns3�aY3K�3���3���3��3[��3;�3���3{�3e��3��3k `3T�L3�\�3[/�3V�d3�X�3�]	4�{�3F[3��+4�V3�x�3Um|3�̣3gB|3�4���3�ӎ3Tz~3�f4́3I%M3�`3��3>y�3�U3�\'3��3�Z�3H*�3H�3޸�3�Ul3�{�3�4mҤ3�o�3�[3\H3�|3�)�3���3��,34��3`4rI�3ǹ-3~�3��3���3��_3�d�3]f3=��3��3���30�l3	��3�l3ڈ,4�Z3�׊3zw+4eީ3C\�3���3O�3��U3�Z3q%34�}.4�˞3@�.3�!�3\��3��w3�:�3D3 �3=ɜ3w��36�73)��3 ��3�s4��A3�n3���3U�"3��C3�^�3oF�3Cc3�b�3���3��3�g�3��31�3W�	4�Yi3M]�3�M3���3hh�3��3���3ƅ`3�g3��:4��3�i�3�h3��3I�3ê3�c�3V�73���3y@4g��3)r4I�93�B�3r�3��3R�4?��3_��3��3��}3J�3�{\3/�P3e�24EŮ3D��347�3j�3h��3G7�3�B�3��3.�3G��3M��3*W�3Yͤ3C�3��3܄3�wy3o��3S��3��3$�3��3_�?3��3���3H9�3,��3e��3	&43�y�37��38��3��3�H�3C��3�c�3���3��!3_@�3�#~3*%�3��3C�g3�9�3.�3�B�3A��3C�53qj3�e4�f63$8�3�R�3��3�DV3�CN3�
�3<�p3��3J4)S4h��3��*3&9�3���3j��3&'�3
_`3g%4�&�3��`4M��3k�X3� �3�x4�u�3�:3�Z�3���3�rA3���3"�3��Y3���3v'4
��32��3v@�2,X3S�3���2���3�`L3"��3	(�3���3o��3u<f3�	3(E�3Hg�2�3cY3�a3�c3#�C3e3;K3�*
3�]u3
�f30=3�T 3��3��3%�2�g3�M�2�Z3�=3��O3��H3�S
3�$38I83�g3��23�.3(�:3�u3e3w5Y3h�"3�3���3(�3��_3�2un�3s�*3��73)�J3/\L3RB3ԑ3��K3գT3�3'S3��3��3��w3�GU3�%i3L��2[Sr3KE3��3(?3 �3�?3
u3Iv3��3�H�3|��2v
�23�3FV�3`y83{�3{]3;Q.3"�3̢�3�3�X+3��z3a��2��3��W3I23�G3U�G3�ղ3!Z63()@3�3N[3�L3@��2�d3��3!�3| /3�Y�3�w)3}3�3#�3��3��Z3�!3'3j$z3�e�3��Y3��H3!�3��3ϕ[3���2�25�v3�3�
3��V3��N3s,53f/:3�3bc�2e,3Ƙ;3��3�zV3rjx3\�_3 
�3`ZZ3� =3��~3/3�^.3�6�3�&p3�1:3���2�I�3̘B3�O3)��3��2�x3���27��3bY
3��J3)"3_��3�3]�33$ 3�!3�bD3�9y3�x�3�(�2K=3��}3'�37I3��'3�2S3��(3�j3�;v3��i2h��3��A3@!)3�?�2��R3��t3Qs�3$�!3`�
3C�3B�W3�y3t�O3��l3���2X_3o��3��c3��3��63��3:E>3��3/?�3�+�2�3L�03��4�3L��2�"k3M �3{�'3��)3O3��;3zC�2<m$373f� 3.�?3��3*�3#�A3�i�2��E3�!�2[��3FI3��3X'Z3�X�2.��3�t!3�3�H 3���3�}�26�03L�3��3�3f93�,I3�ر2oq3�Z�3~(Y3��3<��2�{�3J��3��3Ɏ35��2�xT3.��2"l}3Bx3���3��[3��3H�3~'~39�%3��W3��3X��3^1�3$�3L-Q3��30�3�ڮ3��M3�3��43���2�I3\AI3g͋3ʼ3u�3L\�3�V3�z3��*4}L3�nM3��E3���3v	3�6�3�1g3��%3�(o3�4��3�Sw3Wj=3g�k3ȼ*3��i3A�@3�w3Dv�3<�S3���3__q3�؉3i�3���3�-p3|y379L3��q3:�]3V�3S^�3)33�{�3��3�vs3��a3�3��x3�3�PA3Qe\3�QS3�c�3,�B3毶3cbk30`�3�c/3�94�G�3�k3u�3���3"5t3�J�3ջ4��L3`ܐ3)4��3f3�-3�VM3�\�3�#z3bf3�E3}j�3�s3��3aVl3f�N3��)3��3��Q3�be3���3μ�3-�H3��3��k3��3)�3���3���3�;3�.3}�3?�}3~3��3��R3*|3�:>3�I�3�k3��s3�$s3��3;�v38�3rb_3v�3��{3�z}3�-�3�+T3�8�3���3O� 4�3��c3[��3��3K+3��t31�G3G��3�X_3�λ3�s�3�W3m�?3�Z�3{��2xT�3���3�\3�_3�"z3���3u.E3��l3��4=&�3y$�3-�|3�4�3�3i�N3��3���2�+�3�g(3`Ź3���3 G3Z�|3�Z�3��3�Ѯ3P��3`�f3��3��x3h�3���3���3T�3]��3��3�C3�߶3�{$3UEt3ɗ�3�Y3�\3x�N37L"4��}3�'3j�3�G�3�|3��Q3���3���3a`x3�
\3��r3kP%3zͭ3f$�3��3���3�K3���3�>�3&�q3�Cj3�3���3,BD3��3�^3K�H3�K3704{�3��3�n�3��I3��N3w��3�ճ3��&3��3��3Y�3/n�376Y3�KH3�jy3��3��L3��2 ��3d��3#'�3TbS3嘛3�Pj3U�#4���3�G�3���3}�3[h3&�3�x�3�8�3 ��3E��3?Z�3���3�7�3�	4��3%&�3���3�&|35ˮ3�o�3V�3I��3"]�38��3�84���3�4G�4�;74w��3Ȝ4���3�d�3�S�3Z�3��4�"$4���3��4&h�3G6�3G��3��3��3�$4���3��3��3��[3��4��3z��3��3���3fY�3���3���3T��3k��3���3�4�3OvD30G3�g�3N�z3�ĉ38\�3gb�3y*�3d��3#w4P�3��3�'�3
�4��3��3>�3c�3��3��3�t�3T�i39�3�G%4E4�S�3Z�3mڴ3��3�3�]3j'�3P�4�ۑ3&�3�3d3u�3B��31�43��3F�3�
Q3�j3��3��35�3�*�2+W�3��4� �3�:E3%$73Kt�3J��3kˌ3��3,I�3�9�3���3��4It�3̊3�"�3�/[4���3�5�3���3�j4�ԉ3K<�33��3��3�4t�4��4]��3��X3��3D�3�b�3�I�3@?3��4�q|39e4���3Ub4��3.iw4-�3 R�3��3HA4�M�3�ǽ3��3�6�3,��3��,4�4��3�0�3f4�3"��3>�3��3$N�3��3�M�3�"�3Գ�3��3�>/3}�?4�b�3g$F3�4[3RO�3��3}��3�a4ϝ3�>�3}o4W��3�I�3;p]3�Щ3�w�3O�34[�3`o3���3��Z3044@͞3�CY3�<�3�1�4�X�3�,�3��3=Ү3��3L�3�}�3��[3�۹3��3��	4��3'�3��3D��3Y�4D'�3��*3��
4���3`�3_)u3>Z3tv�3OUC4J�s3�۰3,��3�i&3��{3�3H�4��3���3��4�4���3p�:3ͫ3
��3ʭ�3�0�3f��3�,4�`�3�q�3-�4���3�sC3��4t�3��G3:�3	J�3 E3ߑ~3�j�3��L3c�3�2�3cG�3��3�3���3��3��2D@3iđ3�gs3��2n&�3N �3A3!E�3(I�3�g83
��3E��3��3�\�3�{3�z3�<_3�z3l2�3��3�F�3�"3�|�3[7�3�X3��.3�mi3�b�3Y�/3 A`3��3���3�vS3��&4��)32��31�[3�q�3+�Z3lKN3�a�3εv3C�V3ǉ�3���3O}3��2	5q3bq?3�J37�o3o�53-M�3�3���3mr3���3��3�&4���2q8k3-|32ʕ3+eX3��Q3.��3Q��2� �3;��3̚3�c133�3[V�3��R3h��20��3Y?3�4_3�E3�Mp3=�3�><3ѣ�3~�3��k3�a3nɂ3��y3>�O3�m3��3f�-3�fF37�3��|3��3jo83`f�3s�3��]3�.�3^()3��@3��A3���3궔3��3b�3���3x#�3�&�3o��3ʧ13��3-��3��3mT�3��l3�R:4���3 @03)[b33��3�ȿ31t3��L3�R3) �3v �3��3?%�3��3��@3264��3%��3;v�3�3 $�3��^3F�3�13Y�3�6X4�&�3IF�3���2(ڭ3̎�3I<O3$��3l-3�mp3� p3�4"S3�:3$MN3��30G3���3b�3Wk�3��E3f(�3���3'�2��3��3���3�W�30 �2Y�3�6�3�_
3_�o3)�j3楃3qe3)��3��83�3Ðx3ic#4R^F31M�3E��3��D3T�C3&�3��3�3�a�3�1�3fY�3j��3v�v3z�m3��3KH�3�Ū3�'03���3��632��3��d3�3@��2h94!n3�V�3�Y3J�3�3H�B3�6�3��:3^:�3�~�3t<�3��3�n�2q@�3Y�3g�23Ɯ�3�W<3$�3qȈ3�4dD�3/��2�i�2��=3��2���20��2Ȥ�2�<�2�53	��2�2�|�2�@3 R3*�2,)�2�n�2k��2�^�2Z#�2G�2���2�DD2%�A3���2t��2���2\�3gX�2tճ2��p2���2!�3�2��3�y�2y��2UuN3(K3�c�2Ss2��2�2��2(��2���2���2���2�Y�29�3�C�2��2�LD3���2�E�2l��2�25�2���2ug�2�}2��2o?93�p$3)�2��y2�/�2���2���2��3Ь2�}3�
�2��G3��2���2�k 3�z3��2�K
3la�2S�83*�2���2�	3�M�2D3�2��e3�V	3���2��\23L3u�3�z�2v�3���2P�2��2 �3S�3`�b2��2��3>:�2'4�2��2�
33�p2eh�2b/�2��?2��2�;3p~F3���2���2���2G��2�2s2��2�r2���2��2N��2܌�2�2�H3���2��2R��2��2V�2S��2&Ƶ2�^3�~R26��2LeP3:�2���2���2ȡ2�{�2f�2�-'3X��2P#�2`F�2^c53V��2��2	/�2�wl3�$�2q*3�r�2ӵ2E��2p��2'��2�J�2�e3�d3�Y83~�2��2UB�2K��2ZT�2Z��2��2��2m�2�*3���2�j�2h�2�13�3���2"��2��3x��2�43��2V��2`��2��3�QK3���2�Ō2�E�2p�3O%�2�3੍2=�3+�2�x*3Ix3���2^,�2�Y3��2'T�2�J�2{.�2��2���2Qq�2�ׄ2L�3g^/3�/3�`�2?��2�2��2X�3P��2���29��2��2ӼU3zY3��?2<�33J�3���2Q�3>�3"I�2��^2#�2F1�2�ѭ2}�2Qj3>#3D��2��62�V�2�H*3��2��2[�w2DG�2v?�28�2���2!��3֣�3*߮3I�s3�{�3���3qh�3e 3�g�3���3DG�33y'�3��3վ�3�ʢ3�`�3�N�3�^3�G�3m��3ʄ3�n3/��3aW�3D�3y
�3�h�3��53Gť3�3��3�SM3F��3��3y5F3kZp3���3n�3<�3f�+3�I�3:�03<�F3�j�3B3Mt�3$�"4���3C�3�9�3��3��46�3ع3ٖ�3P*�3d�3J��3�4�3�Fm3Q��3]-�3�5�3B�3;N�2�3��3;,(3��3L�=3��@3�	�3���3�>3��3P�3EF4ɲ_3��3HI�3-7�3�w�3<C�394��_3���38�J4�[4��=3�;C3Qѫ3Lv�3d�r3n*�3�"}3���3�r�3�7�3̞�3eD&3C�3� �3�^c3c�Z3C�3d�z3���3��3��u3���3��3�� 4J�3���3*3��3��3�R�3��3�Ē3�-�3!�b3��3�3�Õ3QYY3�L�3�B�3z��3씆3{;*3%��3��3��j39�/3���3�34׾ 4�p�3AXM3Y��3>��3�s?3���3��F3ր�3�Jt3���3��q3�Q3��39&n4i��3p%�3{�q3�ZB3�i^3˓�3�]�3S�3���3���3x�4�X3�:39Y�3���3rKF39�3@wu3T/G3t��3&�3�,35�3!P83��3�S�3��3u�3�M3�3F�3��4�E3R��3��?4s��3E"�3��R3� �3 .o3eh33p��3��f3��3��Z3��3��_3d�#3��3��u4��3*�3+=�3>��3[q3�;�37�y3T��2�h�3�C�3u�3Y�4>�3��3��3�3t�|3�ځ3���3ڀ36G74LI�3pb�3,�3���4�p'3+�3�33V�e3�x3���3���3�cG3�3\��3�H�3��3�%3q	�3��3��93u��3��M3
4�KT3+[�3k�3�nN3FF�2��(3�I3Ys3f��2TE-3���2��73��3�83J
�2�fd3n�33�j�2x?�2�z3��2>��2���20�2A�3�t�2��3���2AF3_�"3V�q3v��2�9 3w�2ݩD3z��2g3V3
3zq�2��3�=3�J3�N3哦2�d3��2_�R3dH3�3��-3	�2�Dl3�d3�H73\�2��13,�2]��22��2��2�I�2�G)3��2��+3FN�3�`3���2�j�2�^33�2��(3#p�2�� 3o�2��t3"m3�T�2I�C3���3���2K3���2���2�G�2�;3٤#3f�2�F
3�?3��3r��20L�2V� 3N`34��2�7b3��2��2�k�2��J3�3YL3%�2���3�$�2���2�=23��2�83/L,3���2���2`z34%�3�K'3� 3E��2�3D#�2j̗2�(E3�3��
3��2�X3[53`Z3���2	d�3P-�2d,�2�3w=3��36�)3_I3n��2�3഑3E�I3s�3�)�2w.3#Z3��"3m�-3��21�v3���2�`23<�J3#@�2���2���3h'�2�%�2g�3pe&3���2Z�3��2�b�2q�2_{P3xn&3r�2���2O�!3_j�2QI�2�c3���2��43�߻2�1N3F�2V� 3�]
3�a3�t�2�h&3�l�2��24(3Rux3b�3*�W2{3hb&3�t�3xԻ2�!3��;3��3��'3��w3�X3��3��2:�23Ĕ!3���2<�Z3���3�?�2*�2n�3�v�2�9�2��2���22�2�\3J�~3�u�3Lb3���2n��2�D3A9�2��3�1�2w/13t�2�3�8�2���2v�2��3>��2&�3y�&3�l�2�3�Y3�[B3�ˋ2��&3�GY3V��3%m3o��2�&3*3�'3��$3�h2��A3q3`�b3f�2��3X�3�Uv3�3�)b3*�M3�g3j�	3�O�3�(]3j�3��33<g3k �3�	>3(03�]3�63���2�"�3z3�6v3:�	3�ө3��z3i�L3�1�3��3ȥ=3��D3�#3:�w3�׮3H�3ټr3o�I3��33y�3�i�3
�3�T3�>�3(G3vt63+73��d3�|Y3��,3z{M3:c3R�O3�R�3M��3׮E3�`3y1�2�23�Y3d�3샼3��03T093�"�3�13^�3��3��3bS3�3��}3�3ulS3V�3 ��3_�3�3Ń3���3	�3b��3�^3��H3�=3n3Uir3�Dd3��3s��3�s�3�+3O� 3��S3W� 39�3�z3w�33�-�3?�3��3��13 &	3���2A�323�1E3eP3S�3Z�S3�Tj3MH�3o*�2�Q�3aO�3vz38o|3f3۳m31��2���2�qC3�6�2/�;3q�2���3I}G3Q�M3�?�3!C�3PvP3�,3�Wn3#�2��Z3���30��3�� 3�K3Q��3|:�3X>V3D+ 3��3<֕3y��2k63��83�-�3|�k3{]�3��3h��2�3�5�3�:3��3b�3�|35=W3go(31�b38�3<֚3�*�3���3�_3&�2AKI3��.3��
3�R3Co3Jc3��3�4�3]�2w��3�	3�p�3��^3~oY3~��2��v3���2���3�Td30��2V՞3#�3�-b3��C3��,3m�>3u�3�@�2L ]3͖(3� 3�M 3@x�3kS3�R3���3��3lm3��=3`J�3s$3� 03��3��\3�R�2�
<3@ۏ3>4�q3xRX3�vu3T��3�23O3<�2�*�3�V�2]3�-33g:�2��G3��4�� 3�3q83�I�3� 33&��2%�O3e�3w�32��3��3�/f3��2k֛3JC�3cfC3��G3�Գ2��933�<�3�is3��3b�!3�r3�NX3~��2k�3�;�2�H�2�# 3W�3���2*�3��l3s�v3�8m3C3"h=3�0�3�v3�y3��34�3��>3ͧ�3 r3PB3�x�3��3��/3��2��v3$�83ht3Y-'3SC3�-O3I
3�H3S.�3\��3�3�2b��3��3u\$3�Ve3c13�{f3;P3��3
+:3�213X��2���32)[3��n3���2Ae�3hҀ3�W3�;3��3"23�nh3�c;3��03�ج2.<3�u3�eK3m� 3223t�B3v+�2j�3p3O0�3���2���3�3� 93��38b3�[3�o�3�Ǜ3/3��F3�J�3x��3G��3�3���3�es3C#3�z3�)3w��3&�3�`�3��B3�3��)38�3��U3��2�V�2�T3���3���3i3be93,�z37I�3]�G3z�3�3��k3�,U3���2���3M��2g��2YM3|�3�2/3��{3=�3˚$3v�(3�P�3���3%�3N�63E�3P�N3��3o�~3��3�[3��J3�^3�4B3X�3tJ�3<o<3hʊ3: �3�mQ3�<�2�O23�3��74��3��{3��2��3���2���3`�v3��3~`s3��3zn3I�2�/3��3�=3��3�:K3}$3��n3�O�2�r3wU3!Wq3�3�2��4|�2d�2��2���2�R�2��a3��U3WR�2{XM3���3�23�3�s3ka3l�2��2�N3[��2�;@3 &3G�3���2P�_3�F�2���3Q�I3�KK3vD`3H��2o��2�,�3<��3��2�L3�{�3o� 3�}3��63�lw3Nh13À^3��~3�3$��3Ӷ,31�v3��*3!ڼ2�2�0�3���2%�2/�c3�n2�)�2�2�3�y3�Pu3̤�3��3�E3~�2j�T3��3�3c_P3hħ2�O3�
�2��3�z3��=3��g3�T�3z&3��J3�J3��:3ͺ3Q_�3Hd3fP3tET3�.�3���3���3P�2y[�3�u�3�3��V3��3&|3�t3�h�3��X3�+(3�V3���3��l3xO'3���2�pE3ʹ03��3vs�3��N3n�~3�>u3�3�3N�3���2���3��m3�l3��L3љ3YӐ3�83�z�3zN~39&3ZT!3�l�3�E3Sw�3�^y3	�/3f�3�PF3!D�3n�3Zwo3�B4f��3Z�W3�)�2;�3ɻ�3�� 3�/=3��2jٞ3(�3��3t,23� 3@)E3�4]t�2��^3z�p3}�3��3�	.3��3�Z�2�!n3�ێ3���3lab3��:3ɻz3�c�3uHW3�3�'23�w�3�93��U3훃3W�<3��3�4���3l�?3\w.3M��2�2�K3px�3�(3��3�~3��3�3u��2�U�3�pt3S��2EE�3�X53��3_�3�N3X~3^��37oc3�I4m��3�p>3�7a3�*3ˀ3QX36E3N~36�k3�ȕ3�GZ3�g13[�X3_�3��3��3�u\3m��2�q3q�<3Ɖ�3�_?3�?G3C�63�4�< 3�13�3�Y�3�13�V3�x�3Î"3�j$3�u�3�|�3v23[�<3t:�3y
k3��W3)eg3'��2@��3�-3�v3��i3`ͪ3ܚ3��4�yN3���2oJ3��A3� u3/Io3�f3v(3�T�3��3�q�3h&3s-)3&)o3h�j3��t3D��3	��2|��3^�W3A�A3��3
�:3�.3���36FR3�83��3ud3n$3"�2ޘ3V3L�3.%�3N�r3�`3 "3�23|3]l)3��t3�%E3D��3jX@3���3P~33b3)03�~�3��2��)30z�3��3�*W3t�\3�M13�5�2F�Z3[�3BA�3"XI3r��2�n3��'3�uJ3T>K3��/3�][3�y3y�3�g�3��$3[�T3q܆39��2�43v�X3�'	3���2�5�3�x#3�q3H3�p�3"�63g$ 3���2͝%3���2�3|3�	3��3s�2��s3i�.301j3�R3V8�3��3~f3�Z/3EVG3�E 3V�03~\�2c73&�X33�`3`}23��L39�3�c3:�|3z�3x83��b3Ò63��!32&}3Y�O3�	3��@3�U|32g=3 �<3$D�3vx3�,53$�A3=bf3q��2cO3cn3�a3� (3���2�.3:�w3�I�2Y�^3&I3r�a3�\3�y}3o�3�
3@�*3u�3L�3�U$3
kV3�7@3��@3��73�L-3�i2��3 ��3��]3��G3�S3��{3�ɒ3Ut3y'�3_�3	 M3n��3�&=3��2�v3��E3!Eo3ۃ3N�l3���2\�3�3���3#NQ3�m�2?mO32#93n`3@�3x��2��3� &3��!3�E53I�3�X�3��A3�u3{�,3�43$(3�+�3}�/3�Y3)�3ȋ�3ō>3��m3.�73���2�03]'�3hTq3�Gb3A�3��^3$d�3�[3�{u3i��3��{3,C-3E��3f=�2N��2C�.3	��3�30R^3�AP3�,3 .,3|rP3�U�3��2xo3,{4B��3޹3H-3�jX3��3��2c�3��03�3�3,��3'�B3p�U32�H3��3��|3��@3	�83�*P3�p�2.�3�63i�3q�:3集3d�3C�3JB@3�A=3�i3��3Yjf3`J�2AB�3�3\��3`�p3�Y3 D?3���3�D3�N3��x39x+3��!3/�36�d3j	3n��3�Q�3��3J�@3�E3fQ53kBp3�(r3�633�q�2���3k#3֜3W�J3o�2�~�2xG�39�3�3�03@�2sٵ2Q �3A�53�I�2��u3���3��3x3��2nk;3���2V��2��U3���2Y�k3��3\v�3y|�2t�3��2պY3��2��)3�F\3�̅3T��2��3�|3Pw3�3���30Oa3j�@3k�+3v%3p!K3��2��3��83�3G3�Ё3�cM3��3
�C3��3�"3<�c3"�3��3�W3h�L3EE3�P3;�:3�J�3�a 3ϒ3<��2�;3Ш�2�23� )3�\3=��2�"#31^n3�_3��3CW�2̞3U<3M83�x63q�g3غ2�z�2F��3&�2M30�3Lk3�S	3�
�2�}�2 al3�O�2N��2�j)3�;3�Υ2&B3H��22�3��[3r�3j3��37��2�2�3�C3�F3���2tt3�΅3�n�3ngT3,$3q33}�^3[��2
/3yU�2�3뉽2��f3�"3��2�3<��3�03	:3a��2�;'3�[�2�~�2��M3+�2�&%3-*}3�8g3E�2~H�2��?3�J�2.��2��Q3���2ܤ�2%�2(wB3���28)_3]\�2Jф3�3��	3��3�3���2NaV3��73$�3?��2Qz�3��3O�3�\3�v(3O3�R�3��`3= 3}�H3�W�2��3:�3)�2���2fT�3�2�2��3�&3�1�2�f�2˧3x3���2]d13VՆ3�F3�@%3�g�2bL�2d�36��2��3���2��3���2	�b35�D3�.3L��2ڵ�3S�26�33�k%34/�2�A-3��(3��3�3�<3{�3�d�3�bJ3!�3��m3��3�`3|�3࿶2\f3�(3?}�3$�3���2s� 3�C�3��2�3��^3�0�2k:3�o;3on'3�q3�:~3\w3��A3He3L�2:"3̉+3�3?�93!��2u�\3���2���3��03d3���2 ��3-w3v�3Z�=3���2�3N�K3�E3�}38F3�k�3�Up3`Dc3�7�2_�m3O>�2�cg3Ɛ32H"3#j3��2�\�3��+3A%3Ml#3�y�3�Q'3��E3�&3$C3\2�2"Xk3F
f3]	�3"3%��3�ar3M��3��2�;3b_T3T�3O�2<�A3Z+M3��2(��3n��3 =3�JT38��3�+3�e3�!A3G�}3Gc3�-3핒3v3r;-3	zi3�F3>~[3�3ⴐ3f$�3���2?c!3�!.3N�%3�83n\�3��3�`\33�3���3�r3���3��3��-3r� 3���3[�3��Y3�m3e�3��3���3��3%��3��3k�63�zc3�%N3ȗ3UYi3�Hm3)_*3R�>3v�u3��4�[F3� 3��F3r�B3�- 3�~.3�N�3l��2r<T3�3���3��>3��2�LK3��S30623�V=32�r3t�`3���2"�3�+3��3|C�2eW�3�TR3-�3Q�3��;31mh3���3�t�3JT73b+�3JA�3�0�3%�	3��)3���3�1�3�_F3�v3m�R3��T3���2g4!�33W_�3S5�3:�3e3	��3M��3N�I3��K3��3���3��3���3.��3A��3C�P3e��2棚3�D3�5�3V`33���3[	�3N�?3o�~33�3G�(3��(44�h3;�)3��U3�^3.w3��x3Bes3��M3w)73ѩ3�Ә3I3 �`3�z�3��2v̕3�U*3�R�2��R3:�h3n�3L�u3Gy3�`W34��3w�B3T>3��-3��93�T3��j3���3��3<��3v4���3�C33î3�x3qI3��3%��2��C3�v�3���3u�23�
:3�J3���3�G3�N�3&®3��3<�C3aye36�_3^�p3?�Z33�3�4�O�3%3^�r30>}3��\3�63sC"3�T�3�_a3Zm3��-3SJ!3( 63	��3. 3.��3@f�3òx3p<34�z3��A3�pY2ԝ�3�Z�3ӹ�3>]�3��3��3]�3�*T3M�3��O3 �3�=3�b�3�03��B3�uy3U��3 �63���3�|3�߁3��53���3E"~3��3l.B3^�3��3'�3��\3d��3�n3{O�2j�	3�ڃ3�{3�3�3+�[3B�3��$3�^480�34�3b�93�AT3~��2��3�-4Msk3'�x3@F�3u��3�ڈ3��93��3�M3`��3F�Y3�q�3��_3�Bl3\�3�?v3'�}3*;�3��4��<3Im�3��3d�3��3D]>3��b3�zJ3�vp3���3`��3a#q3�]3��3*�S3��3/�3ta�3nRb3�3[4��R3F�Q3�k3� 4KQJ3�M�3l��3���3��z3�{93��3�7�2�,43d@�3"��3�+3��53d��3�B�3~�n3_��3_Y3@#�3��3���3L;3jɂ3�3x�3���3V��3&�^3\�2�WL3�ku3Ǣu3��]3�_X3I�3G^�3�H)3xm�2�^3��3��3���3Y�*3���3*�3���3Ӓ3~�n3�!o36��3S3�e3Ru]3�u�3hcI3�"3�3�3�ن3؊�3��'3=<�3D\d3��E3Kb!3�K3�+�3J%T3)"�3�3���3_E`3�9�3��l3e��3-�s3*73R�135Y3���3;��3GJ�3��3J��3��4���3�J�3���3M��3,�[3Ex3r'�3�=k3��3�3�'4�43%e�3�
D3�<4A[@31K3�jc3?v�3Y�Y3�n�3�H�3c�?3l�y3,�4̷3U�43��V3:��3ᶌ3��3�ڶ3ת83'�Y3Q�3T�
4�)3�mK3�p�3�J�36Pq3wA13�]�3:��3*&�3õI3Fgm3̅3�C�3An46��3�	C3�=%3ǿw3��3��h3��}3�<-3s��3�3K�3��K3���2an3lE+4�3��`3̛3�/3cY�3��3Д3�+3�`�3�(r3害3���3�"�22ӌ3��53H{)3��3{�N3�f/3P�(3��G3�s�3��_3�3��3��+3�b3F��2oȤ3��3��e32�C3` D3�073敦3��93j�,3�	3N��3�S34�2��3<�3H��3R3oĎ3�N3n�24�3�G�3�K/3�n3ydK3!s3N]J3� 3%Z3:*�2��D3:�3�e�3�$a3���25�%3��34�c3��,3��53E  37�3�f73,EE3q��2��2qo�3�n�2SHO3��"3jP33�"�2�w3L�W3��L3��>3��A3�#�3âP3��2O�3^�3� �2/9g3eL3��+3�3fj�3�	3�F3FEI3���3s 73�L~3,��2D!I3D�<3 �33),3Sxn3g�V3$ߴ3 	@3E 3���2�3��f3�_�2IM�2U^3�663�O3��d36G43��3�g>3혼3�F�2��-3�4=3�M3���2��3�Q3 �3lV63�>�3��3-[3���2g�%3�[C373�"O3�t�22G3 �3�RS3��3�:3J�$3�+�3G�3ӳ�3�˅3��[3\�+3}�%3�_3��3L
q3�6�3�؍3��3�J�2t��3�@03ձ�2�K3߼�2w��3£3�"�3-��2��)3��3qѵ3�i3c�p3O��2��	3A�3�-13�`3Ey33��3���3�3�d3���2�V3�G3�N3�/3�{3��3̬�2J�3>3K8�2��G3R�4��3A�3Z�U3��3�)3I�3��43�(3,�r3��3���3z3!�2ⓝ3�^3L2H3��W3Kc�2���2i��2@Y343��C3H3%��3�T3�)3��3�O43�w3a��3d�m3
�\3^_63%��3��3�3�A�22Y�3��[3�B}3�I3�=*3z23J3���3q�@3$�3�6�2�Q4]��2�+�2-3�`K3A3ʏw3Dq3,X�2Dhm3�o�3���3�73�z�2�63��]3[��2���3��3 ��3*�3:�3��?3�J^3q43�j�3Z,3�`3Q.3B��3���2~��3��r3~�2~�3���3��y37�N3nB�2��_3�wY3[�2�	3]�U3��a3�q3��s3�p�3_��2p�H3q�}3kNO3v��3~uL3n��3�2�3�a73LC�2��Y3頫3��3�H93���2.nu3�dl3��3]�3�x�2}��3�73V�R3�	
3MxS3�|a3,e�3��=3#��2�j%3�'3qA�2V31�36�	3J�43>�`3�Y�3�*�3���2���3uW43�3%�
3u�2�>G3���2V�&3�F3�?
3.�T3��3F�P3��g3�\�2پ�2�7B3�43���3J��2@3�Ő3$�S3g3�m2b�23"ߋ3��3䌯3��>3d<3��)3��P3�[3I�3Ep�2�	q3��X3
�*3�"3�3��w3B܊3o[l3�3z::3���3�Sr33
53�D�2�+3b3#�(3NR3	U�2�FF3>�@3W~X3̅i3�:13$=.3J�3z�3��?3�3��V3��B3�u3-�33n��2�i83�i93{Y�3a�D3$J3��#3F�[35�3-~W3\�3a�O3�i�2&�z3��"3r�Q3��2�q4�G�3��A3!*(3*��243�{>3fwO3
��2�0Y3G#�3<�g3B�2=˓2ww�3�2�du3�?3V�2�3�y36ӗ3U'3|��23�3��3}��2��$3��73��3���2��,3���3��83��3�W�3��L3t�53@��2�t3g�_3�3G�3�3�G�3�J=3;S�3%� 3��2s+Y3ŭ4��A3_�*3�ܲ3��3_]�2	�:3~�:3V�2u+^3�lc3��3���3�3��	3uu3I[D3��3��2�Fb3,�K3J3x�i3�vM3�}V2OP�3D�13���2D�2��2%x�2�,�2�3�o�2�F�3�A�3�F3��03|��2��3��H3,��2���3��3�[3��y2�ض3���3vl43�9d3~]�3ۊ3��>3�3"��2&��2iP3E E3��D3^�3��{3x�]3�U03�3;'V3��&3
	3~`"3��3.�3��2��!3i3iKH3�� 3��3��2�Fv3��3�43�)�2@�o3���2f-(3
%3g|�3!73|�3�F�27�83��M3.$�2n��3�!3	�"3=3��3��M3�V3�3(�{3]53��3*� 3#�3�v�2n?3?O!3��2�IM3QP�3rb?3��2H��2��3��396�2=R3e��2nOn3ە�2�C 3�-�22��3���2('�3�_�2]��2!�<3���2Q��2�3fa3F�3�36x�3��\3hl�2@��2�)�2KIr3��3��I3%X37S3!�2��I3$�3'��2�v�2*�3�n�2�<3*�
3H��2z��2�s3��3���2%3�ܝ3ށ3��3YW�2d}Y3&�3x:�2�;"3�+3�<S3@��2�13c�3E�Z3���2U}�3G�3yO3��x3��B3�^�2c�3�tb3$?�2ވ3�!463tC3NΈ2&�`3	�T3�*�2�P3/�2\	3���2	:3�)3qB�2���2t;37��2vV�2I�3N�3\��2��{3�Â3
n�253��3��2�m�2ޙ
3}'=3�?-3�3t43*=�2��2l�2�`3�K3�3&3���27߃3�3tQV3�E3_|�2��
3��	3o9w3���2Rv3v$S3���3�J3��22�t36AN3��43��3� 3j�M3�F�2e�3�P3���2�3�2y�3�$�2/< 37��2�n3)d�21O=3�.3H�2F�3�~3k�/3�+Z3�'�2w�D3�3��2e�33M��2�27��2cW�3Mc=3[�3�Y�2da3���2ĥ33���2��3U�<3%�I3-9�2y�^3X`~3\M_3��2�93�_3Ki�2��2��3��2'��3��"3�%3�4�2��3[�s3Ll�3,� 3��t3�k>3��3"BF31�34{3�Az3�3Pw�3M�3W�z3��I3o��348h3j�2�)c3�-3�h�3�"3f4�3j�V3e��3��E3��4�a3P��3j�k3n�j3��3���3�3�Q 3[U3P�3P�3�خ3�I3���3���3 �3�`3 �Y3�T�3uj3��3�
K3�<�3qr3�A�3��E3��\3�3��p3ڊC3 R,3ö�3�3���3�;84�[�3��y3�p�2Wx3��y3`�*3R�3��3ֲ�3���2��3 �+3rQ�3m5-3W�C4�3�$�3,��3��3��w3��p3�K�3��2&a�3�>4�M�3�|W3O>3�13`l_3�=3�3ف 3Q5�3��?3i��3'�232?C3u3$��3}�u30d35[3��#3�R�3C��3���3�?3bը3�L�3���3��M3.#3;��3?m3Db3!�3�� 3��i3���3�}�3<�V3�M�3���3�4꺇3�k�3�/X3=C�3�a3j�V3�Sx3=�b3��3���3�q�3�3;K3���3�5�3�8"4$#�3�֒3^��3�/3�<�3��.3z�{3F3U|<4�Y3�5�3��r3�]�3�_13-�3@��3�Pm3#!3" �3�*�3{��3�A�2H?�3n��3?x3�Y�3�'3�~3�/�2��4�؄3M'�3$B.3�g�3+�3z6�3��a3243�-=30�3�_�3N�13"�d3�h�3j^�3�̉3;3���3�,�37E53�>�3�<V35��3�F>3l8�3�9i3P�]3�R3��3hR�3t�3��3�U3�Pf3Y�4gl3��r3V�3|�3��34�3P�w3~�3ez�3�mv3�×3�'�3�%4[�`3���33��g3s�43��44^q�3�e3s�/3���2�W3{�3ﰨ3�mB3��3S4ݾ3Kja3&��2�[4�r3���3��G3VNT3#�4�@ 3���3��3}��3��\3���3��3�g3��3�3��83@s3��g3fFJ3��y3��3\��3���2��[3"&�3B�33�(3 b/3�:3@�3��P3ϥ@3��V3+�F3�O3�6�3�-3J 3��<3��h3�6O3gR3�3�3��3Ԫ3�_x3�}3*�3w^y3�ԍ3�M+3��L3��@3}�63p�2�3��H3�FI3t<3{�3_�?3��,3b�37\w3-�2e�3q�3ξ3#�2��3^�p3]C73m�2��3&�V3�V�2l�-3�� 3���3�FP3潁3J�2�y�3�$3g�3\d3te�2*�J3wt3sd�3��73*��3�3q��3r��3E�t3-Fg3�{�2��3��3�'3�u3��2u��3ex3N��3c"3�3��2�s3o�30d3��3/3�X&3Ѐ�3��.3��2u�3�/�3�ݑ3b� 3}��2-��3�:}3�3Ǉ73*�23�33��'3�C�3qiG3~R3��93x��3��2�)]3ɱ4�*�3X�(3�h3�e3� 3ۉ~3�e3�p3G�"3l�B3���3��}3]03�Hc3�x�2��F3.�W3��&3Q.S3�T�3��>32Z�3K63ɻ3�z}3��)3�3��_3��o3;"3�[�3�
48[�3�W3y�Q3�]3�s3�/3<��3__�2J��3���2+C�3��q3�,3=3��3�=3�3�A3�?3l[3�A]3�3��2>�)3k�3�c�3b�2j �2���3�p3�,�2TLp3L�3I��2N�u2�Ȥ3��3K�63���3ѿ�3ϗ3�?�3t/�3��3'~s3�J'3�ˏ3q�Z3T~h3W'�3��J3F�T3_��2��3x��3���3w�$3�_�2�M3��3�&v36$;3��2*��24�4�F3�C43d�D3��3�()3�g3��3&h�2d#3�3՘3|V3�s
3��,3��!3B3"ل3+\�2Ɛ�3jO3M3_?3���3Q]�39"�3G�n3GEk3�
�3N��3��h3?5�3[YH3k��3�FQ3���3Z��3p�\3�w3I�3y�B37�	3���3923oN31�x3�|�3l�3���3�&�3.S�3��3w�I3��3&�i3�03z�s3*Q�3�3�S3�	4��3���3>3���3�ʓ3E3|߈3�>W3{(�3��3��3�]J3%��3�3��
4��o3��3�m�3Şg3�oZ3C<�3�{�3,�F3*�3[	�3���3���2~~3}7�3��S38�*3V-g3�W�3�:�3l�b3���3�634$D3�t�3�@4�#^3�i36j3k�b3G�3�3r3w/�3��93��3M/�3Z/�3���3�C	3UhW3�:�3���2��M3�i$3!T3��3͕�33&Kq3^*+3e��3`J3O�3�g3o�A3�_83[Z�3���3�3���3t:�3��3髚3x�2�,�3$k3f,3^N3��X3"h�3�3-�3f?35�r3=|�3�4�4,3��O3�g/3��l3$͆3�l�3dM^3�3��O3���3�{�3��l3��3�\�3��3�J�3�X'3�_Q3���3TF3Zk�3��`3��3&fH3��4>ڃ3Ґ�3v�'3B��3��k3�G3��3�S�2��3�4(��39[3B� 3���3��D3��M3`C73�L3�Ye3�F=3���3��u3��3���3�v�3Bw 33F23]�e3�V3�z3ϓ�3||3:�$35�63w�s3sk|3`�3z�3��(3��3��"3�;�3�.3ŕ3K�"3��23yX3�.3H#3s�3SG[3��h3��I3=&3IJ`33�Y3ݙ�3�΀3R�o37��3�z 4�xf33%3斀3���39Z3?[73��&3Kv�3<�3�J3Ω53v��2�>�2e�$4^-$3W6)3�3`�M3X��2��m3��^3o�3��H3�}3ū�3k]3^�3�%A3���3�3�d3�4�2�J�3�#3y��3�J3Z{�37/3��3%u13�m�3�\3�T�3��38�3YɆ3�^D3�a�3��3#��3�B�3�K3~�3?G�3���32b�3�3���3�r^3�Ʌ3��}3���3?�3�3<a<3=}�3O�j3��n3���3�/�3qxi3�V@39uE3��3��w3wб3��3��+3P�3��3_9�3c�03�]�3�3��p3�@�3~$�3���3e�3=��3vpN31�3P�83� �3-��3���3�!3ۍC3Oj�3I�49��3n�25Y�3��3�^33L��3���2�u�3P�3��
4̚�3�l�3�/30Q4t�3^�P3ߛ�3R��3��h3��3��/3��>3��}3"��3ӻ~3�f3�E3(s�3Q��3>EL3
�3f�3Y�3WCZ3�4�-�3�.3��3�Z4u3|��3@�\3.Ѓ3�d35A�3,�3�h_3�W3NB�38�4�8�3�� 3��3���3��t3Jl}3�	�2p��3M43J=�3zR�38\p3��3:R+4(ť3�D3uGI3��f3�8X3��:3�63|�T3�7�3(��3'��3]X3�@\3c*3Ks3,A3��33�|3�ɔ3�63̓~3f�F3�y�3KM^3��B4�D�3"��3�L]3��q3P��3M]a3k�V3�_<3�BC3��4@��32:�3ah,3�3���3�3���33Fp3�3�30d3T��3�n�3�Q!3$O�3=��3T�s3��3�ݳ3���3h&�3+��3�lo3=�3g�W3 ��3r��3W=;3n I3E@�3�-K3��'3��3�W�32�H3��3�PJ4�g3En�3��'3_4�ӻ3*�3J.�3ޅ�3���3W��3��3�+K3���3/�3��3uf{3��e3J�3���3�P�3���3au33M�38S�3�^�3C�O3#Z63p	13���3Jc|3'��3�s3$W�3c�d36(�3���3��M3g�=3��]3�J�3^��3��A3P��3>�3t�B3\��3pd3��3�a3$��3W��3p\m3<�2L;L3�k�2��3w�
3&�D3��	3��c3a�53�3{� 3��13��,3��23M7+3�!�3��3S��23�c3��B3�I�2��~3�J3B��2��3ɣt3*3Q�:3�3}��2�3�D38��2�C3��X3'�3�A3�[#3B��2���2U3F�+3,� 3bܿ2��53IL3�P�3�a3���3�
�2���3�%X3[�3��#3>��3� 3�	3
�3���2�t3�y4��33��2 �2s�/3�23-;�2 �3�F&3��/3
!�2�l3���2�{	3�3y��3u7�2�[�2>��2�%�22��2�|3L�^3�@�2��d3��38�Y3�b�3�5�2!]�3(�*3�3!5;3]��2j�?3�3�<3��3a
3�-�2���3�{R3��d3�h�2�.�2ӵ�2q�{3��N3V��2�7,3?��3eF33�2s�3�;43(N�27.�2�'3-R�2��3h�3�}F3@3ȻL3�xs3/�w3Pg�2� 3��\3F,3nW73�3~I3a��2�13jM)37)[3�s3fF�2H�83s)L3*Ǚ3i�_3�83�_3jy�2C6�2�M	3��39�2�6�3;�
33��3��3DԀ2 �J32�&3�Y3��3/��3'�3�3`�2��A3�N�2X*�2�T 3��2F=L3߃�2�ć3 p63 �83�093"`�3�3��%3�2N��2I�/3�[>3�0$3���2�u33n�v39�(3��U3ܖ�2Y�A33�!�2H),3�*3��s3���2�j3�3�@Y3���2���3��3s�'3�'3s,�2���2��M3+�239��2Ƽz3�o�32tz3�Z43-7�2
[j3�633�V3��3�6�3�f�2��3��37
g3t�2��3C3�t3.�3	�3cs3A�3bJ<3zԺ2�c�2�3I3>�23��2�e3S�3���2��a3ڲ�2��F3��2�}y3��3�̧3˻73g4�3�z�3���3S"3&��3�Z!3ǈ|3��X3�#�3��@3;�3$��3w�m3�M3~�x3�y=3�v3)/(3W�>3 �3��3���30c3���3��!3�r4Ě93��L30;�3��n3~H3�>�3�GT3؅K3y�|31�3��3�x�3_�3���3O�B3�@�2v �3Qܒ3c�3�MY3{�3�}~35��31�
3���3jAP3�8�3?ro3��3��3�m=3�X�3"?43l 83]h�3�ͼ3�o3^�93s�3�t3B�(3gZD33��{3m"3�#�30:T3�#^3(�93���3�E!3�&3��?3y�j3f*�2�V�3�٥3�%3?�P3��3���3�L3�3/x�3Nʙ3/3h(`3�jo3 �3�n83�v�3i��37�C3�� 3���3í3=j�3��R3�x3��a3�GG3(�*3ɗ3\�3��3�83�~F3�&$3�ق3��n3`X3�r�3l�!3 w3�X33�[v3�aL3 ˆ32�#3@��3
�43��13ۍ	3M<�3�G$3h�k3�X�3��2 y�3z�3B/{36)�3�&3*�3A�3���2�t3�a3G��3�R43%��3�M3z/�3+�>3�3�E3�F�3��3$#>3�V53���3�7�3�2!3�5A3���3L˱3�3��13(c�3��d3���3(��3oH�2Ӻ�3��"3�x�3��Z3�߹3��e3��33�d3�`b3�93�33F3��3���3�+3p�31G�3���3�e3
�]3�s�3�pl3��34�g3᱃34JI3b�@3�� 4���3�{3�A3�@=4���3#;�3%Y�3_:3p��3s�^3e
\3\�3(z3̀4GK�33zJ3Mb�3��3��R3�FA3ZlI3)��3&p3 �3ZIF3�qQ3]�3�>�3�$	3��K3�b�3�Ǧ3��2��A3C<3��)3�v?3镺3���3l��3��3�X�3��3d�3�3[�2=3[3�TQ3㇐3�3&3�3��3	3�33�K3͕�2X@93cR�2���2`�+3L,\3]E*3/�H3}�	3��3ctX3��o2<"�2�Z3��2�y3�u�3�	m3Ś�2�+3(u�3���2?5�2�#3j��2��2Q�3��\3��3C�[3�
a3�o/3� 3f��2H��3qo3�×2�X3��f3i;3��2��x3C�p3��83/�2,��30�2�Y]33�2��23�`3��+3t�3�N3�i3��k3��2��3�w3�4+3���2��V3A
�2��Z3��.3\c3�N�2ͯ3nZa3�̻3��3�A3+�_3T��2+ve3�f3>�,3�X33HWI3���3,!3��3N 333g3<�2o�3w-3)�+32�(3͑Z3>\�2x�2�0�20]v3���2�a
3� 3O3\(3T=38�H3�V�22��2O\3�}^3�'3Γ�2�Ą3H�
3�2��'3ί2�3�u�2��3��3O�m3�33��3��*3�E 3t�3|x3�3*3 +3E�2,3"Ʉ3
�234@�3+�2�>3��=3��2�IY3R�37�d3��3���2׸�2��!3�l�2)K94�W3aO3�#�2Ӡ�2�3��2԰�2nt3�J43f��31cJ3�3U�2-o3��2�ɧ2J%o3<��21�$3*\13��3���2b�3g--3>�p3Ʀ3�3�c93�M�2H��2fP3)�237v�2��I3��3�J3�[r3z\�2q�y3�-$3a�2%�K3A�3�23�3�
D3m�3�>3]f�2�[�3�8$3*A�2��g3�`%3	��2���2w'3�53S�63/�'3��3<�53b��2�rY3�`3��(3S3$��2�rA3��2ok<3�y3���2�+3Fo4/��2.}�2�B�2�?�2�_�23C 3r�83O�2(�3�T�3��3��2��o2�)'3-�23�/3��3�׏2���2'3�2�3^3s��3l�^3U��3f�A3���3$�b3r�U3�U.3�a�3��V3<ޏ3*{)3�4��3=e�3�23�o�3�M'3e}3�.3}�3m`R3��3h2�3�c�3t4~3VV�3���3��37ΐ3��d3���3̭h3i�_3�9�3��S3軅3��3��3��3�0$3=$�3�3qq3��3ߑR3��q3�{�3�	�3Jq�3JL�3��=3�w�3���3w\3X3:_�3
D~3�V�3wN94MX 3�e�3��4�3��C3Go3!V�3�b�3#Q3puh3���3|,�3��Q3��3��!3S�a3]�b32��3�++3��S3���3�Ro3�@"3 �L3��3�&&3��3�4��3e�3�M"31�i3���3�Z�3
03�(3J6�3bR3��3�)!3a�)3u&N3�G4A:3�D3��%3Lg3��p3Z��3-�373���3�i�3\1�3_�3�R3��30W^3(�3%gZ3#�K3�Fk3�53%!�3�%�3~kY3VkH3���3 %K3�g�3$�A3Į!3�@3J�t3Ƣ�3��3��33��3p�3�Fi3�73#b�3f8�3_�3i�3W�F3��3�YC3>+�3k�3��3WZ3�=4��o3�OR34 �2 F^32UZ3Cj�3[Lu3�Y3J4Y3�j 4z�3kDA3�r�2+Ǆ3��p3�>/3	K�3*��2�b�3�v3^��3��t30�l3m�S3>4Y63BNc3�X�3s��3�S�27�m39k3f�O3�uZ3���3�k�3�`R3o�3�:�3��V3��13DՆ3-B[3�؟33!��3�H3D1�3�`@3�P4� B3N�n3%Y�3}/i3��
3�L�3�.�3��3J��3��3*��3��3+�23-53��3��R3v1�3.,33$~3AS3z�3gw�3ZD3�;3�R�3*#J3�/3�u53o3��3��3HM�3R&43�GN3;��3t�3Ak3�E3�)�3F��3�~93�ע3@3i3��:3��3M��3�i3��z3�� 4�r3@�D33�J3#VE3��3�i3��3%�R3�+3Ȳ?3�4�y�3J�R3��I3���3,tI3�YD3I))3�[^3��F3�x/3K��3o��3v�3eת3�m4�{R3Tn�3?z�3��p3�A3^�{3�z�3�D�2$�d3�3��y3�p3���2k��3$��3%sl3Sf_3�B@3��43	�+3_'�3�,3�}�3;�K3���3��%363):3k�Y3,x"3�K[3��3���2��73o��3n�l3��3�X3�l~3��:3��27�Q3�m'3�3�rJ3�O�32/3 %3"�375�3_�/3��]3y�t3��3�i/3Z<�3��R3��"3v�3�L�3D��3cc!3۵3��3�Z3)=�3hD\3�843R�3k�H3��3R�&3�3�;53q^=4��3�L3��H3lt3qA+37��3zX�3_s 3 �q3F�3숚3�A3H�2�u4�}3
�N3�.3%	+3�
�3+�3L�3;\3^D3�*3Z�3'W^3�223�cG3m@/3jƁ3_1�3(U�3��G3B1j36��3��M3��3��33�3�|3߃
4:}�3��$3�-�3�R3�(�3YN3�Y3�Q3�i84��J3�x�3�?q3�I31A3��3��f3��3)�^3@i4�@3߾{3�3��x3�|3G�3v�3���3���3�D�3Y��3�R3*.T3QO�3`��39i�32�v3s�\3͡3��A3[G3d��3��`3g�m3��3��{3��H3�+83�9�3	p�3��u3�s3d��2��3O3i��3��3��3��S3���3L�3L��3k�3�dj3��H3iu3��
4�N3��83��'4�W�3���3��3!ύ3D;�3Hp�3��F3��3���3/�3�ܜ3(,g3u�3L%:3w^4qp63�~3zA/3@�3M�3fl3���3ť3��W3OV�3,҅3�>�3
6W3+b�3�fe3��3Wcq3��3��
4.qj3��3��31�3t�B3�4�3�3��B3�543�4�3��\32�3|ǁ3�M3�Ik3�,�3���3 �3wO"3өo3��3�AF3�hu3�t�3��13�m)3��3,Ȣ3�T3��39P4J�@3L$S39�M3�z�3�z3;��3�؇3��2�]�3��~3to�3�Bb3�n�2
[�2Iۥ3G��3��]3`�I3̓�3�5p3�gi3ÿ3��3]3e��3�ʌ3�U*3-�3�3S3-v�2*=3��3��2���3o�3L��3=F�3���2ͯ3ï(3��@3_v3�� 3�1�3)~�2�w�3��3*�3�?t3��4�p3�u3�3U�~3<=a3��P3��T3m�3�+�3�q�3��3O�3�S"3fQ3Ca3�T3��3��3�lh38�+3�dg3�G3�'E3߁93(��3k�I3lN+3��?3��3�.3��3Ե�3f�`3�'�3�&�3o�3���3�B13��3��o3�3i�e3-�i3��3w|{3=��3�۔3��13ەO3e�)4VX[3�$~3�035�3�Y*3T~�37�3��B3��[3j��3"��3�*3��t3;�R31}_3���2u�3J�5311�3�CE3��r3�#�3g�p3-�3k0#4�?�3���3�r�3:ć3l��3�V�3X~�3��=3��v3��3SM�3�:�3X�3���3;K3][3�Z3�L�2���3�73�X3��^3��3�j�3�|)4J{3*+�3�׸3�l�3q 3�!�3y�c3&�3*`�34��3I�3Z�3lz93�4`3��3�+3�K�3s�?3na�3�fB3R��3RvE33v3���2�t
4��[3E|3�}3�p3��3��3H��3,��2]M�3�ݎ3�۲3���3�s3XE3���3��3Ջ�3�]3[�3r#3��J3��z3$`�3���2]�43��2tv53��93�7a3���2?l3]��3��24��3c��3��3n�X3�[�2&��3��^36C-3��3MV3�:3��-3q��3&�>3E$�3ζ�3���3U\{3H�;3���3��e4.J�3�x3~�3�]3,�3��4��3�Y�3�`3��4�I�3���3��l3��p3l��3�m36��3��3���3���3�{4<�v3GŔ3]��3�Ϥ3X�A3�w�3QР3�[3�R�3�*�3o?4�a�3���3'�4�2�3NĐ3-��3�\�3��3V]P3���3���3���3F��3O�04ʘG3*�3��3�J�3��3o_R3�>�3_I�3���3*�M4��4zpz3�3�3
>�3s¢3�n46��3{�4͚3 �3��33S�3�3�O4;�J3X�3��3٫�3t�3��3qO4�3��3N�41]�32��3�EW3D��3�%�3��3Il�3!y�3��4<�3>�3z�3��z3�w�3�%4���3��3�M�3��3�H4Iv�3���3��r3g�40K�3E�34���37 D3�|*4�;4v�3��3U�53:34BiQ3�w�3��3�k3���3�O4-h3���3w4�3%��3#��3�F4u��3�*3O{�3;;�3�v�3b��3$x+3�,&4��3뀩3��3�S�3`Z�3�"�3�Ɯ3�Ԯ3MN3��3~x-4�(�3�b�3���3��3�d�3,�3y��363B��3x�4���3f��3Ȋ@3)�3�e�3��3�I�3��U3�^�3uU�3$�3`��3Rg:3g>3Gl49)�3M=�3gݽ3��3Սi3W��3��3�@�3I՘3���3�r�3%K�3\�3��3Kz�3Uʙ3i�3��m3��z3w�,3-�4ۏ�3)ֿ3x�V3�R4��3�s3%��3�ι3�3�p�3���3y�l3�[�3�i�3e�3H�3h�;3���3K�4�ׅ3G�3��3_K$4��L3�*�3��3��3w�3۫�4��3P4���3Juv3���3��34�4(��3gY�3�W4��3�{4cR�3v{3Ίe3S0<3��3AQ3"�A4#��3Ɖ34�b3�`�3V� 34�J3eZ3�#3��`3l�-3��2jLO3$�3y
3ڐ�3�{3f�3��3�32��3vy3P�2hP;3�K3�U3��C3�z�3��W3��_3���3�&�3��<3�@3���2x�3YI�3��3���3�F3�PP3$��3LK3V�n3��E3� `35�3}@3F�3��3�$�3xa^3��3��@3ݵ`3��,3S�3O�:3��3f�3��>3ʣ�3^�e3(��3��
3:&D3<g�3B��3�_23w�
3U�m3;3�3��&3���3�)3��3���21 !32�,3��>3�X3�|
4!#a3s�Q3�43���2�q32�3�׀3�\�2��3���3�\q3�Ȍ3SG�2���3�uf3 �3-53,�33��3�3�v�3
o�3 -3��J3�^m3�153~�2$'�3�l3k�3l#�3��I3c�32�E3�3��_3��?3�U�2b��3��e36 3/H�3;_!3�\3Ǜ3� �3��g3��M3-J3��	4X�-3���3a3�2��|3�|3+�3Ot3�)�2��53��l3mS�3W�3�-3OC3�8w3�35��3�33b3�|W3�s�3e+Z3�<*33��2S4��2c113^�g3Q�3�cR3�}�3 �n3u�2��3$��3�L3�Bh3n�3)?33��J3e�2)a3]�3O��33$j3��3��3�3n|03���37�(3.�3x��2�3�o�20[]3�I63]�2��3�<�3y63q`�2kɿ2~3�G3�k�2�*W3Y�/3؂3��3��3��3��3��2.4Ǖ3d�53{�A3DH�2�:3qzv3J�23��\3#73��3���3> u3��-3/DF3�l43��E3�`3R�!3'z�3�3b�3!�3�3��3�4���24�[3b3z��2��2�k3�BO392$3�W�3���3�fE3�3�6�2��X3�G<3��3�q�3�\�2�Ð3�:?3�o�3f�53j(w3i�3}��3�|3!�Q3-�M3pӼ3��3�1�3��3O963��3���3v�3;��3W�W3�)�3�<�33�A\3���3:��3��>3j��3ӝ�3�C3�Ƿ3��3�PD31�3GOI3�1O3���3��H3H��3�[�3p[�3m��3.d�3v�3�E(3���3�3K;t3��r3Ў93n�S3�(3QZ�3|,3%y3�_T3$
4�Gv3�3jE�3Q��3�Ԙ3�\[3o��3X�3��|3I��3J��3\�r3ns�2��3���3�y3Bl�38IE3߇�3=xW3T��3^�|3��3Jń3�	4�x�3�q3-�3��3ot�3#c�3z��3�b83ɣ�3���3Ơ�3g|3��3DU�3O�3&5m3��3�[3���3nS3@B�3/��3�533t4��3��+3��f3Φ�3P�03��4Zn�3;V3��3Ǿ3w��3�M\3%�W3��C3.��3_�m3T�3N+�3���3`.!3�	�3(�3��83oQ	4�!4�c�3�ɍ3�ڱ3�|�3���3�`=38"�3e6e3P��3=�4M��3v��3�S�3�vS3�3��#3^qp3G�e3焺3�I�3��e3ï3�qS3��3{�47l3��p3�e3�V|3G��3H�53��376�3��{3��"4ۘ3e�W3hq3�S�3�R�38�H3М�3�3�ӕ3n�R3ב�3��s3ڔ'3�i36$T4��\3���3�n13�ne3��23w��3 EH3��_3k:�3Q�3��3j."3��2�%t3�ҟ3�F3X<�3$M63h��3�3�g�3��o3�3�,a3a934৞3KΚ3���3�!�3��:3�T�3$r�3MP63�fT3�,4�m3�r3�'3^d;3�3���3�s�3]5W3(��3#\34��3>9�3��:3Œ#3�'4���3���3��3!/�3O�}3�ڄ3�%�3�3��l3���3�r4���3��r3���3�Q�3S�13�(�3�2��3�K3i��3�aS36��3�7W3� 4b�3R�3���31��3�3��4߅�3A��3C��3&� 4���3�n�382m3*�4��3~TR3Uw�3C�3�94ePq3���3���3� 4�u�3�Ql4fө3���3E״3M�4�4�3�"4���3m��3�4�3�#4�04r�c3U�3��4Rd�3��3gO�3<�3��4���3�"4��3ޱ�3G	�3�p4W+�36m�35��3��3ys�3���3���3�'4yt4��x4��3�c�3�|:3�!;4C�M4�3!%�3��3� �3�3�3%^4�$�3^�3{k�3o�74��3i�3��4�54ѣ3N�4c�4�K13� 4��4��34��3�E�31{4�3��3�3��3F�4~��3��3A�3֌�3�4�(4g�	4��3�4���3�$�3�4+�4
S.3�i4��+44OO4�/4<�3��4W��3B�3��3���3$�	4VZ�3JL4�4~�4B�L3�@:4.�3Y#4O�3�3�37G�3Ě�33þ3|�q3Ǳ�3E�4�m�3dL�3��3��L4]�3:,3�3 �3��4Yb�3i�A4*ˡ3P�4�
4ׄ4�;Y3+�4*B�3�)�3�B�38`(4N
4㩆3v54�<4�u45�24���3���3�3��3���38�3�,�3]z�3��4�/�3J��3w{�3{'4�ճ334���3ۡ3=�3��3�(�3j��3|�G4k4C9'4`��4��u3Ց�34�2�3 �4�۶3�$�3m4V��3r4h��3���30ؔ4k��3�[�3�*4�O�3�]�3���3��4t�M3��4$�48�4qG�3/��3h�3�o4���3M$�3:��3�D4��3o�4?��3�ƈ3��3Eқ42�3D��3E4�gR3#%�3ez�3ک3�X�3��4��4��3���3Q>�3��3��3�_�3�D�39,?3�4��3���3��3?�2��3��93a��2���2G(�2a��2��2���2^�-3&�3��2ڞ3�+3,�2���2t$)3��2�!�2(ʞ2�3�3y7�2�(A3 �+3�b�2.�2}`3�J*3�=)3�$3ZB�2e��2�3�K3d��2��2��z3��O3r�K3�V�2�83?c3�K*3'�R3ޣ�2SH3��2H�;3��3}��28,�2��K3I��2��2U�3�3�a�2�3��3��3y�3��3�[3�P3���2���2_|O3㓷233ƹ3B3:S�2tC3(u3�3>�2�p3�[�2��3>'3\�%3�G�2%z�2���2p�2ʧ#3Ѝ43r-30A13���2�\ 3��3�e�2o 3=��2�A3�@�2X�G3��2�)3SC�2�}�38��2|��2�N�2�Ғ2]3��3�p3K�3Gf�2� w3�3��3ϓ�2��D3�/3'Z�2�ڇ3'�31��2�i(3aC31: 3?043^^�2��&3�w3a��2�6�2��
3�Q�2���2��
3�L�2P��2S�f3�%	3��2�`�2�N'3��3-�3���2��3���2���2��3�M�2,q�2�3���3|Ž2���2��2�O�2 ��2��2F�2,Y�2�v�2ar3��3w+�2F��2;3$3�3��22<J3��2U�33Fz�2��3*3�2}k�27"	3M�3�23�b%3�B3��03��
3�3�<3\��2�H�2��h3�Ϸ22U3Rh2��2�
3��3�|�2�˥2q3o�2��3�s�2G�2PD3:<�3S�2���2� �2�ѩ2F�2U�3J�2��2�U�2#�f3�t/3���2�^2~N�2}3��3��2���2;3���21p3��2T+�2���2�wa3�>�2W��2���2G�2��2k3���2���2���2�"3�.�29�&39��2\�3\Y�2߰�2W\3;/�2=��3��2G4�2��2��3Uq*3X׹3��,3�H33�3�ȋ3���2�D83`3̽3��-3M��3��r3:Y=3�Z	3���3��@3��z35��3��>3�Xu3&�38h�3��>3\f3��3���3�3�t3��f3?�K3ZoY3�63�0^3<[<3��\3��3��3��_3'�3���3s�E3��3�(3�#3u�3A/O3��c3F�?3��3�!F3��3 q3��-3�i)3��3�3o� 3Ʋq3�3�>L3�Ȇ3��-3�v�2s3�Nm3D�c3��2�k830[3);3�`�2��p3�N3��:3��93�D�3�B3=�3�!3��$3�u3�%3�nH3�E3��E3�,o3�;3l]M3]ܷ2���2�Bj3n�-3s�.3�d;3q1�3Z�3h�|3S�3��3�Z(3�1�3h�K3F�x36|3߹#3�)$3��3��J3�f43uN3���3�À3m�3���2�i3q�2��M3Y�3\�3�K3�43�<�3C�*3s�3�LI3�4{.>3Ch�3p�?3�O=3.W3f�/3�l�3	)g28�83u�C3��3&V3c��2�3��B3��o3$�33
	�2N��3ǻR3`]i3�ޝ3'q3ܭ�2���3,;.3�<3��@3�$)3�g3��3�Q3`�3���3!HY3�O�3�i3o�-3���3;L�3�@g3<[3#�2�NP3���2�Jy3��83��3H�j3h@�3�&�2d73��63�z3�e�2S�?3�WJ3�83�X3Mc�3���3��H3��2��e3͓H3fh�2]�33�:�37�]3�D?3�y3��\3��a3;	4L�3Wk3e�T3��03o�3�^30�:3��2#�E3:�3�3���3��63��f3�S3�h3�I&37�:3ʍ�3��\3�V�3�*3��2n��2�.�3:�2��293�2|�3�43R�3�(�2Ѐ�3���3H!3�
3wǚ2�~�3 S�2'�2K3��2�Z�2` 3}�3��&3��738?�2��3+�3ˋT3�I3I@(3�
3��36�=3'�2=X"3ˈB32� 3��T3�x�2�K&3�,	3d��2�13�1\3ע�3s*�2�sx3��33��2mx3:y�3H�T3��?3J�230�'3��C3	s3��P3wX3�VS3�+�3��[3��e3���2��3	K-3X�3'3.�J3�?3ӄ"3\ɫ3'�d3[u3)03�,�3�p�2�u3��63�g3|^�2�y.3���3Y"+3b?	3� c3�u!3I�3Q.3�jZ3��?3��'3�.=3.�2R3s3f;&3ά@3��:3��83��'3�u�3i�E3�3��:3�3,�T3�23m�i3��P3F"a3�Qc3��@3�7.3a��2Sp3��3`T3=1@3�3��m3�F�2b8N3�3J��2�N3~�3ˡH3�#3�3յ3~�)3z��20$f3��i3Id�2��3,�$3b�,3��2!�z3��3�I3[<3SwR3�23m�Q3��3C"+3��3��2N}�3�g3��U3�#�3o�x3�`j3|3�="3��b3!�03�+�3��Z3ࠀ3W3Y3oJ[3��*3�3�e
3[�3���2W�<3U��3H�3:��2�)4r��3�AM3W�34�3��13��o3ki>3ˬ^3�|53M73��Q3�!3��2��?37]3�$`3W�E3&ӿ2�jR3�!L3m	S3�C\3>sC3gG&3���3>Q3a�3k�3G�`3@%�2�mJ3��Z3���2|Yc3���3--3r�M3�'�2�3U3tz�2��B3%�C3�p3���24FK3Wx3��J3�w�2�F�3��3��s33��3H;�2�u3v�U3yŇ3Yhm3�ȗ32\y3F1:3_{�2��I31kW3�D/3�33��2��3&��2�[?3�e83��	3��22��3*3<`"3@>3�03D�3��>3W%�3+��2��3���3Z m3�f+3$��2�C3�E13��3�s3��2��3���2�mE3�GH3���3��O37�3�Yk3��$3h23� 3�36CQ3��z3�T�3�pU3K4�mb3��$3�^u3���3h�(3��3��>3�=�3x�
3 y�2�g�3m�f3�3�z3c˟3�CQ3���3yC=3���3�]B3�1s3[��3��3��-3F�c3�"�3���3�3�e�3je3���3�K\3I�C3�t3�aN3*��3"��3�lf3�(3���3ˍ�3��13�Ԙ3��3�G�2sC3��3��3�My3.�4N��2433]�$3kK�3��23��3��D3?�3�G3�U�2�E�3�`39\P3�J3Ho�3%\31h3LIv3^�Q3�(3~#.3h�2n3���3��32N�3� |3���2�-)3ŴR3�jQ3R�]3�A3]t3�?A3/�|3j�B32�K3�d�2'��3��3�W3�u!3��3�֚3%=Q3G��3ʵ+3f��2��3n��36�3�R�2�[�3i�P3 �23�73+hC3���3ά�3���3�B^3���3�lu3W4�3�3���3$5�3Z�3�w*3�+3��3��3�(3д3T�33>�S3�?�3��3�s�2�~�3.��2ͧ3��3hE32�A3;:m3��;3���3'H+3��3P�53�e(3��p3~>t3�W�3Z�3��13���3�&�3�3$]3���3hv�3qC3��W3�@3z��35�z3���3 �n3���2�W�3�e4�;'3>}q3(�u3Z��3�|53А3��3��E3���3�4�3C�3mt�3RC3	�F3p��3f�3VL3�37�k3�q3M�3�/03f.^3�id3�Ϊ3�
3y��3D3"��3c�2�@3Syp3��=3Xx3i(�3��3�4E3kF3r�3H3��P3�g3!Q%3k�\3R"3���3���3^��3��3�64��2��3���3V]D3���3q3�@_3�<�28]=3l�O3_�3r�u3���2ꀃ3EF~3DP3���3X�2q>�3�J3��3(8~3���3�Kq3?�4��g3���3Z�`3�H3*�&3��3 X3�"3�o3--4"�3E�R3�!3�O�3��63�^�2��T3h�t3�\�3�g3|4yI�3�� 3��3[4Иh3W��3�Z�3���3o4HI�3[�3�}�3EF�3��4��3���3�F3�&�3�3JF3U�P3��=3Z}�3�W-3#]�33�1�38y�3���3�k�3�Y�3L��3��3�R3�-b3�.�3�m3m�344�C�3��3Br$3[1�3��i3
�u3�z�3��3�ݮ3/\t3s��3��3��~3��3ÿ3/�/30��3oX�3�׼3��m3Ѵ_3���3=63H6g3s�4	|�3RЈ3�>3E�3$�3W�D3��3�_3��38fR3JY�3�_x3�&�3t��3|�)4_7�3ն,3���3G�r3�Y�3�N3�H�3q�3+�3	U%4�b�3v\�3G?v3G��3�-�3��3��E3�>J3o��3��3l��31l=3j��3�˹3_4C�W3��i3Z`t3�g[3���3د#3�|3W3n�3$��3p�~3���3!��35��3���3�3��3��3:*�3��C3Y�3�L�3v��3�6�3�r4��3�3m�3 ��3r{�3�3�}3�WO3E��3Δ(4�]�3�z3��r3I{3w��3vy3v�3���2s�l3�Q3>}3�H�3�A36�3]�;48T3�N�3��$3k�3
aR3΍�3�,�3�%3�7M3%r�3S�3�0U3��+3��3��s3�G3�n3�_3m-3���3-Q�3%(#3k��3N��3��+4Hf3ȋ|3bZ�3dFU3�Uq3Aj�3�J�3oJ3�S�3�4���3��3��W3w/�3�3q�93�c�3f�73&��3|33c4��3��W3��3��_4^�63��3��3�1�3��h3-��3hG�3I�G3��3sF4���3�r�32�3?�3>��3Đm3Wˈ3q�)3�"�3ΞI3���3N�3�X{3���3���3�843ʢ3n6�2ų�3jF�2�I3�&3�|3�`3��b3��3�3�3�2\j3��.3�Ĉ2Tƞ2�>@3�~3P��2S��3���2��2L��2�J3���2�|A30�3�(3BB�26+33ל23'I2��3th3ZA38��2?j�2�V3�3�*�2�/3xq:3�G#3�M�2+`�3P�E3��2HG�2	<�3�J3i��2em	3f83�c#3�Y3o@�2WB�2�>35�f3�H3�� 3>s2(0�2�Q3�3K�13�p�2�|3L33��(35M�2~V�3&��2o;3I��2��A3K93 �73�� 3\�2��h3���2�y:3d�3�(3E"3	\�2�3D3u��2m�73@�2��p3���2H��3q�?3�3؋3l=�3)�O3,�U3�3}3��B3�	$3C�`3�k�3.�3q
3�IA3C��3�S3wH;2��_3��3w�3��3��u2�3j�83>�;3��=3��33�!S3)*{3^�`3p��2 �3��39S(3b)3��2&3�3n[�31�Y3�~3�$3��h3g�3�̥2h�2X��2�h.3S9U3�M<3��$3(3�%3��3��3��a3�	_3��2�}O3tC�3K!332�	3��2��3}ƒ3��@3e��2p�53�T�3��38: 3Gm�2{�+3��3wkI3B�3���2��P3��3��2�"3�̸2Xj3��H2�d3�AP3���2�e-3e�G3�3=@3���2bK[3��3 �
37n
3C�t3i��3���2L�3h��2.��2��13s�V3� 3K,B3*g�2�3]�2�3V�3};3�3"3dC3Nm3 .�2��2/>�2#�3�A	3'�3��2�=3س�2�P�27�+3��`2<�2U�3<��2l�2*3+3�H�2A�2T�!3/��2U�/3�
3��L3C�2��2wk3L�3Z��2`�#3�j�2�-3�8 3 �3���2��3���2H�h3�#3��Y3���28`B3xV�2�8-3���2�U@3��3�_53'>"3� *3	o�2���2j�J3�-�2��3�A 3�~�2�3�2�vW3U�23��3f��2z�3E7	3s�i3^�3Ws13):&3H��3v�43��2��N3qr�3��3�4C3+�2'Oa3D�c3��3+� 3���2��3�%3y"]3./3�E�2�+�2�Q�3�T^3_63�I3m�83�F3�f)3c�3��3=L3�Q�3���3<M3fַ2w�r3wA53���2;A3�>�2�JC3�U#3O��3�x�3��3볙3 *�3:�L3�j3�a33e�53j�%3�rG3�bI3���2k�I3��3�8�3��C3;�J3�P#3o�131��2�`3��53/�63�/3�Zz3E!3|�3�$3�_}3���2��2!�3[�2��"3hYi3]�J3!�3y�83�E�3�t3��2�	35�}3�03/�3�m3�*
3+��3"�2(Ȁ3Q�@3�3 �3R?�3��2	W/3��!3���2��3���2{�2��2>�$3��3d�3�pS3"��2��63��3�b93��3�}�2y�+3p�)3d�V3D� 3s�a3�=!3�4�43)73�|h3
�S3��*3���2��{3��2��"3町3��?3`�@3���2��F3j�?3$}3�3{l�2=�63���25Λ3z�3�c3m��2��4�\Y3�s3�2.31�B3��3]na3��_3h��2y��2��37�3�O3�35z*3
)$3�93jGs3{��2�v�3���2L7o3]gM3m��2^}|3N��3
�3�d%3VX	34 #3s\3��U3�a&3���2��2w�P3<�h3r#E3���2��;3�3��3�F'3�2{M3���2�RI3�t'353k93!��3�3>e.3l�R3�?_3|\�2"&3�˖3 ��2��3��3��3
*3"p(326A39�u33G�3Z��2͜<3���2�8�3��(3�k4Zi�2��3��3Nd�3�3fխ3�3���3�8�3�	n3Dl�3�24ri`3T(3x��31#�3�܋3�d23l6j3qB�3h O3j3�}�3��93�3�3R^�3T�24EE236�83<�\3��s3���3ƞ3���3�[�3^-�3|c�3�_�3;�3�� 3T)�3�K3+�3�o3��3�n3܇;3:��3�H�3��_30�3�}<4J�!3π3�݌3���3�H3�ro3�k�3.K3`2Y3�_�3���3�<3D"3<EB3#��36==3�<�34�L3�'�3�3�g�3��3� 4��V3�$4���3��3�ӎ3�P�3>3��53�B�3�&3:��3��4wܼ3P�3	Np3�T�3�j3Xo3n�3��e30�3^D3���3:g3P3y1.3�4?&H3Z��3lz�3=�>3MU93�w%3��3"13�ā33�3p�3��3�/<3�Z�3��3;�g3a�3i�K3�-�3���3��a3��3��W3q�83b4^33�k3��O3��3�@�3޺�3�P+3�v3�4��3 4���21��3aY�3��D3�'�3��d3�$�3��R3�i�3�2i3T�i3�7G3�a4?�>3��3d'�3�M�3�x�3�2n3�ǃ3=3���3hS�3��48?�36zU3j4��{3N(3���3��-3�ܡ3[Ѽ3x��3ΈZ3���3��53�j	4�Q35��3��3��/38��3�3��3��3N��38�
4e��3 R�3��'3%��3{	�3@3���3�>3��3�
3'4��3�ub3�z3|�4�߁3,�w3��t3�Ga3��B3��Q3/[�3t�3���3���3u�3�
�3��=3Y"�3\6�3+��3'H�3M@Y3�R�3n�\3H< 4�L�3|�3�03�4ug3V-�3���3�B�3�oU3��[3�4�3��O3�4<_�3��4TB�3Q�3#��3��3���3��o3ٕ�25��3SD3�߆3l�4�U�3u}3sÈ31;�3-D|3��d3��3�u,3��3�P�3�y�3�Z�3���3��D323c3�g3��3�x_3�3|n73̋Z3��3I�)3���3�d�3��3dW�3�rN4{�L3>�93��3�δ3�V�3T��3G��3��2C�63&v14$�3�S\3ת3�%3�Ti387�3|13�<a3�ؠ3��3|�3��3K�]3�3x��3^�}3>��3�x�3a��3�&3�Z�3t��3I(C3�Ro3l��3'6�3A�C3ĉ3���3�;�3��83}��3��Z3���3Y�R3|��3�n�3��N3l;�3$#4)[43`3�**3z4�3R O3�k{3>�L3Yc37�13�Q�3E��3��3�� 3���3,~�3]ve3Jl�3�0�2�ˎ3	�j3���3wŕ3�?[3f\3!4�l�3�
�3�-{3<sI3��3��3�pV3`i"3�M�3���3��743-`3W.�2��3T�3��[3:"3<�=3*�3��B3��3�Ѵ3ׂt3�^�3��Y4�U3��3#b3��}3^��3a�E3���3��2���3�{�3�f�3#.�3�L�2�3�3V�3#GM3��3Z��35��3���3�E�3�P3���3�ۇ3cq>4=�3l��3�Ө3]��3Ҙ�3�!�3ь3�e+3�ѩ3�44�3Sƈ3�γ3�v4.C�3>�g3���3�3ڑ�3$�3�V�3��3!��3eDj3L>4��3Ҏk3���3��3ЋL3ǈ�33ky]3�x3�л3��3�7�3�T3��3�93GqS3��3D3{��3c3�64�n�3�53��N3��4�3���3���3~�]3��D3�(3�B83(O3�a3�"�3Uٴ3���3�	3~�3/�4�g�3�w�3:#3�|�3��|3���3��32e�3��%3�K�3|V53��`3�4s3A�3���2kw�3���3�3�8�3.
4 �3F��3��K3k��3���3��3��3{�B3b�3�F�2��34+�3y�4�,�3�4�'�3�{3��j3��4�Ku3�U�3��247��3�3���3RY�3��4�n3&��3���3H�v3���3��3hG�3\L3�f�3iQ4_NF3���3��4툛3ح3��u3c�3� 3��3���3�3SBw32�D4^�4&s}34TS3���3���36�3Ǝ�3h_�3�3�3�h3#_�3���3%��3�%Q3;�&4Lu�3�+�3�Ų3�N3ex�3	m�3���3�G3]��3:�E49�3u�3�w3~O�3�Z�3�ώ39��3b�3���3��3X�3Wm�3�� 4�L�3�54D�3���3V�3`_�34K�3;K�3�d�3��3�4��4��3���3��*3�4��3�H�3T��3Ui|3��4��^3�e3�f�3�o3��:3��:4p=o3�J�3�by37:�3Ma�3\)�3R��3��30P�3��04���3�'�36��3A��3	�3߭�3�S3��3�J�3$D3\=�3���3o8>3}�Z3 �@4.4z��3-z�3yS�3ĺ�3c*�3�I�3�;�351�3;@Y4���3܎�3�s3>�!4=��3�(z3�)�3�UZ3��3���3c��3�d�3yѶ3��P3@�3=e3�b4=��3���3���3,	4;\[3�)V3�ǉ3�_14@m�3�e�3� d3���3��w3�?�3#54�~3��3@<�3Ú�3`��3'T�38��3��W4yD3��3�)�3b�k3HhT3}��3��3c��3̏�3-4�Ѻ3��3Cz�3��3k��3�503�t�3� �3o�3�\3�>4��3�:�3�oj3AqM4�e�3���3� �3nt�35�@3PJE3J�3[�F3��k3B84\�4E��3x3���3ڃ4�TC3���3�z3���3'D�3M�(4$:�3�83�w3��j4�@�3�A�3�M�3�:�38R�3��3�q�3NRC3��4���3�X4g��3n7F3�Q�3��3_��3",�3��h3��4׾3G��3<|41&u3W^343ei�3�0L3�)J3��[3b�i3�4\3�@?3^�636�A3��3DIS3�A83w[I3��s3;�:3�3Z��2�a 3��3×3���3|0o3�3��[3�m�3�L;3�~S3�!3|��3�4�29�3&��3�*�2��J3���3Za_3�3�Y3�A3��2�Z33�K3�,3��n3��3��3�Y#3Փ�3�*3�e�3	��2��F3��^3qDe3.��2˅3���3�A3��I3^��3a�3�53�83G�73՞F3�4�2�f3��2��38�K3F�3ǘ3��i3Z�-3��*4C�3�63ZI3\�i3�	38�3cˀ3�a�2�$p3�/�3^|3e}3Ag�2�F3i��3׀�2339+3vE�3�3��r3�Z3��(3%@�2N*�3�WN3�=3rR3��2�Y%3rKe3|r�3~:}3�-�3�+�3�h3�/3X:�2�t3d�w3��=3��J3O�(3�]?3��3���3rϘ3^�301�2�&�3D3�M13�ň3ı+3�v/3j��2h�j3�3V�53�F�3~�^3VH(3��3o4.3���3�w�2]�g3\353O,�2�=3Q�c3��&3Y�3��3�Q3y�@3�f430ˀ3Y v3 ?38'�3��G39di3!�3v��3��43+M�2��33|�f3�3+[3�Z32}�3Nl/3+�3��%3^ 3ѥ3
�3��3Vt3=3ޡF3O3�҆3;�3�u43X��3��3p�z3�#3T��27fd3�3^��2�e�3�H�2��K3Z�3)Bn3�J3w~T3���3k̼3�>3+��3��c3�c�3:�J3�f=3b�P3��383=��3σ�33s_3��Y3�>K3!Y3�=b3W8�2 #�3���2&BN33�"303��2�܋3��\3�:3.�53V�>3�33D�!3p|J3���2TyC3�3`Z�3@b[3r\�2�ۄ3�\31�U3�3�U�2|q3o��2y�3.3�H�3��K3d
84#.c3:�3�P3�@93��3�3o@3�)3+Gj3���3zsX3��3f�a3���3��.3���2�1,3ai�3�U�3p=r3_��3Q�3ހA3l��3�,�3O�R3߰_3��3���3>�;3gD53��3<<?3%fV3��3 ��3'�3
�2(�383�Hv3Y=�3��X31��3,�t3��3;��3o:�3�A�3�&U401E3�u3x`)3�R�3%z"34=�3�$�3s�K3��3�x�3jè3K�3�^�3�}J3�?�3��3�S3��C3{��3ۻ3�L�3�v�3��g3���3bm�3�ނ3~Ie34W3�;\3f]<3gm3~�3�[3%�`3���3|��3�B�3�Z�2/�3=�33��3Հ3CF�3<��3J?)3���3���3h� 3��3Z�R4p�S3�#�3�[�3x]�3���3J�3�}3F�03��q3��3���3Ju�3SN?3���3L3�3�x�2b��3MC�3�3V �3M��3}��3K3�X3��/4[��3͓�3��3 wI3j9�3�+�3��H3w�3\4�3+��3�o�35��3Pwy3x�k3���3ݠc3��3,sH3BvE3��3S}�3	{3��3�<3�94��3R͒3q��3J�3ib�3O��3ZŦ3d�$3�3��3
�3��b3�]c3���3P�3��3���3�">3��e3�TX3�@�3GK�3�N3�ލ3��14p�)3�&S3z�3��3m N3M�^3��y33�3s��3 �3��3M3�G3s"�3[�t3��Q3�x�3�Xo3�H�3Pv3c��3O�3fo,3�1^3�(4&5�3�wh3zr}3��3�{�3B�-3rH73W�$3O�3��3W,�3��p3M��3=�I3Oc�3ڄ�3�?3���23D�3�a[3vN�3dm3�{-3)�3�249�&3!z�3�+�3�gY3_}a3���3���3�i�2�\�3@��3��4	��3��3���3��3y'l3��3�<3c�]3�,�2O�3p£3��`3!73�^H3�M3��3]�3��3>��27\3(�3f3��&3'e3)93�#3��2r�/3�on3BZ�2��3ø.3j�@3���2�23�w�3��G3�R�3��y3��3���3�2\3}�+3F�L3b�:3Z=�3���2��3rO3�P3���2�Py3�U@3�'v3��>3+��2���2E63�K3ڻ�3wi3l��2��3J )3'$?3�|B3��3���2�&y3/�43�c3�G#3�O�3s��3v�3cM�2g/A30��3�3��M3Y3(�>3y�3lk3�/3s�G3�	3�N�321�2�V3i�3"�3<v3��%3�'�3;��2��H3s�3JU3B�3�:�2��83�3 ��2}�E3�I+3��3J'3��\3a;�2\�,3��>3��3[m33&�H3_SY3�23u�2��B3�-)3 ��2%_$3)Z�3g�3�>&3��O3��c3��J3W�3�%�3�Z3�b3�3�N3��2�3��03���3ݣ3��2o�23�%3Ү'3gn53�13��2=mu3��3:g3_�#3+\�22�3�j3��2b�3�03ܼV3��&3�̃3��73M�"3��2i_�3V��2U3L3�W3)�73��231�3��$3��436�3�i3@��3�83;��2�p3��2-2�2��w3˘�2@�;3���2���3��33�n3#�A3 ��3 �-3�E3��3h39�B3D�w3U�m3</%3�*;3[�}3�ޙ3��w3�H3b)T3��!3z
�2z[�3��2�4&3s��2�j3��83��#3��=3��4��3��E3�J3�,�3}t<3T�2�YH3߃�2�C:3x�3�І3:�J3 3��2���3/�2Q�~3d73�h�3�3��A3}�j3�3�2\+�2[��3�T 3��>3���2qu23[�3��2_��2�q�2;Ϙ38]�3dEZ3�D<3�ކ2�83��N3��73�L53�Q38�43��/3��3J(3(H�3�53-w�3R�63�13�<�2u5�3mg�2�Q�3aG313x�`3T�3�433�-63�3t�3�F3��3��3"�T3�3���2	�3`3LY�3���3K$�3t�F3��83T�3��3�I�3J��3�N�3դ�3@Т3�`3
_4(r�3ĉ�2���3=��3�33��3FD3��93S8
3�S�3Vu3�&m3h-3f��3{�43�T~3�%3�D�3��f3�-�3��k3A3�Ǐ3�gU4��3"�93�M�2x.�3�d3���2�ht3F�U3 :�3W3�4a�F38\m3x�U3û�3|��2+V3ë3}\3|>3$�3裣3})�2&E�3e�3�|3X&M3��+3��3�W*3��G3Ք 3��$3L&�3�&�2�3!ʓ3��3�
53�3�3oxe3 �3�\3U3ё:3DVN3�31�73N%o3��3寤3ΑL3��53��3�Ջ3Gn;38��3T<]3T4�3�4�3_33(�Q3<@43wۓ3���3��3֎�3Dn43���3���2�ǐ3ڏs3��2E$S3)�3���3Ě�3:�53�E3v�E3�f53p|3���2�M�3NX3�}n3q�3��Q3��2�R(4�C�3�� 3�3943A�3�~3L�x3�?3k��3Ϝ�3��3S9<3w�43Y��3�g�35�3��3�.3|Dt3$53ץ�3�ic3t�3[C3�4�B636 3�l3y�&3ԧ>3�\M3��i3V�3��3%��3�5�3�a�3��F3DZj3��3}�3�#r3U;3�;3�=3��3�Z3Taq3�I=3�4i33��Y3w�3��o3�;3�-�3�"�3�"l3_�j3AY 4��3 a3)3^Rs3	r3:tE3��^3�-37�3iz?3�L�3ش�3�:3� Q3)?�3C��2��3�|3��Z3�Y 3�	:3?|�3-,3ox3�3�3}�3��S3�#�2d%X3 V3��)3��13��2}У3c3Y>�3�o]3]A�3-{y31�3�F�3?��3��L3�{�3\8_3�Vl3�04�:�3Pg�3�u�3�]�3L��3�U�3���3_��3�Q3iyQ3�:3�(�3��3F943��3�z3�(�30l�3��3妇3Lѐ3�Ӧ3kS3'�3��3�H3k��3�4���3���3p�3B��3)W�3߈63Dι3-m�3�U�3@�3`A�3v��33�3�Ƃ3��4�E3�F�3ieN3^��3��]3e��3;2�3hB�3 d334�3��3�-L3���3�]�38�_3*��3Q73�	4�3U�Q3v3�3�;3FW41��3���3�3�F�2��#3i��3�#�3Z�(3�&�3K�4%l�3O#3��3�.�3�ؙ3�c�3K4.��3HϪ3r\43`��3��3ɋz3���3݊�3��3A9�3mϸ39*�3�[y3��3^̘3m�13{3���3ԏD4�MI35�-3@ǡ3x84r�83@r3U�35��3�	3���3H��3��J3�xc3��4�܌3�&�3�g]3`�3�V�3a��3�3��93�"�3E��3�r�3G3N�83\��3<�3�-3��3�rT3��3�ʘ3
5j3� `3_�3=�O3�A4k�3�0�3|�3��3� �3ȼx3���3K�[3�U�3Qr�3� �3�!_3(� 3yz�3CY3fAP3�	�3��C3���3C1�3#�3�z�3��3￲3T�-4�L�3(��3�JY3�T�3�Q�3p�N3�2�3{q,3�|3�%4j�*4��33E�2۳�39I�3S3���3H�3|(�3�y3�?�3�`w3Fn3T<�3k��3���3m~�3���3��83.zo3V*�3׭�3o13�Q�3�K.4_G�3S��3��3[�3cǚ37[�3Oˏ3�V�3��3ð�3�f44��3z�3jB�3�o�3��e3�<�3��3��y3Q:w3�6�3��3_�)3�4���3�
�3��3�n43���3��3��73.6�3��s3%��3� 3b%�3�χ3��p3��3�w�33^30^w3���28O3أ�2��p3��i3�;P3�� 3���30�83673Lc�2|�3��$3���2�v838�23��k3�43�{�3�'3��3PAO3Փm3�)3�S3+�\3��3�33��3��@3�ۉ32�3�;�3w �3�z3�G3���3	3�I
3��<3�2��3�"3��3�$3B13(��2���3�V
3� �2�3��3b��2��B3�&p3\\3YeC3�q�3C�3-3M3�\3��3��2��G3*D3S͋3�
c3�*`3��J3� 3��+39!�3��3�Z3R]3�|3  f3�4<3`�3��373� �3�3�%3��27�3��D3Д 3<�3���2�pH3��n3�1�3��$3{h3�)3J��3�� 3[�L3o}3��P3�!3�:�3���3�P�2���2�t�3��H3#G-3=3��-3��43i~�2N\�3��3Z�v3�?23��w3!�3��x3���2���3֘3�3+�i3vrp3u�3�M3���3���2�p3T�3�d3Wk3�r3��z34d/3�C�2��3ȍ!3dQ3dJ3�Y�3��.3�F3��@3Z^�3�3�!L3���2�:S3:r�2�3�h=3g�3��(3��3z�=3C��2܀�2�wb3���2��23��3	��2]� 3���2��3
�3���2��3��35g43��&3�3 �3b+(3�A3�8H3܃3��b3Z�3�T3#�j3S��2��F3�813��&3�H�3�/�2��Z3!m3�=E3�8N3���2IQ�2�r�3��(3t�q35ET3fO3��3j�=3z1!3�o�2��$3K3`k�3cO3�3r2;�i3UK_3��t3�PU3^�2�G�3]�"3b?�3�B3	�2�E�2?)�3�BM3�A�2�+!3�23���2��2���3^�2}Nm3�t�3�S3aɗ3�Z>3��A3(�3���22Q3��(35�F3Cy3h�3��D38��2�{�2�;P3dF�2� 3�/�2�b�2֮2��53%3:�3�26�j3�o3�"3��35�O3�23���2vn83G3	�2b23jY3�w
3��t3x�P3�ϗ3�3�63DA3��e3ɾ3b�2w�J3tz�2F3�h3�3;A43�S.3��/3�1#3��:3z}3y�+3��3a3��g3�)63�i�2���2?~3�3�2�2v�<3���2N.3
�H3�,*3Ts73Mu$3r�83T�3ޅ3T��2��P3�!�2ˋ�2�*3�(3�g!3Y�	3��63i�2k03��2�@3�<�2,�3�޺2��2�,3%�34qT3fh�2�tz3�:�3��<3]��2�>�2��(3y<3���2�
3���2�.13��2uP�3���2 ��2�'�2_�[3'�E3���2�<y3���2`y�2���2�d�2g�21eq3��3@-;3�3x��2��3�	34�2�-�2���2��!3_3dp3sj3ٞ�21��2J�3!3��I3T%3;�3,)�2�=I3��P3HԱ2�A3I�x3ocv3�v3�y2Z�k31�=3P��2Z]3et�2SE3��3+�`3{1�2��"3�_�2"��3�Q3D�.3���2`�93�{I3mJ23�u3�}�2�0�2��g3�@L3���2T*�2�K?3�53��3o�%3�E2m�)3�� 3�T/3�3��2�c3�C�3�3s3��13�M�2��53�Gm3A;03ˑ�2�"3-b|3��]3�P3ܗ�2ޅL3d�"3�V�2�d:3!��2N�3ƈ�2Ż33
p�2,��2_X63M��3�~83gf&3t3f��2��2U3�iH3r�3�33#�A3�A3��3yޅ2��
3g�j3�3׏�3���2��2���2`m$3��"3~�2��3z&�3�k�2`��2%�3�n!3S��2�V3˄-3w��2>v*3ۢ�3�Fr3�*3I3��3b��2a��2;�D39�12�ce3"R�2! }3�3c��3zg3� 41]3#��3�3�f�3Y�83]
4q<�3Ɖ�3��3!��3���3Y��3NU�3p��3k�3lC3���3ZK4
�4�RT3qR4�z�3�%�3���3A&F4��3�C�3?4k4�3��3g��3E\�37�|36��3GR�3�P�3���3��3�4>��3�V�3|�3�Ǵ3!x�3�4���3���3}b�3���3��R4(7�3g3��3�S�3��s34v�3��3ZY3f�3W(@4�N�3u�[3��3��3���3��3�4p/l3C�4���3�4��3Y� 4��3&dY4[X�3���3A�Z3���3��3}�3�]�3i$f3Jڷ3��8454�r3<��3 �4a�d3���3{F�3ͭ�3��3-�Q3Ȭ4[�x3�!U3��3��D4ژ3�W�3]�3��}3ꇥ3��3d�4ˢ3~^4s�j4�4�ߏ3�$3�,4ڗ4���3�>�3ѕ�3sx�3�rm3ɲ$4{Ք3��3`x3D,H4�ì3O��3�4�{4�̛3|��3%��3ş4�H�3]�"4|�$496�3y�3�:�3���3��3^�3�S�3y�3\f�3��3bѲ3���3�L�3��o4�uB3½�3�i�3���3`�3���3�e 4��/39#�3{�4��3�)�3��3*�Q3��3�3���3Ţ�3�n�3�w3��4!��3L?3?0�3�Q4�3>=X3��Y3�*�3��3���3�N�3m'�3�{�3�K4���3�\�3u3B��3eV�348F3q�4�e�3�ܿ3S��3�04n�3C��3E�3�+84��3��3���3�� 30��3sO4z��3���3��3[4�R�3�{�3�N�3H$�3[�3?ȁ3%^�3�[36�X4V=�3U��3c3�v�3��2��
4H�3�\4�C�3�L�39��3Ԩ�3�-�3���3���3K1(4x8�3)��3Ѱ3�;�3���3��3��4��P3���3t�3SC�33T4�;�3hC�3�b�3��g3"�33�b353��|3� �3�W3?�D3#d3��y3gײ3w�3��u3�K�3�m�3�`3��K3a�93j3��3"��3m�3�S+3s�3�|�3�Ba3�F�3<�m3V�i3m�|3u�W3b��3s�q31�3��37��3~~�3�&3�|�3L��2�-3�H�3�q\3q^j3��p3���3v'}3V�{3��3Xd�3�K3,�3��2"D3svP3Z�O3���3t��2Nf;3Fj�3	�3#)3ݝ3H�}3 ��3�3"�H3�|p3��g3"+3�8�3�[&3�3mhv3Y,	4E03�s�3U"3i3�%<30/
37�3J�36�3���3��3��m3��3�*n3t�3���3o7^3��2Ӄ�3|I?3��3��a3�M+3fb�3�H�3�93r�q3�83�/;3�Ϭ3UG�3��3�,3�`?3`�3B/�3�R=3"�3�]�3f�3�A�2K�3�X.3Ş�3Dj-3Ydb3J�B3gWL3�a63��3EHA3A?N3�V31vb3[[3�O�3�4j3N�+3RD63��4�ʵ3]73��3���3�{73��!3XW�3B�3�34a3�?�3�M3�:t3T�<3���3l�>3��`3k��2L�43�ݎ3��3⏑3��3 �3G�4��3��l3�H3��3ܒ*3�53'C�3��3" �3^Kn3���3�31KY3BT�3�K4ˑ+3�3ʸ�3�u)3*g3��B3T��3�n�2��F3��3�̍3���3�)3[ʬ3T�j3��s3�U3��3\��2�X3���3+jp3#�X3r��2l�3�;d3N*]3�t�3�&f3�&3�Z3%-73o�3m�r3�3���3�J�3{|�2�v3/O�3k�Z3�zn3P3�/x3�23\W�3�73��23%�#3c�4�r\3��3U��3��3�3~{�3�V3�(3w��3!��3�4���3�n3�tU3=�3��3��3��,3��3<;3MXS32��3ݾ�3�Ҿ3��S4ci3�S�3aH�3���3�|3w��3Ꮅ3�x�3�2�3d��3D�3 i�3լr3Bf4E��3|�)3S��3e�^3�ǈ3S;3�k�3(�3\z3,�3��14a�o3��3£�3k!l3h;H3g+�3%�31�v3{ũ3a�4Y:�3�a	4|�D3e!�3t=�3J�3�}�3�`O37��3�p3/ �3g�n3>@�3{��31h�3]�!3$4�3�g�3���3M�3��z36�3�X3M��3�4��3A�}3�@a3Q��3ϸ�3��	3Ӱ�3�S3���3�<3��	4s*v3�^g3tn�3�'e4	:f3{�3�Y�3��{362�3	�3�I{3�3Vi�3O�L4��4���3��(3���3hJ�3��3֝3�4M3~��3�A�3i4(߆3/Й3=�f3d�/4;1�3?b391�3��w3�3� �3�4ֈ�3]!&4�+4��4H�[317O3�54-�4��-37��3Gͩ3;�3)j�3��4?>4�@�3+g�3Y�04�L�3l�4�t4�N�3�@�3�3e��3�W3D��3�[�3F�!4ơ3W��3)�3G�/4�F�3f��3	�>3y�3:�m3M�3�]�33z�3��3��4�`�3�\[3��z3��Z3�8�3�@c3EX�3�'q3�@�3��3��3�3�z�3V��3Eu�3��3iU`3>^M3��3E��3��3*�s3ĉ�3�"�3�
4�i�3%4�i�3���3���3���3K��3��3~1�3V��3�U�3���3��C3�l�3	;g3�9t3a�4Qs3sO�3p�3�e�3w��3,�3��31w4&�3<�3�L�3Y3��3VS4�.�3s�i3�ܫ3��3	�3Em�3�]J3���3_0�32�3��3c�"3%L�3�τ3��4Դ3& �3��N3�nl4�ɝ31u�3;C�3�Yj3;y�3uHi3X�4���3aΤ3��;4-zv3�'�3��.3xy�3I�|3E	�3���3�\@3�`4&A*3\��3�X�3��.3{(3�V3>��2$��2=�3�?3@ȹ2E�$3�~�2�#�2��2��b3��3��*3��2�P3�]3SM�2�03��2�w�2>K3ZN�3<;3�3��U3{��3v 3�W3��3ť�3��3��x3��?3Ų333��3�j3��l3��2YY3s�3���2��3��2`��2��*3LZ93��3�3ػ-37��3�ֻ2��3#�2�y3�Q�2���2�7�3�1�2�Q3.��3樄3�3=�2�*�3�U3�$3O3,�3YhB3��#3��K3��/3��c3�M-3�}�3a�3"�3xo3U�=35�2�{3ʕ*3AD35l3� �3�p`3y�c3.S3t��3��?3Ϋ2��(3w7$3�x.3�ǳ2�
�3���2#��27�3��3��F38)�2R�3*Ci3Nz�2�35Cy3p٣2y�	3nG�3�a3h_�2���2�6l3�3��2�i�2�ó2^E3���2��3��3�-13Fqa3�n�3���2EL<3��O39�3��2e�3^�2�3�.C3.�3���3̡;3�f3��3���3��F3�gM3��2�)31�3��2���2���2M��2���3u��2�@3�I3��"3�C3�C3��83��2^F*3`�n3t�P3a�13L��2�-�3��M3���2e�P3S�2��37w�2�%;3���2\³28��2Xv�3��	3�c�3���2���2|� 3��N3l,3}��2̓$3�l3A�3_�3߆�2?�3??(3�ո2<F(3�3X�33��2��;3��/3�n3���2�G�3�&3B1j3B=3���2���2A@�2p�\3}]�2.3�Ր3]'3?m3�2�B3�T3���2��F3ᵏ2Du33�v3o�3c��2"3���3�E3�S,3��{3�U�2ԇ�2�3o�3���2�3E�3U�3mq3�U�2[33�3-y�2e3WC�2��:3��2*�3�(3�T�3�?�3�e�3��i30B3]V�3髤3 �=34��38�3��o3��J3 ��3s^�3g�U3�K3v��3;�3(�F3:	53d�{3kb3~)r3ZG�3��3R�/3xQ�3(�3�@3���3��t3��3AĠ3|�3*�L3o:3L�W35��3���3���3��t2!Ī3KP33m��2)PS3LR3ːK3�3Ė�3�3��33M3�K�3.
\3��"3>��3�*D38V3f�N3��o3@�3���3�#�3ͺ4��3��Y3A�.39��3��M3�/�3�K73ȃY3�W:3!ݚ3�<w3 %3�6I3R45�M3F9^3��Q3�F�3,�\3Z��3Pd�3%=�20pB3�3U�3;T3Ш<3W��3e�3�:3��3"�`3}��3A,�3�9 4��=3��y3h�d3�u�3�k`3��3�M;3eh37/3�U�3_3�b3���3�4��i3X@�3��3F��3���3�|f3w��3B�'3�3��n3�+�3_83�V^3J�"3�X�3KlT3z3�C�3��v3�H3��3�s�3��73(�32��3�D�3o�]3>3躻39�3):3*+_3�A73�)�3ɂ3���3��T3Aq�3�83m��3'5�2hl3�y3��3�bA3M�3��c3��32p�3���3ϗ�3x�.3C3=�3U�3�Y�3͎�3N 3C��35(�2aͫ30UE3���3Gc3��)4�qh3eӑ3�B�3�f�3�b3&��3�3?Mz3$r3�J�3M�3��_3%<>3���3á�3�_3��3��3�t3�R#3jd�3%��3453�-3�0443��3i��3P=O3k�$3��v3��3N3�*�3<'�36�3�
�3V�Z3!�D3lg�3�|�3���3|3/3��3�|3�I3{o�3io�3߫.34�83���3��13f3�3i3n�3��3��3(��3i�3\-�3�QA3[]�3�S3y-3	n3&�A3���3/8
3�B�3b�R3$�3Z�j3�x3�T�2R�3
K�2��3�>�2��3<�3B��2i��2j5k3�%3	�h3��73�63�3%'3Z��2�Y3��E3��2>7�3��/3��3��v3Z�3��3�3��2GMA3X]�2QW3�% 3�I3L�2^�}3c<3�,3�6�2��3lR53H��24�3Qz<3f#]3)D�2t��3�A3�f3D��2s��3��2�23ф�2�z�3���2Z��2�73���2(�.3��3�B_3ѻ3n�2�3u*`3Oz3ٝ�2�3�2dd3�-�2�{[3���2Z^K3�`�2 ��3RS3�SZ3�
3�A3��2!?532�-3@Yf2��	3�_�3:Vl30 3��~2�n3!"(3���2o��2���2��_3CA�2���3�>�2��/3d`3��3�tl3P�!3ũ3\�3R)E3X3��3V{3�c@3��D3ף}3�e3L�3��^3�3
 3Q��2R�2x��2��&3äZ3��?3I�3��(3W;�3�m3S��2 ��2�3�3�f>3�&*3���2W�3~�R3Ght3�QF3$��2��Q3m��2���24iP3�S3�cG3�&3�.;3Z.3�9�23k��3M�
3�n3'493y��2�s3V�53/�3���2<3 '�3��3�3P�23�p3(F 3Ύ3�,3�V�2�\63�j>3�\33��"3(�3cRo3i�3�n/3� 3��2{?3k�.3�3��E3l��2Hqk3���3ߠ�3�FP3u	3�*n3R�43��3أH3^��2�3�@<3��3n�_3Z�2'�3���3t%3��2�w:3���2���2*=#3~m�3�C�2~^{36+�3�<s3d3�\�2���2��i3��2��3���2-�r3?�K3S��33 3'D3�L*3{4U�2�/3��2=�2�� 3t�3vU53���2��m3�3�)3SpV3��2��L3�`(3�=	3��23�Y�2Y��3+��2r�W3sp3E3��3��3��34C�3�(3��x3�G`3���3��?3r�D3JH3��3*�3�O03$a3~�3�d3�213j�83��Q32-3bD3v��3� �3��>3�g�3Y�3��-3��3b-G3/hW3�13���3�ҩ3�|�3NC�3�8�3��3�7D3���2�o�3QR|36h3�^c3�,63K�3a�y3U��3[�3���3��3�,4�lY3���3��A3]]3A+3��3�Z�3m3�Ƅ3��3��?333���2���3�~�3��2�hi3��P3���3r�>3��3�@3uM[3�<3(�"4f�3d�3.kz3�'s3�3�3W��3��!3���3jl�3��]3��-3h��2�ſ3�& 3"��2�3l23�fq3�Z�2n�3� 3� �3�][3\��3�9w3�H3p�3sË3p�@3��3��B38)�2y�`3x�3ګ�3��R3���2�b3+ve3Nv�3�G�3�֤2���3g�3`,�3��	3^�i35|W3tU+4LZ�3-�3��j3�X�2�h�2 х3
He3:��2lp3mʵ3�ɡ3��G3��'3�}r3�%03� 3F:3J�3���3�g%3�:�3�xC3(i3ʔ3���3/E	3�#'3j�e3Ƀ�3e�-3-5�3��<30�#3��3���3:�)3q3N�A3e��3��53PA3U��3P��2��3[�*3���3Ѱ
3zF�3S�l3�y
4�3+�C3tZ>3.�3��G3"dY3��b3B��2�E/3ó�3`�3�a�3i8�2OǞ3�'W3�3���3y5E3���36�3y�35�2�	3:e53aL�3ϡ,3�E3J�3PD3Ĵ3`)�34�3q�<3u3�M�3OԐ3��W3��2�q[3"M3KX3A�G3�fY3���3��)3뜴3s�m3b��2�C3к 4��>3@u�3���3��S3%�3��3i�l3�_3ɼ3� �3�i�3���3�	�2�P3<��3v|�2�8z3q�3\��3�ZE3q�93%��3�
�2Z�:3�[J3��2��.3)�3�P3�bt2t�830�3�2��2���3�?3Px31��2�
3�,�2��2��2���2��)3��25�53Ω3�x3L+3Gi�3�'A3��3�j3��U3��:3�|�2���2<��2��:3Yc3�o83��3�`�2�D3z~�3��?3���2��?2�]3�y3��}36+�2=�	3A�>3T�z3���2u3���2�k.3��2Y��2-3��2C�3T�3��2���2(��2��f3��3y��2��\3��2ɮ�2`�2S3�'�2*0�2>�3�XW37�3���2�7�2|J3�&3� 43��*3v0�2���2��3�q�3��Z3�+t2N�33s�3�]�2�O?3-�$3�K!3B��2��2�K�2��2U&�2xf�3l%�2�43J�	3�l�2�6�2��
3Z�2���2�?3fz}3"43D"�20	�2g��3���2 ��2B��2n��2\hL3��3֛)3��2�H3���2�%o3��t2mS�2[�n3$M3c�3�)3�*3˙2Au3�2�3ڊ23�.w3%�2��b3��2Ǽ�2{�!3\�2n=3�p�2�P3���2���2�b�27̘3���2a��2�� 3��2C(�2�� 3��3B7�2f63�.�3��a3�f�2#��28�$3ޭ3T��2�&a3���2e4�2���2M�3��21�2��2�ū3g�2�b3�3D`�2Q��2�L 3��3j	�2Q�!3�7(3��3}�3���2�7U3��2D�+3�T�2�2�3l�2I3�E3`J�2�g 3�u�3��2��2c��2�D�2�ɽ2;�2���2��2^�13T�f3�ph3UU�3���2�d&3.!R3��2��2� 3��*3Ci�2٣�3�>3�շ2Ԣ2.�~3�tq2� 3�2\0�2h��2%�2�3a��2TeL3Á�3Hf3��*3�đ2pd3u�2&�3jMM3Є-3׿�2���2 E�3ٹ�2���3¿�3p��3��03;£3�%�3���3KҐ3M �3@�31�r3s��3�� 4r�3���3	83�g43z�3�?�3���3R3O|�3Xi:3k��3�493p��3;��3�%&4y��3J 4P�3!��3�q3У�3���3p�p3�1z34��3�W�3��23��3�o�3��o3C;�3���3��3�`3��3�l�3\��3��Y3ob4��3�W�3��3/�z3g3��3,��3H�3K�u3ZU4���39xy3��=3o�3���3k�%3���3aj3vL�3@|3294/ˏ3�X~3%�U3*�4���3�g�3d1�3�a3�r!3���3���3��:3�X�3 ��3I��3��3O,3b��3U��3IhR3E�3�3���3���3��3��3uO`3�Io3�4>m�3�Ҙ3��R3��v3Cx3.�3�3��i39��3���3��4gW�3�;<3#��3�3�C�3`pp3��O3Ԇ�3���3Α�3�h�3B|H3뗘3h�3(��3��x3bG�3M�3�˅3���3u*�3�;�3w�3�M�3� �3+=I3m43"U420N3�9 4�f�3� �3�?�3�^k3Q��3�0l3�H13���3!c4���3���3��3%Ș3=͔3y3!��3��O3ה�3��"4�/�3���3��N3l��3	��3\�L3�k�3+�M3���3�[b3�ڻ3��I3�ʜ3�D�2��4��I3W_3zɌ3ݮr3V93ң�3j��3oq3�+�3�}�3OA�3!�3�]3���3�t�3�#,3��3��M3�U�32�b3k��3W�j38�Q3�Po34wLG3o;�34��3�\e3_��3&R�31�3vՈ3�E�3�c�3ڎ
4���3D��31�3`Ռ3� �30ʷ3#C3��F4I�3��3k�3S�3&Z3t��4�3�Ŀ3�E�3��3��c3v�3!�3aF3���3n�4��3�]�3?i/30B�3%N�3�]?3uŬ3Y3Rs�3U�W3�4ry�3uɎ3!�]3d�3��3���3D3���3�73*
�3�3��I3V+3���3&��3���3�D3�|�3�YH3�I:3�h3��x3,a�3�h	3�3�3�I!3�B	31.�3�13B�3
)�3&�3�3�T�3/?>3 �37�73cG3A��3z�]34��2Rz3Em3v�3!��3�/H3%{_3wQI36�P3(�Y3�-�3��3�43��2q�?3�e3�c�2�m�2k�2u�3�@73�IT3Ǻ3���3es	3���2
�63R�3�\3ث13�X63�i�3.�@3���3�%'3��?3���304'�2��2�Dv3�ں2�W3�23��3���2W$�35�3.��3�63��:3�Ȏ3,�^32��2�D�2��3pA3�-�2zP3u�M3g� 3��3PM�3�3��3��N3A3�e83�q 3�؆3ٿ3y�?3���3zJ�3�d731�3�{3�&3Q�3�cm3U23Q��3�(�2s��3=/3�IW3�iv3.B�3�h3ٖ3L�3��3o)?3��83��\3�V�2�%73=ͯ3E%�3EYH3=ƀ3Z�F3+{�2�K:3�>�3�2H�#3n�2c`b3�-3j�p3%�2�k�3v��29��3e:3�͋3{�%3��g3��3N�#3�q3���3oe3�`V3���2�^e3Ѥ	3��2�+�3��3\t3I�_3�U�3�{H3��"3��23C'4�0"3~9�3E>3G�[3�3JC37�x3:��2��$3�,�3���3I�3���2:3�2�3��%3V*3Hik2�:�3M��2�83`Q3p0J3G��2���33�f3qΏ3�ә3x1j3d�d3z#3zK33�V3'#13���3�y3
�3a�3�2w3#$�3�)3�X3�	�2a��3�c33?�3�x732׻2��2���3Y�3$K>3�>�3�^38�3Ѵ=3&CM3�F�2>��3��3�a�3Q��3���2��3n#�3�X3��Q3ҧ�2Hr3��83��3`-�3��3���3�?4(�@3s��3��3��k3��	3��>3+�3��{3��3ӌ3)��3.pE3�=V3zy�3�)�3��C3�)g3�F�33]3��3��3��{3}��3�x�3I�3̠{3
ާ3r$�3�,�3$��3p�j3{��3N�A3�hk3��L3&G�3j�`3Iyf3mQ�3(�3L&�3%Ȃ3�<�3;B�3 �33C�3b
�3v�L3�JP3 �3{��3�y3s3n�U3H^�3h��3���3�ǖ3?�n3 [04�
�3(g3�Ξ2u8�3�P}3��W3��3�d3�"�3ف+3h��3mn�3��z3�X63{sX4�|3YI3�=3*�3��n3�'3�)�3��"3"�3�s�3np�3�ۓ3&�-3�L�3"�3�V3PZV3ri3�j�3�N3_��3�[E3��a3ձ83q�R4�\�3g�D3�+�3|�53�H}3�;�3���3�K3Q�3��3�	�3߽�3��?3)�3�h]3��f3�J4h��3��3l��3�A�3��e37Z[3E�3�4w��33�3��h3�9�3�gD3��3)��3χ%3�$z3o 4�&�3_/�3yi�3,�3,�3��*3,z�3|�83��3t�321�3�Y3�ŭ3�3�U4�à3���3�Y\3��d36O3Ӡ�3i��3,�_3=��3�^�3��3�Q�30�D3�L�3��H34�H3gZ3f�73A�3z6�3�v�3�K3{�E3��_3Ya�37ʅ3��m3�R3R�3�5�3���3⣕3��37��3ˁ$4���3u-M3G�83�ك3ˏ�3��*3��3��
3|Ӎ3'�V3N�3��F3O23-9q3u%4�"03�~3ӓ[3��W3���2
�83=;�3t/3�λ3�_4���34�t3��>3�!3ide3�6G3�~�3903KMk3�Z�2v�3���3��~3q�3]�54j:�2H�3F]z3��3�i}3�N3��3$)3مZ3�84�4
�3wV�2�	�3=�3�I�3-�3��2C<�3o 3�x�3�{y3�O3
;?3��3FG3�@W3��32�'3���2��3�33�2g3��r31ٲ3���2(��2�*^3��2�3��!3��2��W3�:3dbe3�;	3��33��2塁3���2�s 363Uj
3�y�2�9
3��E3���2�3abz3yT3��2>�2q3�~A3�\3��03׾3�T3bj 3r3��3-�3�h3}��3 �2̒3t=i3ې%3~�$3���2�Y3~��2��	36�3��3P�3Ii�2��3c�-3�B�2m�3c	3�83x�3�Q3��2;��2ľ3I�3��2S|�2�VD3�RG3���2���2,K�2?�2NR3��3�<3i�2�״2���2��3���2	>23��2틊3@�3В-3�GJ3[�2h&�26f�3V�2��3"S�28�2���2��2A3�Y3;��27�b3��)3�I�2��2ț3��33,�3{�2��+3r��2��3%K�2�{�2��3b 3�13�2Y��2��3p.3�t3*'3��263�h@33~�3Le3��=3b�3���2�/!3���2v��2�f�2�]93Ir�2>=3L�3v�31p3`�
3�Q3f4�2<��2��2�M�23ۤ2g3F`.3OI=3Vm�2b�2��3��2�ܖ2��2�B�2w��2�y3a�.36��2Y*39��2�Y\3Eb�2ʵ93��2r�2[L�2D:.3wg?3�}3��(3�t3��G3�=&3:�2��13��2wv�2g�D3���2�'3L>	3
*3k3>$�2�b3�}`3R2�2ˍ3X063FV�2�q3�|�2G 3���2 �*3ҳ13}�{3���3B��2��3��3~��21E3�3�2�v3�538n�2�3{�2}�3Y��3�83^��2���2�!3As�2J��2�7�2�Ra23�3�|�3g43b�3��2��3+�}3�p�2���2A��2��I3�F�2.��2i�2Q�3�y�3�F�3��B3Gi3��Y3�~s3(�3␘3Fan3��/3��3��3zj�3��3�3�X�3{�c3�H3YkN3{Y3���3�	3�ե3�J�3b^�3�i�3�ֹ3X\3=Ff3��V3r��3��63rie3���3�Ϣ3�5`3w��3���3JR�3j�.3��3��E3t`3� 3�]^3�6�3��B3���3�m|3��3��3���3�8�3�uo3�M�3ށ�3�J3!�>3�L�3'��3Ҝ�3��4E֘3:PJ3�OX3:�z3� �39�D3���3O�|3N��3�So3bů393��3�93��4n�33�a3�q�3���3�Hu3���3Li�3��=34׆3�B�3���3�3�N3@�13��43XU3�:�3�7.3�+�3��g3e��3��^3�P�3��3��4W�3?+3��d3�1�3���31�3f{�3�#(3w�3k�3zd�3�ח3^~.3,o�3��3�
x3�P�3�d3�2�3C43���3�ā3ҡl3�43��3p�Q3�hV3U�f3�L3 ��3�63.��3_�3�D�3cl�3��3|�F3��[3�ڜ3=.�3�R3��:3ll.3�3C�3h�3�k�3n/!3�533�4�3��3m��3ӁB3-fq3�q3>�g3�T3�\3Rh4C�3���3CO3�C4(.g3�q3|�3X�'3���3�=3�F�3A��3e�F3���3�)4LW3e�y3i73�W�3Yvs3h.�34*e3�5,32J�3��3>��3V��3V��2�\z3Las3�`37��3��x3�/^3Voo3���3�&3`�Y3h�V3Ë4���3*�3i��3@ �3�M3�Q�3�ŗ3��J3%}3���32��3�F�3�l3�U35�H3�j�3�"�3#?3���3�^33�m�3�ɀ3o�<3g��2��3�p�3*�3�$�3PV�3�^3��;3�#�37� 3�I3Bv�3���3�D�3-�3�R�3�'�3�5W3�z�3��3;>�3�8�3��3<}�3��4�8�3U�f4���3(p�39%Z3�Ԁ3��\3�a�3�,�3��3�a�3���3144��3�(4O��3��F3z�3���3<�3V��3�}�3�K�3
�3J73D�@4�_�3ɠ]3O��3���3xê3�Ư3���3m3���3��;4f��3��3�ɀ3�4P�f3�J�3SW�3�X�3푖3O��3Ʒ�3���3�=�3���3��W4@�3�/�3��32��3^3�/93$N4��3���3@X~4(4!��3&F3���3��;4sB3	I�3��j3�T�3/7p31�
4*	�3	��3;پ3_�`4PK|3v��3U�3V4/3�3{�3R�4�:�3��3���3s��3ǃ�3�[3��4� 4�G}3w�3D�3�O�3xL�3�D�3B#�3��3Q�3��S4D�3Xs�35�3{��33��3���3�?�3��3K��3GR4�T4��3��2���3&^4z��3}��3�>�3��4n0�3*N�35��3���3;R�3��v4߆4P\�3Ʈ=3Zu�3���3��3
��3'��3�4�3:�$4��+4؟�3���3���3H�F4V��3u��3%��3q�4a�3H��3F;�3*
4k�3�!4�s�3Xe
4��3��3��3�W
4���3}ǲ3n�3T44K��3/r74���3eq4.u�3��3���3��3�s�3+��3ro'4 JV3�4�6�3�Y4 ��3��3�5�3��3���3T4�Q4Ŋ�3ѱH4^l4/4�=4�z3��3��4�β3�84~�3�v�3�4n3d�,4��34�34�v3U�=4�)�3nZ~3���3ԕ�3��3Fv�3�\�3#J�3�4 �	4��3��3ۺt3�32,4Yn�3�Y�3�y�3<�3r��3c� 4�[�3?ԁ3�j�3��4���3���3�;4K2�3�Z�3�[�3�J�3+i�3>�`4�+E4.H/4�->4��m3X��3�4�w�37�$3�n�3��24ڙ�32�^4n�4���2W��2\�3B�g2�c2e�2��2�,�2�{�21��2Ck�2�_�2g=3��2�=�2f
�2h{�28�2��\2�2�2L �2m��2Lrw2b�3P�2=&�2�B�2/R`3|�2�T�2'��2��2vR�2�R�2��3��2?�2ٵ3v� 3��3AD2��2i�2�OG2KN�2�ݵ2���2��2��3�m3���2̫�2n+3q�2��2�B�2�o�2�24ߥ2�q�2�v�2��2Ġ�29��2���2�_`2V[�2��2��72��2��2/W�2�QH2�2'E�2I�2��2�A83Ŭ|2ȵ�2{�2a��2Ůq2H��2��2��A2���2��	3��3ٔ�2�'2��2��2v�o21��2��2�2��2��-3���2}�2��2��3xy22�o2~ɜ2���2Zi
3���2�i�2��d2h?3��3��2F�27Bh2��3
 3�2���2�	�2��2ea�2%�73�i�2���2	�2�3�s�2	d�2$�2w�2���20��2f��2/�a2�^�2y�3�3@�2r�2$��2KS�21��2�V3W�2�W�2��2�)�2�H�2x�2"�&2\�`3?�2��2�#�2Ζ�2s
�2qc�2�Ez2㙧2���2W�b3x��28��2�2|2t�3j�2b}s2q��2�k�2U��2Qt2�33F��2�k�2?��2�V3
f�2��2���2���2�d�2�J�2�3�(y2�	z2�[83*V�2�%�2`�[2d�3���2*��2��2YrI295�2N/3��3	��2گ�2���2P�K3d:�2_3�I3հ�2�2���2���2�c�2.��2*K3Q��2���2��23�M�27��2=��2�kB2�23�i�2��#3+T�2h�K2�]62��P3��T2�Z2wp�2��2?�2"7�2v2��L20*�2V� 3}��2�2H�~2�@�2�R�2L�M2���2iw%2
73�n2�\�21A^2���3��B3�% 4�e�38��3��3NJ,3e;3f�^3�KX3���3�{3�4���3$n�3�=3�m�3d`u3�qa3+"[3#�J3�C3�O:3���3�0�3���3Z�3��3�G3�y33�o3Z�3k��3E�B3E�q3>s3u5)3FΣ3ҵ�3+[�3۷V3��33K3+�W3�{k3D�.3k��3қ�2��3B-35�3"3,��3d�T3e}�3��&3'��3�X�2ki3��3�u�3��A3�UL3}r�3��3 �3�\�3ե�3M3(��3�4"3���3H�a3�Y3z%J3�\�3�_�3�%4�!$3���2�2b3!x�3�c 3��3m;�3��2��t3D@4��3�aM3J�3w,z3���3F�#3�:[3G�>3,��3=�3ʨ�3~d36xB3�;�2���3�wZ3�a3��34�M3_�k3{|]3ע3��2�Ox3��3�δ3�'*3QB�2i&�3��3�3o�V33�T3���3Φ3>�>3Qu35�3��3
2.4 U 3V��3��3��a3��#3�;3=~�3��$3�F�3Uڙ3W��3T�33�\3�۠3�U�3�v3A�/3+�3?=�2��3/ք3��K3�ۗ25�4.N73OL�3D'3w_3ͱu3>I\3{܀3��*3���3�4�Q�3�@3'�"3Z_l3��%3"�$3[�3�	3 �`3lt3�Q�3Y3Ð�3�m3{b4g>o3�!�3�3�P3�+3���3e��3�2=2?3Ed�3��3��R3r�2�%�3�N�3�43�U�3��3�^3
3�+�3�v,3�v3^�3���3<<3S�\3F�3�di3��@3*V�3X	Z3S�3�U3��;4�P�3��A3]3��a3��73�S3^PH3�,31��3��3.�3ɐ�2��*3���3ż4�^o3R]33f}3�&3�D_3�Ȃ3��=3��2��3, �3jބ3�&W3��T3��33^U3553o΢3�T3O�h3� 53�B3�J"3RL�3RT_3^�4=h3��v3n�3ZA�3���3�l�3(�83��3��3c��3O�3�`4��3O��3��3WoY3���3Da32'�3�C{3��4w�3��3"�3�ՠ4"�3��3)�37��3}E3��4�3�<�32��3�r�3�#4�94��3��D4۝�33Z�3���3%ʻ3��4��3o|�4E4�3ah�3_��3�ku4���3�Ω3b�3�X�3�m�3�{�3�4(�3�(�346�<4�F�3���3���3ϖ�3�v�3.�C4Y3g�!4.��3&*4f��3�Q�3��3���4:��3 ��3�Z�3��3��3���3�u,4��=3���3��4��4��3IȬ3�Ͱ3�F�3��3�]�3RT�3�,&4�$\3�4c�P3��x3�x�38(4���3�!4��4���3@��3�� 4y�C4�g�3��3��Y4���3���3���3�{'4��48i3��34�i3qA4�$p3W9�3���3��3�jU3՟4�B�3f��3l֞3�Ъ3p=Y3���3���3�\�3��3s4�K04�@4�Fv3���3�4Tf�3D��3$��3Xy
4)_�3��3#��3'�3��3�o4��3E�3鄞3�x�3�!4#�-4� 4�M�3h��3�'=4'4�M4��^3��#4��3Hx�3�+�3��3B��32��3�$4�g�3 ��3'�3�%�4��3�<4�P�3�K�3d߾3Ć�3�4[z�3jh!4��4@%4��3�@3��3���3���3�-4��3�o�3]sg3�#V4��4���3� �3��_4v�44�3�]4��4m��3�,�37�4�`3α4$��4�;4���43�~3���3�KZ4E�37.4��4�(4��3,�4Ά�3<
�3�3�˅4�3 4��3�Q�3��3'4iŘ3o>3V�4`��3ߜ>4C�H4!Þ3W�3#�4�(w3E�4�_�3M�L4��o3��C4� �3��J2T�&2Rw�25��2K��2��O2!�O2 =2�2VX�2۳2�Q�2i��2�>D2�̒2咋2�-�2�2��G2�1�2W��2�Ϡ2)\2��2.x�2���2O��2��2��L2��2�2�u3�+2'�2(��2�Ȁ2A�[2��3t��2{A�2��1ۂ2!��2�:2�`�2��2�@�2~+G2yw�2�ȵ2��2*2�U�2ǎ�2��2r�28[\2djj2C�)26�2�DX2w��2�M�2�U�2̵2�� 2:��2+��26�62��$2�Pz2��2�Z2̹2�|2�t3Y�2F83}�2�e�2HHw2��l2���2|:�2F�2o%121D�2��3|��2$*2$Z2�>�2��=2�42���2~�:2_Lg2�t`2���2�z�2�J2�G 2Q��2{l�26^2�n�2"�r2!�J2�2*Dx2��,2�]�2�W3�TR2�72�@2�ݷ2�ϣ2hC20»2���2�O@2�-2��3��z2�([2 ��2��<3%�O2O��2�g2�!}2��25�E2�q�2�Y2��2�)39F�2��2���2�2���2:/{2��,2*S2���2]+�2ye�2l��2��g2�[2��2^��2m�B2���2�b�28�32"�2��2��2q�2��3��2"/�2���2֎�2���2>H�2���2C4>2׮|2�%42W{3�~Y2�[`2d�]2�8F3���27��2E��2��,2��22��2���2�i�2s�2�.�2r��2�#�2��W2D�2��e2e�#2�Ď2��Q2�f�2N�a2J.�2�ɘ2m��2J�2i�-3�mD2��2�
"2O282Nʇ2�]w2|�i2Ɣ2Ӹ�2��3�1m25�R2|}�2�_j2�lN2��2�C*2�m�2~��2���2�e�2�e2 �2>�3�2b�02G�212�CG2
832
��2;�72�Ut2]k�2됟2޶2{D
2 �2Ħq2p|E2z��2W��1Ϝz2V22l�2GO�2��3��2L�3kr�2�S�2��&3#"3�C�2_Q3A 3�P3�#23\T�3O|�3�23��2�б3�Y3 ��2]�3��2F,3�2N�3 TD3�A3SP@3�ܥ3��V3t�e3�b33�S03�k%32o3��3i"3w[c3|r�3��3��C3 '3�ֵ3��3<��2�AB3�H3�^e3�M3�k�3,	h3Q��3��3�ߕ3�I3��;3\kM3�/O3GZ3c3��,3���2
�*35��3�wn3C�j3�t3a/23�Q�3@!33�3"A3��3��
3r�r34kD3>/3x
3��3j�3/T_3�I�3�IL3�*C3�.X3�.N3D<#31^3���3GRG3��i3��2��3���3�3E�3˪�24�3�h�2w�3b��2��3��f3#}�3� ]3Ȅ�3�	�3ݫ�3 �3ŰR3��3OY�2x5K3?lm3S��3�}73a-�2��R3���3���2��p3�#�2��@3"�3�ʓ3%w737�>3��=3{�37�2��3��3G:�3�B'3w�3�_�3���2iC3�[�3MN�3�3�H3�uD3R/3r339�3Ig3d�3�O�2�M-3j3���3_�U3,��3W��30!33��3�m=3v%k3eVZ3t3?M�2ٵ&3�c�3PC�3��23��3B!3��Q3s,3��3�,�2's3C�^3.f3�_3��43׮n3a��3�o3��g3ȑ�3Ç3	3�y3�`83^�3ӵN3a��3��3m�W3�A3.o�3��3�A3��\36�3�.3|�3 ��3��3]!)3��2��4��=3��@3�N%3�|3��:30^^3�|33�A3G�k3��3r3��73U��2;�O3��b3E�2�J�348$3n�3*&O3�b�3��3</�2��3[�3�3.3��33��26aI3��<3TZE3��#3o�3:��3$�{3j��3�t�2/:3�=3�;�2�3�7�2-��3J�J3��P3��U3��3Z�2�:4ʶP3�ۍ3��3.�4>(13,�V3��F3�U3���3G6�3(o�3gC�3��i3|�v3hyV3�P3��C3y�3�i3X��2=4��3� �3�<�3�Q
4�F3���3q�3�G�3�|3v��3�H�3��y31�~3.��3^=3LGa3��3VW�3_�p3���3Ϊ�3�h�3�Wh3h�Z3��3yͥ3L�43�B3��4��<3'o3��3]ա3��43��=3��3V�3L�w3�	4 *�3 Z3`3�Z�3
cK3��2Ur3Sp31kM3��_3�N�3��53�b?34�3x�3�);3S"3�3���3�%<3P�33&�3�5.3yb�3�3Xz�3e�f3�A3�S3�x3���3ש�3E93�-%4�E3$pw3p�(3��_3��p3{34< 3���3S1^3`�3�X33�B3l��3~3�;b3��3���3^Cb3�3�m�3��3�p_3�
�3w63�7�3^8�2ڔ�3�3�36H3�5�2��3���3��T3=�3(�3a�>3���3�v3���2�D3<��3O��3�B13��43)ֱ3���3��3�3b�@3W�4@_`3�?�3j��3U�.3?�:3x�4��j3g��3ϋ3�3�{�3R�3K(�3��3���3��3q�3��3�G&3T�3A3['�3ɹ�3 0!3�у3�q3��3{�p3���3�w3>�
4_��3a8�3���3���3wp931��3��3���3tՊ35��3r��3��3�gZ3v��3j�3�Ɂ3�i�3�l�3�-�3� �3�}�3;ݩ3�vt3	ob3�ߠ3hz3=m<3Gܚ3#13�d�3�p3i�{3>F3��3�W�3(?�3�ʩ3	3G��3���3��3�Zb3��y3�31:3-[�3�H�3�,
3�Z,3й�3�z�3l��3|�3�*t3�%3�@�3$�30h3��3H24���3��3X=3�3�xE3�3���3�S3:��3�L3�Z�3�
A3)�}3ҿ@3���3�53� �3�`13�B�3In�2ͪ3�d�3L2�34�!33i�3��3�+�3xL3hW�3]�s3�2��O3��3X�3h�/3V\35�l3_D3el33���3�7�3ɯ�3:|�3���3YX`3X923�L3�0b3;h�3[�3�r�3��a3`Y/3h�3�QT3�@h3ߙ�3`33Hx{3T��2mG4��393ƜQ3>�*4�5^3ܑ23���3DD�3��#3@�03AE�3�,3�ge3q	�3�ճ37!3�2��c3Vd�3�3Ոj3��@3��h3�>�2�hl3bE3gO3jSI3s4��3�q�3��%3.3�hL3�3��T3��d3�J23R@�3a��3�MK3��@3���3w#�3S��2<ɓ3.�n3zH�3�Z*3��o3�.(37�3Y�3�v4ҁ38%v3>�%3�I�3��?3�O`3EX�3��43'��3�I�3HA�31�2�_3Q�3S�3Z �3��G3 �3v��3B�:3��3P�3�p3���3��s3723>T�3�Wa3G�3 *3�Y�3�p�3��L3�z3�q�3CX�31�3�Py3�-�3��3�3|<�3K|U3��3���2�wu3���3W�T3��3��3�\3�3��3�3�F3�13~�|3\�3g3�3��3I��3��3�3Gb�3���2��3N��3�2O3'FB3g�4�v3��:3G6�3Ug4Yx3��}3�ML3^�33�3��`3�ȱ3%A,3��3�I�3#�3bEo3W&�29%x3��3Va3�P3k�3�!�3��f3���3��A3d^3��R3S�3�N3C�3Au�3^&3Y,3%�U3�3�3)'3�D�3}B�3N��3��3!S�2��u3�Ӈ3�JS3(063�7+3�=�3�mF3I��3�M3p�53w3B4�+3v�I3|x3�P3x[>3���3�F�3��2K�3:f�3G$�3Қ�3��2(0�3�Dx3Ϻ3n%�3�	34b�3ڍ&39��3�si3#`�3u��3�T�3?l�3�ǲ3�Us3��4*~Q3�M�3���3	�3�{�3}�4��3&�3�"3q��3���3��"3�r3��3��3�~-3�3)��3���3���3͗!4���3�=�3��33E�3��32S�3�3k~3�l�3�!4���3+�3r(M3�B4��3���3)��3�2�3_O�3<S73�E 4橙3@��3نq3�(k4���3��3s��3c��3��]3\��3�t�36�o3�$z3��3M�)4�]�3��?3�D�3�"�3�]53�l�3̳_3}��3of�3�:�3-]3��k3d��3�M)4�!�3LX�3z}�3�74�at3���3��3e�&3�D�3
�4+��3���3�KU3��3���3B�3Ry�3�P3=)�3Xa�3M�3n��3�܂3c?3S�4췙3�	�3�3���3t�z3���3��3�!3��3 �4� 4�3͓Y3�f�3R�3� b3L`�3W�3���3�5H3���3�?3:�T3tH�3�>4�3+8�3�m�3��Q3(�3��3�,�3�ʖ3�Z�3��4r�,4U�u3ؾ�3�s�3�/�3�m37p�3��p3P?�3>˾39Z4��3l��3�@3j34��D32��3O��3�u3">�3��3��}30#�3	˃3���3q�4�W�3(x�3��35�3��3u��3aŅ3���3�Ư36 �3n K3��l3c3F34��3��3�Yd3�KX3���3��l3-�3<�3�e4�=4�' 4��3��n3@s3���3Wj3�y�3��e36<�3� 3�4I�3D�3�wM3�mK4�v3�К3���3�r�3��[3Ɍ�3٭�3�}+3�۷3�%4��3Aת3f3*�i3���3�<�3�޲37L3���3~
13���3��3"03�:*3r"4��3���3��a3�؎3k�39��3m��3��3�w�3,a�3�A4uX�3h�+3��3�'�3���3�G�3�B3��3հ�3�3���3��3DJ�2a�E3a�3<��2Ke&3 �3Z
�2���2��	34z�2�Z�2��.3(�3��3h��2R�Q3��3@=�2���2�3��13�{�2�<3��3���2�e�2jxN3��2Y3}{.3x$�2��|2���2G3��3C�+33�.3>�39,�2��03��2��3�O$3E�3�H3~�2��23��3�73�k�2E�c3�e3D�63*��2�e�3�#3��36�2/�}2���2-O3�f3	�2DK�2�F3�B3à�2 �3z�03dk 35�2��
3S�2!�2��	3q��3~	�2w�2j!3��2���2W�2BQY3�8[2}�3�"V3� 3�3a��2���2=1�2�+�22>3"��2��2�F�2g�&3���2x��2�Ƭ2��3�3"��2��2K��2��2�^�2���2X�2"z�2ƲI3,�2�|�2IR�2��24\�2��2Rm3rF�2Sm3�l�2�
3�@�2�Q�2���2'�3���2iJ53b}�2�(�2��2}��2s�C3 �2���2k~�3'G23Y��2Y��2+=>3���2��2���2fo�2�H
33�:3��3��3��2���2E��3��2,`
38o�2�-3e��2-�@3��53�12v��2��g31�M3|�3���2�CS3�'3��2j�3���2]�3��3�q^3֖	3�Խ2tb�2>֦33�2o��2��93�L3"��2���2��!3$�c2Қ�2/�N3��'3��M3���2�3��2$��2a3��2��<3���2ϨK3��3���2���2���3��2���2T�3Y�2��2*t�2gY�2�;�2D^�2�&3\�3*/3a43�7�2Ѽ43� +3�R�2��2z.$3(�2�*3��)3Y;z2+82��l3��2H"m2�g�20�3�R�2��2�W3��2�~�2�y'3��:3��2�J2���2���2z��2�$3��2�@�2�ټ2a�J3m>�2r�38Y3�*	4y�V31k�3��`3�d}3c��2rk3�Zs3w|!39\o3��3|�u3���3��W3
q�3-��3b9+3в3VN�3�<�3�f3!��3 �z3+��3��[3�Z�3E+73��D3��3⍖3΄B3��3��u3��
3G8Y3��3�_3��f3���2}3˂U3%�q3���3�#831��3t�X3s��3�5V3�r3�
�2*�3	3n.�3��2�$3�� 36l�3]�3�G3�yt3l��3M[�3'�`3 v�2Ch�3*kF3M� 3�[n3�a3�y�3m0�2�3�[3Ű{3593]��3�C3��:3|��2|�[3�:3_1O3�֎3y9M3��X3��3�b3��m3�U�2@}b3;R3jm�2a�j3}Y3���3{3~M3;Ƒ3�63��c3�H�3-i�2h�73}�3}L3M�>3wb�3�Q�3w�3���3�d�3&k�3JZ>3@1�2��3�	{3Y��2@q�3zv3a�h3U[l3��3;��3�C!3�~'3j4(�3��3�j�3?>�3�>3�3��3P% 3?+_3$�3�9�3/��3��2tGM3�l�3��03_ك3$�3ci�3U�$3xj�3��]3|�3H13�k24��`3s(�3��3p[�3�Uj3�JO3�^3T�3��b3<�3�hr3wk3Y(3��N35�+3]�3�l3?>3�Xq3��z3QX~3�@3�x�3��I3z��3g9P3�ד3��n3/�U3*c�2jN�3(��3+�3�vt3���3���3xʿ3��3���3��:3�g;3�V�3D�A3�+3�H3�j4U<3_G3v'V3m��3+}35"T3�Yz3}�Y3��3�33�KP3��,3��P3֘3�E�3G-u3YX3G��2�j�3\3��3�4:3^e�3�p�2��(3�I3Nf3�W�2��4g#53�Th3��3q3�%3�U3K�3�7�2���3?�3���3�M53z,�2"�f3�=�3ac!3���3�"3���3�F3}ȯ3z��3u,23A��2X�3Y�73��R3UU3��>3F;3�f3B�)3�R�2�\43BI�3��93�,c3�T�2Ʀl3��"3]-3"��2X3��*3;�2?��3�D�2��x3�l�2�l3|�B3�73&�3�kq3�.3@F3�]3��*3#o&3��Z3��_3l��3���2�p^3�3�}3��13���2O3F�
3�Z3H$3�cA3̿ 3�R�3)P-3�D3�*3�+C3�
3��s3)�&3��3 �3�΄3?e�3��(3J��2Psi3�'30[Q3��-3�m)3)�3��2�ib3��3�y73��%37��3{�63��S3��p3�V"3�A�2!3�2`H3��Q3��X3��3�w�3�-3��3G��3h4n3f��2QE3�?3�E3%�3Kp^3��'3|+T3��3��3� 3��3ݫ 3�p3��2�73�303���2�3�K3�	E3S�C3�I�2N�3	�2SK�2g=3��l3�935)3��w3�A	3ݰ�2��3,d3_�"3�b,3��R3��3[�3Z��3�03EV�2r�!3�{�3�3��2�43��3��<3b�\3~23�=�2�g3T3�c3��63�*#3���2�3�ق3�3�3qQ3��2�>3��3)�3n&�3*��3Z�#3�v3���2���3J:3��2�>l3"~�2�d3�r3
q�3�-�2�4 3�3"�:3�� 3�zD3t/3�/3b�E3_�-3��]3^��21B3��X3���3+W^3]?3��3�MY3��83y,3'�X3N�|3��;3\v}3�K3�T,3�'
3���3;�L3�!;3��Q3�=3�T3zpP3R13ʇ3��3� 4mL=3��3��v2\�83^6�3�	3��,3�r03��}3A��2���3n�3D��2��d2��3�%$3�M3r43��{35Q�2���3HeO3��23p�3�n'3x�r3B�2(�X3�
?3�m3�z*3~�2��U3�v3D�03�3_��3�E�3L�4"x�3�D�3��Y3ȿ�3�G3M�}3j��3��B3��:3
��3�L$3���3,�3��3�z�3N�_3z�U3ٌ�3�3Q+l3IO�3ﮒ3��T3��>3ϧ�3k8a3��|3L�~3�3�(b3U�3��3X��3��)3O��3��E31�`3� 93���3ǃ�3ƕL3�k�3��Q3�i30��3��4�G3�v$3ݦ\3�24Z��3f�X3E3�zr3�W3ި3c�3�Vw3��v3���3g��33	U�3WK�3b�n3���3Y��3�2d3>Ƴ3�)�3�	�3ON�3n��3�Q3#A.4��f3d�j3yE�3zY3�"B3�}�3c�3��2�[�3���3�j�3�>3��3zQ�3.z3�rB3�3m�3�ݾ3�q[3L:4��73�L3�&3�4m�3�њ3&��3f��3�	3�{�36o3�4d3!-#3к�3}��3k�n3G�3��3�M�3��M3�Y�32�W3�ƈ3��3/z�3�ф3;�q3冩3&�4�?33�|3+�3T[�3[�e3���3wW�3��3�}�3���3���3�P�30Cw3�N�3�1�3bA?3x��3m��3ƺ�3u�3�v�3p�3��i3��3*�%4�.Z3H��3�53m�]3k�R3?�4'߬3�`�3�S�3���3��3O��3߅�3���3�݂3��A3�2�3: �3�3��3��3ٴ�3/M�3��s3�!$4�c�3!�*3a�3�3m�w3��3��3��35��3Z��3��3z'z3)�#38X�3�O�3CS33��3�1�3� 4�/�3���3]�p3D �3벽394���3خ3�1W3�i3f:�3���3���3�:3��i3��3�i�3V|3��v3�`W3���3�g�3rF�3�aY3�߻3E��3�(�3�^3��=3��Z3V��3���3�#=3y�3���3��]3�mh3�͢3T3/3�(�3�4-�3>��3ZC3�.�3���3]�e3�7�3j@d3j��3�D�3P�4}Ӭ3'��3�E"3�d#4�؅3hq�3TW3�04:d 3��3g�3'q�3��3�Ҋ3�X�3��3�Y3r�3��W3�3��33ޥ3�Ic3J#�3~)�3��3��36a�3̦3�P�3��3���3�σ3��3'��3�Ɵ3�k�3a4%��3�14�v�3o�3g�(3$@"37�=3%�3p<Z3D6�3�!�3�[�32��3ȩ<37�4<p3�C�3h3/iH3���3���3h3o�3���3�_�3E��3���3�L�2��3��3�Y3r&�3��H30��3|b�3K��3��&3��3��3P�%4��,3��3k9�3A�I34�13�Ն3&��3��i3��d3��3��3h�3T$32]�3���3<�3/a3�1�3	.�3`�I34�3�j`3���3jZZ3)�&4�.3��33�^3b�U3Pa3}��3x��3�#3��}3�2�3k40N3XXK3ι�3�G�3t�3D�3#�93���3i�3��3�=3fq�3���3m�4Dɀ3w��3/b�3T=�3Q|�3�\@3cx�3]33 �3�L�3Kc48F3�v3r�3R�3g[3G��3��C3ȼ3d9�2��3�EG3��N3L35�4��3k��3���3?�Q3�:S3 �3N��3��f3�$�3/L�3S��3?,�3�m3rl�3��F3{H3"�4��<3�X�3�_3b
4!@3���3Hd�3�F�3��3@��3y�3q3I3���3��3�k�3�U�23L3��3��4>j�3�3���3�Ĕ3ݣ�2��3��O33�S3�o3��	4��?30�=38 3��3�\?3­�3�)4�3c3#�F3Q}�3��L3���3�X�3�A�3>�3ǟ�3*J3W�3� �3'�3���3�s�23�L�3m�d3z�38oL3K913��3��i3Oܡ3֝3v
�3�^3�jR3˅�35F3��3���3�3�+�3d�)3��3c�L3�RD3p��3
m3Z+3�13���3���3�u3�ǁ3b_�3w�3�V�3Ñ�3!�N3@Ʉ3���3)��3�*[3ᇄ3m��3H��3���3�[3���3��B3�,�3Ͷ�3~�t3��3<k3c��3���38�3��3Y341�[3I3�H�3�X�3R'`3|�v31��3�+30�3C۴3q4#9�3fE�2���3[}3އ&3�'?3�"`3�N�3�RZ3w �3�4�3��3,3a��3� 63Y>:3�J3�~�3p!=3��3�ǟ3"3_�3r�3B�3���3�c 3��4�R�3��3Ğm3Dk3��3ݏ3T�33�*3�x.3W 4��4\��3ci{3��[3sx534ѐ3E^�3��	3}�2�j�3i64�-�3�N3�[3��J3n�f3��E3�#�3�1�3C��3y��34��3�2K3�o3]��3���3�w.3��F3�u&3)3H�3�n�3 �3O�53mx�3���3�y�3'uH3��;39e}3)�3�
3�v�3��3|��3<ݬ3}��3G��3z�U3qȪ3��4��2m�q3�ۯ3㋓3 ��3��3�Ҩ3;3��_3(:�3��y3u�m3��R3��`3�5�3Rv.3M�N3�"B3���3A�X3�k�3ڳz3<tP3Ad�2�4��r3��P3`�[3�S3�93�`K3��3�U3>�3���3ֺ�3Z$3��2��h30�;3�#3��\3ދ�2�@n3��3�oy3��C32��37g�3Q�4�L3[f3��E3�CC3��"3X�3H��3<3R"�3CO�3�Q�3�}3R�V3��3�3`3;3@��3Y73���3�==3ɨ�3B%:3�|�2Mb3��3��=3�t�3N�3h��3͙S3�V3Hs�3�f3A��3*�3a��3���3��2�O�3��3s��3�D]3��3l�37|3¾�3�|�3��I3cL!3)�3B�T3���3D�X3L�3��3IL3\�34�3d߮3};�3�w�3��y3Y3,��3��33_F3i�*3>��2NJ�3
�3�Mp3I�33&�3��3���3��3l�E33��2���3~3ᑑ3��3:�[3��3pT�3�͐3��o3H�f3<1�3�DZ3�2��83�gL3��3�R�2�3�3�j}3���3�J/3��4C,3��c3�s3?L�3�{H3���3�X 3%I=3�%*3}�3i��3�K�3���2Ř�3�`R3��O3�w�3�CS3MbH3�(#3��3H:3X?'3��z3C�4��(3$�3<v3!!3D�,32R63��Q3�_�2�JR3��3/[d3@�a3vP�2�;f3�M�3��3m�363t/73`�3�W�3�r3�)�3��53�3��u3�z_3�3?�k3vR.3�{b3��3�� 3e�|3��$4���3w�U3��H3F��3s��3��J3�}|3��d3�%�3$39ܞ3/@3K,3'�W3��-4��Y3�υ3U�3:}p3��'3		R3ο:3�3J�s3+�3�T�3ǟ�3��3��u3��3�
36n=34b3�ڍ3��F3�L�3�h53Z�Q37�039(�3��323��T3�j3�F�2���3�#q3�u3��3g�3�%3��g3��-3a �3�3�Q�2b��3:;3�}�3t.,3�*�3��X3#@ 3�]3�C4u�3e�3o�'3�E�3��^3���3���3��?3Sَ3���3ti�3
�R3SsI3V��3j�_3�A�3-�3 �3��3uqK3�_�3��3m)j3�13��3�b3Ӌ�3�T�3�
�3�83{[%3�3�m%3��3q�3_�3zɒ3\�'3 ��3,�83���2�[�3j`53P,�3Z�3=��3�R�3xY�3�3;+4���3�H:3"�3[�3�� 3�*3���3'��2���3��V3���3�R�3���2�|�3�4��3��3��E3�F|3khf3�̮3�؅3|53T3�q�3o�K3�Y3O�03��S3�z3�t�3[��3L�3�4d3�/�3S�3`�g3�r3�?^3�3BQd3a�3�3�2�}�3t$3��{3K�c3���3��3��34a~�3���3�v�3=r3��E3���3��3譲3�v�35Z4u��3J��3��3=��3��m3|}3��-3��3��4���3���3���3O�3+�3�w4�-�3B�4���3�F�3���34��3���3�p�35d�3e�3�κ3�Ώ3sџ3=Ҩ3!qx3�{3q��3�}y3+��3ώ�3G��3g&r3��}3��3BB+4)��3�M�3���3�(�3�+]3�i�3� �3���3k��3�y�3=��3�f�3�kx3%��3Z��3Pqo3+�4@�v3�|�3`5e3���3z�3�F�3��3o84�E3B��3,�3yG�3���3o�3_ 4�0 3 ) 4�#4pk�3���3�0=3Dc�3���3�}3�Ϣ3"@O344+�3ݱ4�Ys3�S�3^�F3�X48<x3�~�3���3�P73���3��3-V�3m�c39�3�+�3R�3[M�3��n3X��3���3�7�3��4��3�ܳ3�S3B�4��#3ʿ�3��3t�
4��3�e�3��[3�D�3�@�3v�)4y^44��h3�o�3@"4���3��b3�	Z3�46��3r��3Ԫ�33�23�5�3��3�B 4@�4z��3���3`�4]�(3��3kZs3�#A3���3_(�3��3�d�3�S�3O?4��4;W3A}�3��3
ȥ30�T3e��3}=e3�Γ3Q~�3�L�3��`3�Y�3aBf3�T4rrb3 �B3q�3�\�3���3�A�3�3�3�;�3�U�3�4x��3��O3y�#3ҙ4g2�3{�r3$��3�R�3���3|SB3�14\��3�	�3x��3WjX4��Y31�36C�3p�*3`�3>%B3@��3{�53���3�k4��4؟�3�!�36�3ui>4���3D4�30��3<S35��3�l4�p3�R�3�)�4u�4G�3=~�3a�3��23!Fx3��3��73G�3�B`4�4�3?�3��
3,ܔ3���3�N�3o�/3)ID3/.-4��T3Z�3���3���3oxu3�� 4s�H3��j3�L3^k�3�1�3��3y�A3?��3k��3�Y 4�u�3�b�3~�$34G4k�3�)3��3軄3�k�3O�/3��4�33b��3�?�3��4J��30�3m j3ご3sEm3ƙ3�>�3��3tՓ3�4�3wb�3ᇍ3}b3`3(��3
�R3*�3Wc3���3���3��3�)p3ɚ�3��S3B�C4H�3���3A&�3�Rj3�n�3�3�3��3�S23a��3�J4-��3�9�3i�<3b��3-h�3�E3ИV3�83�X�3��3�Ѓ3�2�3���3j�=3G64�;_3��i3_F�3#t3ߒ3ڶ�3\_�3��3֨�3#�-4��3�2^3|�)3SN�39�f3�Z;3�U�3��3n��3�X3K��3�6?3n�O3��3���3�o�33\�3E�3�k�3%�33ݞ3H��3��d31�3:/4�� 4���3H�83^�)4�)�3]��3�84&�?3[�3�և3Hn3��k3��73�8Y3��4ڪ�3�|3�>3�~h3�L�3��r3��3�ON3��x3�W�3�}�3���3�q3H��3p��3�3L�3\�63y�3��K3�.�3/T�3�3���3D�l4fxg3�`3e�3?z�3x4k3�F�3�d�3aq3��3��3�1�3��3P=3�΢3�3D�131�3��3���3��83��3�=P3�%3���3�d�3(n�3>��3�6Q38�T3�aG3�R3̻3�8�3_�k3d�4�.�3&#�3IZ�3�-�3�3D�a3���3?��3%-�3nYW3�'�3$��3,�i34/�3[��3.(�3E}3�ߓ3\��3M3]3e�c3�g3�݆3�3Xa�3X��3u��3�3�Fu3�it3�џ3Ugr3���3�3��.37�4:6=3zuu3ks�2��;4R#�3a��3�K�3"U3�3D��3���3�3#3�"�3���3z��3 M�3;-3��d3�S�3��p3幧30?i3vQ�3]x03�3�"�3ۢ3vƀ3�3z؉3�C�3=�y3�j�3�My3$��3���3�� 3"�K3��3W�30�4#C3]��3�3)[`3�n3ֺ�3��v3��O3��3��3�3�3��33�L�3���3U��3G��3�ɂ3y�3���3͍�3@�+3��3�{�3Y�t3Q9�3Kn3H9�3���3Ne�3ݽ3U�[3]��3 Γ3��36�3+{�3ۭ�3_@4�^G3]K�3�893�:�3.�3���3,�4�f3�)�3��4���3�E�3��F3���3��G3i6s3s�3};�3�qb3S��3�k�3���3=H�3�M�3�ü3�)3G�3�	�3�H3�PU3��3&�3 3*��3HV�3���3�!�3��e3�հ3
��3?s3�֭3_13�ޏ3�ʂ3���35Ց3L�O3�7�3�<4��3��-3F~Z3Jɿ3�B3�J�36��3�(=39��3��3 ��3�Ke39@3r��3Z+�3LT3=d�3�ц3�:s3��Z3`4�0n3݈i3�y3w�F4A��3���3x��3�x]36�3�ޡ3���3�_a3���3`4h��3��3��93̶h3��$4#&�3ݨ�3�؃3y~�3��N3}q4���3Q�f3Q&N3ľ�3���3��P3�~�3"�h3lϔ3���3Z6�3�5b3Bg3n#�3�%�3؍3SH3ea�3g�3<C3C�s3�b3�U�3bM3u��3��3�Gu3ՙ3�4w�l3e�3�W3�v�3�0�3%��3�O�3�!3m�r3Z�4���3+��3��3�9�3h��3Gc�33�4)C3�W3�6d3��#4�<�3)9�3�+�3]��3}�3\�73���3!�3�=�3Nw�3P<�3R��3ځ�3G�3�[�3�Bq3���3C�3T�3G�I3�J�3Cڔ3�]�3�-3@��3?VZ3���3���3��4h`3A��3��3@(G3�!�3��3f4��h3k��3��3�4I�380+3K��3)�a3��)3�;�3��&3p�4��3��3��3h�
4N%�3�ͻ3;ɝ3�w�32ѡ3$��3<�3��3 �3�Ռ3�3��4��3�44�3�-�3���3�k/3�73�$�3ފ�3MR3L��3�P�3�4I#�3V4S�31u�3�jj3Կ�3^
�3��3
"�3B�u3o�A3��3ȉ�3��3�#�212�3T�g3(#[3��31�3jQ�3��b3�4�.�3�q�3�a;3�n4r1�3K&4��\3}ƪ32r3�[�3�(�3��3ɯQ3�4�u�3'aO3��3��3A�<3�sV30u�3�E�3���3r��3S_ 4�9;3]�3�%�3�E�3h�3��U3@��3'.�3��U3�ܘ3��3*�~3���3�4Uk{32E�3�)E3�k�3���3�a�2^��3aQ3w24@�>3a�4ɫ�3Eq3�w3t�3e��3P��3�D�3�/o3�qz3�3���30�'3%��3�K4e�3��j3�/ 3��4�f�3G��3a��3_�D3l�S3�LS32lh3X`J3�R�3�G�3�r84B3O]�3Ϣ3w_�3�rA3N�3Ǹ�323���3��4�X�3@�3K�w3s�3+=�3���3rw3��&3b��3��$3}��38@�3��@3�'?3L��4�4�3+��3A)�3��3��o3�23*r�3��&31Б3cn4)x�3�O3q�*3�5h3<�V3Q<73��3�(83T�3\U3���3I G3Lǯ3�-�3i�3믲3�D�37��3��3SЂ3)8�3с�3K�3�%�3'U�3���3~��3��3*+�3�qK3B��3�'�3��O3pI�3w`u3)�4;�3V�v3�'3��#4��N3�.3=m3?�83�Q3�N3� �3(yQ3��3P��3[Y]3v��3��=3�3<��3��/3QT3?Pl3�Y�3c43Ǽ3M�F3b�=3��3ٜ14̡�3m�>3��n3٭N3�f�3��3!��3�[a3��3���3��3r��3��3���3�C�3���3Ɵ�3�`U3��40�(3JΤ3���3�=53�P3dc3L~3z�C3i��2��2̎�2��&3Q�13��3���2Bմ3�dV3��X3���2��c3N�K3~�3|�2��%3�3�v35Ų3 �3�2N)@3� t3�23��(3�%F3]�E3(�(3k73^3��2W�h3^nD3t&k3I�3�i�2uǁ3�c?3� �3�3���2A�3Gl 3)�3���24e�2��3ε3巧2��2PM33��2)�3j�2$3���2;9<3fb3�3Nr�2�M�2�3.3��*3��%3�33[z34�S3���2jP:3=�%3��z3�A3.�3a�3�S�2�3�3�=�2�R93%�q3 �2�3\�3'�*393�@�2�v3�u_3)3��2X�73��F3JS�2q3� �2;2�2��3���3�>3�j�3�0�2��'3��J3l�"3�I�2!3G�731�n3�>3�03=�{2j�'3��2� 3�f3��3"B=3c�3�+"3P�3�43g�3�t3���2G83 ��2��<3z�2=�"3�[C3��2�38g�3�iO3�Z3���2a�"3��:3u�2QJD3�	�2��]323�(�3��=3Y�2��3�r�3���2��3@�2���2�'3h_3��o3��3��-3�Fn3�i03g��2U3,13Lg%3Ue�2��i3Dc3i3��3�IH3̎�2���25�:3�/�3��3��:3���2��
3ð�2v&3��3�G�2d�3�k3nG393e��2�\=3�x3�3H#Q3�3���2z3���3,�3I�3��2�{<3ƇK3���2 3 �3�3��3u�3�3`x	3�'39�3SV�2A�2��3�D3"�2��I3X��25�3!!�2:'}3:3�3�<3�4���2'�!3D�
3�6�2�e3�S3T`33��2�ZJ3H�3G�q32�%3/Z2=yQ3/~83-z�2� 
3}�2ơi3*U'3H�#3��3��37�>3��4���3U�{3��P3��3�S23+�3IM3��~3Qr�3䫵3S'I3ⱀ3���2��3���3ݤ�2�g�3�G�3W�3�F 35c�3Y#t3@?�3h��3m�3e3iC3Y/r3V+�3H�d3��s3a��3W�l3O��3�\�3
F�3.��3�3<��3��^3T3�UN3��<3z]3@��3�I�3o�3�5�3G�3���37U35V3�V3��3���2�y�37Jm3��3�yK3�4r�y3��E3��3��3��03=(93��n3{�:3��C3�A 3�2�3�T 3�F\3��4���3�'3��L3[�M3�)3\%3�rt3�R�3���2u?�3�v�3��3�=3�3�?k39�33�UM3v�36�37D3�2�3H�;3��'3�9�3xX�3BG_3�yg3\3 �03/3��\3�q3��2��F3'�3\x�3>�p3��2�f3�3Qj3w_3k/30|�3�e237��3F�C3���2�W�3�4s#3�PO3 a�3�yc3C`3a�I3�O�3
�:3��]3��3�v%3�m3#�&3�
�3@��3K�3��m3y?�2aL3��K3�(�3�f3��x3�R�2��4mp�3S��3�BF3�3��3H<K3�ח3}�,3QC~3�z�3�Ϟ3���3O�=3]3�^R3��U3���3�M�2�ԑ3:~-3D��3�_73j�H3��2(�4oJ3$�32dL3\n�2@[R3 �3<3�l3�13�	�3��3�_3B��2BH3v�3��2�=�3w`g3���3O�23Q��3� 3�\3��~3�S�3HV3�?�3{�3o�3�'43z��3�M�3�� 3�I31<�3y_�3{�33�2nϽ3��31z3�:�3R�43>3#*3Y�i3��o3˷#3�3���3�q?3��|3{�3�k[3=M=3�`<3���3�h3AP�3-�3RI}3r��3��34C3���3�GK3���3J��22}3��N3'�v3Ns3'׋3��A3G �3�q3�(V3"�3�ю3�93a�3u�c3��63�53]Z3�̐3���3In3C�3)Lo3���2uk3�3�֕3Y)3���3ʭ&3�B3�83߹�3��-3$�L3�QC3�73��2B��3_y�3Юq3�r53��3�}3�T�3|f>3�3�Ս3��O3�Zm3V�3�3u�3Kn>3���3>,}33L�3��3��3S�63ղ!3\^,3'w�3/\3�Q�3���2��.3�+�3��3]$F3�� 3P�3�Ha3�_3��N3f�3M҄3$�k3Eh�3�)�3  ^3~Co3�Q�3g�53�|�3�M3JFT3�� 3떵3�߭3���2�9�3�h�3��f33!�3��03���3��3[��2�.�3�X3T�"4�j3��38l+3�";3�E�2�,X3��N3��13�1P3 �3kFg3���3Z}3�ed3R��3"41f3��s3�2G��3ȦH3i�C3&�g3��	3�Ѧ3�3�K�30P13�123Q��3/�3��Y3��e3gW�2ZI�3��b3�g"3�j�3o4�2Ẃ3V)�3P�3.uS3���2�3�3�h3V�3�t3�30�3�3�3wO�3~d,3J�e31p3vT�3[�0323A3��<3?�3�3�1�3��]3�?31�W3�2�3�x13�3Y�03Pj3��<3�3F�3���2���3�4	3-D�3_�C3�I,3�3�24�.�2�3I��2��A3��33)��2�@3T��2{g3���3V��3��u39d�2C3�7q3A_�2g�%3�13Nc3��	3��3�p3ϭ43�q�3ߴ�3�S3N'3g 3�f�3YY3�UG3���3��3P�L3Pe�3�/�3"l�3��?3son3���3r�73�9G36��2�dA3qp=3��3c�23��37�(3Nn�3�m$3/.V3�x3��{3���2JA"3g�_3��3��34<�3��3�J3얙2�=(3;H3�=E3��b3�u�2�8�3�?3�Q;3�X3��3yo�3��4d}�3<��3`�3g��3���3‟3��3��39�3V�4�K�3���3�|�3=a4��4�[39�3K�3�*4E�l3�6-4e:�3C��3�"�3�64)4[��3,��3��3o�3W�3�f3_H4���3Gc�3�.L4�;4��3���3ԩ�3e�3���3-Z�3�k�3�[�3��46��3@ŉ35�j3e�4�H�3��3o��3x.�3���3��32��3��3��3�W�3���3��g3H��3���3���3"w@3;��3��3y��3�B�3}4���3fN�3�4��W4ߔt3�9�3#ظ3�"R3ꚝ3L�3s��3�W�3��3�G#4�n�3r�?3a0P3V��3�f�3�7�3�?�3*�3�X�3��13���3'��3Z:^3��3w�/4�]�3T@�3hY�3���3���3�~�3t{�3�?�3*/�3	4��+4E�I4�}]3K�3dm
4�!�3��	4���3�.�3�Nr3���30#�3���3"�3��H4�إ3���3�	�3�H�3�l�3$�3�>�3��\3k��3!?�3���3i�4)&-3���3X�3Č3TQ�3Ϲc3<��3�]�3**�3Z��3"J�3wx3��Y4s�3�ʓ3�%�3�U�3cǤ3l��3��4<��3�ض3f+R4��3��3Q�3^b�3\�3u�337�3J�3ŕ�3�d�3�i	4\ݔ3�3�8�3=aL45
�3��3v��3��3��P3���3��24�d*3�A�3	�P4.y}3z!�3��Y3
|4n$�3t{3���3���3�c�3�GR3	�4��3*[�3Ʀa3ޠV4x��3�3�Q�3�'�36��3�R�3���3�c�3y�4��3V�4���3��3��3]��3ښ�3�a�3�N23��3���3�)4rӱ3_�3���3�.4�Ze3�4٧�3�31�3�r3�3wh�3]��3��4@�4�4���3��4w��3FM�3[��3��#3Nu�3���3��3o��3�3��=3I	�3ԸA3���3�MT3��c32�E3,�Q3f�N3�%13hc;3�H�3�ۉ3P�\3(}n3�%�3�u@3_Q�2��3�F3��;3u�3�<�3��~3��3t�3���3I��3m;�3ْ3=V3��z3��`3$�3�ym3���3E94m@3���3z�3�@84c�3��3aވ3�53�If3�"3#�3���3�{�3#��2��3r�3�7�3 �}3���35�3m%3/R�3>,3+�O3���3L�3	��3	3~c�3k��311Q3��3b3�l�3�a�3�G�3A��3c�3U�3���3 2�3�u�3�`�3�Ņ3_3�~�3ҜD3S]�2uZ�3��3��3��3)oc3t�3���3P�3WhO35�g3F��3<Sw3s�3�i�3}P.3�f�3s+�3��3٪�3�d�3?[�3(Y93�9�3Qg@3�x�2]��3�;�3[x�3��~3W"3
��3]�3�G43b��3��[3덡3�GX3���3d3u�3u�3�(4E�34P3�f3:��3�AC3�3T��3g�F3 �F3b/�3X5�3�T3L;�3��F3��3��	3�43��&3gt3<&j3���3�ց3eÁ3�(3ךh4I��3�B�3o�O3��O3�m23�Ň3Ʃ3�H3�T53(O�3�'�3�Q3�e�2���3R��3��3I K3L43j��31�M3O%�3G�?3��d3&�3:�"4t[93��N3%�&3��3dz3u�F3���3�w43D�c3�#�3�o38�3H�3�Ja3�>]3��P3��w3�Rd3��T3Q	�3���3hd3��3�w%3��4l�3�3�1�3rݔ3�X3�3�g�3v-)3Wq�3F��3��3FǴ3�.:3j�g3�n�3On3��;3 Z[3J��3��U3�8k3��3� 3�V3U�3��!3l)3�]3��t3�I
3��e3/�3X�3�k~3{�4���3�B�3c��2"�3B=o3�d3�-�3�<83��_3n�c3�$�3M~f3=�B4��4�<4Y�3���3�}�3�.4�lk3��)4u��3��3���3IK4�46A>4L�3Bj4{��3P"�3�%�3}�3���3�J�35�4��3�ý3\"4.�d4�3!��3��3y�3Ջ�3�~4Ȭ*4��3���32`�3+O4��3:3�E�3ls�3G��3%; 4D�3z�43��3�Q34��3R��3�r�3��<4��3$@�3¨$4��3��3qѹ3�%4��t3��4s\$4fG�3�ј3G3�3(�4h�3G~^3�D�3�-4�q4�T�3T��3)��3f��3w��3k'�4?�3�f�3Qm�3�!�3Dϋ3��4�f4�k3��4S�4�4���3m��3;��3}��3�939x�3�xF3�]�3�%r3�44C��3!�3J��33�^4�-�3y� 4kb�3���38{�3G�3X�3�ʊ3�˿3\"#4�#94�=�3|3�3�k4i��3��3@Z4 �3D�4YT�3�14���3�p�3ή3�<.4���3u�	4���3@�d39J4��3��3��3e�4Z�44b�4Ǒ�3�>3 �4�
�3Ó�3� �3Vx�3}*�3SP�3B�4��3h/�3��3 ��4��3�|�3yd3G��3d�3���3��4[r�3>�<4�[J4=��3��3�_3(6�3�p%4���3Fv�3�͙3�d�3�{�3b�@4	��3o�3�ڵ3h�94ٞ4c��3:
4�G�3��3�c�3Ɍ�3g��3s��3=� 4�f44{��3�ۉ3��3u�3@�3�F4IE.3Kx$4���3�4u�3LI�3;�3?�R4ࣩ3�3�4�� 4d@�3���3��4�E�3 �4�,4��4���3?3#�3�;4k�3��3q�3ǲ�3C��3�@4��45��3��3
��4�,�3��4q�3���3�U�3{l4��	4p�3+X4�r
44d3�3�nf3v�3Hו3z��3.��3e��3Й�3�a�3�/
46ò3P �3E�3��3��~3��3H_�3� �3N�&3&��3��h3zL3bD�3>��3��e3N�z3Z�73�C�3ה�3��2�33��u3�O�3��3r�3(X�3QW3��36�%4}?3���39��3=��3<�3���3���3��2i�3-��3�U�3�1�3V23T>M3�%X3�73��3��3�M3
@+3���32͊3�x�3�'?3���3��3�y�31�3}�?3�d3�b93 �3eF3��3�7�3披3�s3�Ar3N&S3^7_3�DS3x�a3�3@u�3Z�35g3�AR3�&3��3&t4cpd3���2)�P3�vb3?xt3�Ev3�3�A3ˀ3�Y�3�ǋ3��F3��3���3A%_3��g3Z��3�
3��t3)z%3���3��3�223�g�3���3��w3x�3�TX3с3Dʫ3م�3��@3�q33Ne�3�u�3�J�3C3��B3=o�3�"�3�l3��W3�33��3w53p<�3�y�3b\P3�M3�g4��P3��L37�=3�H3�o�2{�j3��3�3(׈3�׵3̔�3٘3`�'3>�j3|��3-1]3i��3��K3:Ӭ3�3SŤ3|_�3�Lf3"��3}�4�N�3�+n3��A3�+B3Ӱ�3�$�3wv�3�On3�3�3�Φ3?v�3�cc37�3y�m3�o3Y�s3��3��h3�c3g'3�s�3�Li37�U3�@�3���3�sv3�M3
vA3�k3�x43�V3_ts3� p3+��3�+�3�}�3d�k3�k|3�0c3�o3[�	3nۢ3EV-3��3��V3���3�Jp3Bv3��2��3U�*3K�3�u�3)�3�;?3�=Q31�K3��a3:�3��3/ޓ3��t3k�3�ł3�o�3Rgc3[֪33���3�{�3�3��t3�ϋ3=�f3�14�63��3�Y�3-�A3��>3k�i3�,�3��3}��3m��3�ؒ3;t�33o/3��n3��'3��E3�{3b�3���3 o3�43Ȁ{3�3�3�h3q<�3:��3�]3Ҿ�3���3��f3e��3 �r3�'�3Jf�3�X4�1�3�E�3�3t}�3u2�3l7-3m�3���3���3V�;3���3շ�3[�3Og3O�43%�3�i�3U�3�u�3�__3�%�3��3Ɛ3z]�3���3=�3�׊3��F3��3�U3���3��U3`Q�3r��3��@3��4�N3b��3�y3�74y�3���3Sn3[��3��3/}`3ZW�3 �'3%�e3X94ԙt3�OV3��3
JW3E,�3:�	3�(l3�f3U´3�xh3�ި3VB�3�3�ty3?4If'3�R3��3��3t�/3�z�3a��3}�o3�@u3�4 v[3dπ3�Z\3��3�W�3�C3��y3��-3���3c3���3�/3)Q_3O}C3147�`3u<X3�53�nF3̑3.�3���3x@3:��3�P�3��3�b3H�L3���3�UR3� 73
�3�xQ3�V|3j�3�4�3��3U��3 ��3YX�3�+]3��3IK�3ŝ3��X3��3�3X(�3O@�3���3�+�3�*/3��F3␓3� 3��q3%%Y3B��3K�g3;w�3{۠3/:�3��2�,>4g�n3l�3��739}U3�֗3�6�3U!�3�xw38x�3E��3[��3��?3%�93h�3��3�7F3�;3V�3P�3}+3��3��3��}3�n�35B�3�K3X�d3��332��3^_3�ׇ3��3�o$3d�3��3(�3%�3rW3�'�3ut�3��43`߰3W33藡3�z�3�y&4:y�3�T3�:3��-4P��3A�)3��3>�&3Gl\37~�3v`�3KI.3Lڇ3��3�3�l�3�-�3�3S��3�7I3�/�3(��3��4�A_3���3��3�X^3��33F943���3\�3�p3�u3��3O��3��3�3���3'®32�3"w3c6�3De�3{�3L��3R?3��3�3���3�؁3Ơ�3��[3;�3��3+63T�=3��g3o��2�[{3 C;3�B3��S3?8�3��l3��D3��r3C�3�3�<3b�L3�53]'K3��z3@��3K6o3J�3IƸ3=��3LG3�L�3TX�3|��3�3��3֖�3�p3��3���3`@~3B��3&��2�@�3:��3��3$��3C0i3?F�3R�3d��3���3_]�3��m3�1�3��c3OX38U>3���3�xr3�w3Zt�3�N137:�3���3��3>R3��22ZL3\}53h#@3{m3�I3���3��U3�ʟ3;CP3i�3�p�3�Q4��k3��I3��[3�[O3P(A3��3�+z3d)3��3�e4Kt3oX3"C3�3�3⒞3Y�:3�kp3���3�wX3�t13�2�3Z2#3YH3�O-3C��3F�>3�^3�_u3�o�3J�3g��3�@x3�(3\�03���3"��3�J93i�2X�3�	�32a3�[�3TTc3N�v3��,3@ߊ3f�h3�Y3% 63��4t��3}!n3Xp3��k3�3�c�3.;�3��2��23F��3�մ3�$�3��3
�3*=�3��I3']�3�/3rђ3Ä3�x�3al3�J�31�>3���36�3X3�w33��H3R�~3�%^3j+�3\�_3Fm�3��4L��3�ʇ3)n=3z�3G`3|U"3^�3LM3���3�r�3 ��3Hpe3	��3�03Y��3ܠ3��N3���2yy
3�!�3_fa3,�3)�-3H��3�4�؏3��v3��3���3���3�~t3�j3=�C3�~3a-3Q��3�KP3U3�b3ͻ[4��z3�F�3�)k3�{h3��/3ɟ3^U.3���2�7�3�3rM�3.S3V�C3e�3�ZB3��^3�Ҡ3��2��h3�&3�Z4��C3�a�2|3�]:4�[3
y?3 �3��r3x�3"�3wFa3%t13���3���3/��3{�3 03�'|3#2�3}D3�0R3E/3 ޾3�"W3\j�3��3g�3P�3��3`�
3��P3B�03?*3�3Go3���3M�T3.�@3ך�3���3��3���3'3���3��3��83�FV3/?3��2�P�3�C3��e3/�H3�c�3Z>3�|�3�3D3sl3��3k�i3挆3���2{�33k��3�)�3�Vc3}3��3'3E3�r38L3N3�U3�Z�2�B�3p��3!p.3�e!3{��3=5�3ÇX3��33�73�8�2q�(3��;3�)3��`39��3&��3	h`3�?3R�3|n3���2��Y31�3w�3�3F3��t38�L3ni3#6J3j�3�(3ޫ$31*X3�{03�v\3zzV3l3x�3\k3���3\|�3��e3/(�2�R3Y��3��37)�3$&3�f�3X|I3k��3�Xe3?�13%�y3���3>�343��3;Oy3-�3��3F�3��:3��e3mez3�ݡ3�S�3@�2���3�]�3�fk3Χ3GX�2!��3�C~3�83���2�3tT3���3UC?3��~3��43��3/ L3z�3���3��2I�,3tB�3���3�>3�}^3�{�35(�3�3d�3���2�h3X�B3�	�3
3}3X�*3/�3p��3�i3���3�L(3�b�3N�3�Z3�R3S3-�.3dM�3\�3'nl3���2s�u3Xvm3��3��o3��g3g�3H�3��3���3K��3��/3�3��@3�o3F�C3_�C3>�,39UK3y9W3X`3IXH3׫�3�n�3g�3W7;3��3�?�3��3c.33�(3��31�C3���3JY3a�3�,3X��3�A\3:b83UT�3�})3��	3Ρ�3�.�3�$3"|�3�N3�;�3�_Y3�	K3g��3G�z3��Y3D�<3�A3��63��
3�B~3RY�3��:3�3���3���2_�r3�j3�n?3R�!3�&t3S�3π
3Ԕ�3���3�K�3�]a3�t$3��3�
3��/3��f3Um�2�{M3;M3.}3&�"3e��3a$3��3M�j3t�Q3��t3N�3�X3ٜ�3)�:3{gh3�v3�G�3��3��3��&3H�R35�\3��E3X�3�Վ3d�f3a�3�ߢ3�8�3uj3ϸ�3�X	4��3t�3Z(3!Zh3h��3��3��3��G3P�3|�3�h3զ3�37��3��
3���2P�B3ﰼ2�˝3r3A�3~��3ƙ�3�^ 3��3��p38�l3�B3Fl*3�v�3.?3��x3kt�2�)l3=�3}��3׸�31��2BD3�![3�Y3�[\3i�3V��3�34w�3{�p3��3�3u+�3�.3�B�3Ү�33NO3	OU3�Z3���3��3'Ts3i5�3��3'3�f,3H�3]�!3�3���3�@3�'3H�3a#�2jtF3�K�2��"3�3�e3���3�=3xD|3|T3+"�3铊3�O3�ex3���31/�30��3r�(3��3�~�3�x3�+W3���2��t3�3Td�3�_r3޿t3\a*3��L3�j�3d3^3��Y3�J93Z�3�63V�_3�b43K�$3�9�3j��30^?383P�83�¬3��@3��~3�#3|D�3��Y3�j�3��:3�WJ3��2|4���3� �3�.3�� 3y�3���3�j]3��F3w3���3&&�3��13� �2�{3r�j3��d3Γ�3*��2fN�3�3+�3�8�3��3ӗ-3��3L�l3�n43�Iz3��3z�H3��@3��p3E�3�>�3��3��{36��3}��3�u3��533ݼ29� 3W�3B�d3Q3���3_Qp3�%3�o3F�3r�3���3E�i3�c�3���2EJk3�w3 3�.�3럕3���3R��3�E�2;S�3�d?3��3���3~�35��3�̂3pЇ3�23Y�<3%��2��3=e3�93���3�Ʌ3h%3<IR3:p3L��2"�^3~'�3q�3�z3Թ3z	�3$|3ZL3��3w�3p2d3C%3��\3S�3Q�3FUj3aG�3qvT3U�#3��3��U3g3�*39&:3'݃3�Q3Ý3�Q�3 Ť3��2�AR3W333MD3��\3���3n,3�M3�c*3���2��s3�D�3�NH3菔3�3=�&3��3n��3�V3unr3n�3N��3�S�393��2��w3X�Z3'�f3}�^3�2㳔3�53���3��3��H3I�s3#�3*3�2\3}�<3�B3��3��3�h3M�3A�O3��3}KR3+Y3RW3�f�3?QP3҄37�O3���2�N�3&�13Kt3�.3� �3�ߒ3�\�3r3��	32"3J�_3��.3Ն3o�3^3�2��g3�'"4Qq{3�C'3)6�2>��3�EA3�^t3��|3I�3<b�3Fz#3��38/�21*53��@3��4G�A3��3~3H$C3V/�2E��3�P3�2�!3R��3B �3�� 3P�2�ld3PD3�2��3^�3��43�s�2��B3�x@3 43�F3�B�3�̛3�b038�!3�7e30�A3\�03�"F3<�336lU3��33�|�3��"3#Ӏ3n;�3��/3Z�~3f��2#�3	@3�s[3��%3P23B��2��3��3W�-3'73�,R3n� 3zA32`�3�'�2�o�3 �3`�m3�zF3�k�2��a3#�u3���21��3�.�2� 3m�^3_�3�}+3Jy23�F"3��3)��2��o34S3u`r3N~�2r{�34]�3��3g�3�]�3�3�؍3��3"(�3|3C3!3�E3�R#3�t]3?�4%�[3�d3h܍2��4/�3��B3��G3��l3>l3�H3�qe3x=3mC3�Γ38�3;�b3�"3�js3�/p3��3�B3v3�ݘ3��(3	�f3��-3�Z�2��&3Ό*4��b3 \93�;�203��>3�m3�6i3�?3_�3'@�3��3�3m�2��3�;3qH�2C73���2[Ξ3�X3N��3�bs3��3��N3N8"4@�|3���3_V3�C�3ܰ03fr3Hdo3�Mt3fz(3ݩ
4!��3q�3�@c3��G3}݉3�L32��2���3���3�%3���3%+�3D A3)�3Lv4y_H3�x�3<��3z\83�3O�3k6�3��(3ʐ)3=z�3H�3�3��32��3�S�3T�%3Ђ3�,�3��q3(�03�+�3`�3`_T3W�3�w�3�W.3�3�6\3�|�3�z3�#t3$'�3��3�c�3H�3�\`3!s�3հM3�(i3j"�3j3"�3�3��]3w��3���3A�{3봫3&�3���3��S3��>3�w�3�<93k�3��3O�3l�3�a53�R4e؍3�K3�gV3qg�3D��3lܚ3�rM3fg3F��3�;<3�a�3cK93�~]3*3�V�3��E3��S3{-�3*|�3�3��3��3}��2�֑3{��3 �3U��3jr36�3HHE3�%3T�3��3c9�3B�E3B)�3Xpa3鹌3!�@3v+4��M3��b3aA3�g:3�>E3���3=��3DQ53��z3DS�3<�3��s3.|32�3r*3!!/3�3�w33π�3~�`3V5T3�;3SK>3U?$3��44$]3�K3�&q3|�O3��?3���3L�i3#\3$~�35�4q��3��:3�G�2ޑu3I�3�_\3Ǜ�3��[3�{3�e3�Q�4^3G�F3��3d�4:X3@�l3��3tS�3�.3 y3��y3]N3Ъ�3�c�3]�3z��3s-3��S32"�3�)J3��L3q;�3���3�:3�3��c3:h3��H3�'�3"�3��3=�q3h`3�z!3~�m3 ��3_�"3��V3��3b{3d�y3��Q3��3��37��3vk�3��2,��3��3�:�3�Hh3��e3��t3�4�(3��A3� Z3~��3��X3�e3�!�3��$3��K3T'�3od�3T
3%/3xF�3K��3�;(3�b�3ѡ3���3���3�ۥ3���3�A�3Z	v3�D�3q�j3��3��3�}�3��o3=v�3�ݻ3��S3���394�35�3+>�3/�3���3n�4�5�3qu3b�~3+Gs3�7w3��3��4�;�3�0:3���3�و3� �3�Ew3��3;��3׳31�3dC�3F^�3}��3��3 y�3]�	3~e�3��3V�3��3��3oy�3C�33�&4��a3"��3���3|l4琐3\��3���3AS�3��34z�3K�3?P\3��3���3���3қw3�ʏ3;��3ٵ�3X�3�~�3�j3"�3*�z3�s�3��3��3�q�3�f4��b3t��3 ��3p�p3���3aI�3��3�\�3h��3g�]4sO�3��<3�*3���3uz�3YQ3�$�3j��3���3͋�3m.�3jØ3��L3�?3��4?Tg3O��3!^�3�T�3�*3���3IW�3��3@V�3�ծ3��3Sh+3n�A3���3:��3E8�3	L�3:P3�?�3�^3�� 4���3f{�3h �33�4N��3��3"�3[��3;͗3bƭ3
-�363>3ݶ�3_� 4*:�3��3��+3<�3<904���3q�3P�3���3D=3���3vJ�38U3��93��P4G�3ki�3h�3_d�3O@J3�Ѥ3���3��j3�@�34%�3Om�3�Q�3r5B3�?�3��3I9�3��3�73g/�3ہ3%}4��{3m��3`dG3��4�+C3n��3���3���3�G&3�;�3�49E3���334e��3�k�3�/3DX4⑈3��.3���3�3��83�>34wB3۠t3�Ft3��G4E~~3(}�3�i�3��O3�t�3L�3���3��53��3�)4�h�3�}�3L�3���3�i�3 J~3�3�3!\R3�s�3�eu3Ǣ�3-�38ڮ3��Y3_iC49z3V��3	��3 �i3�i�3��3�C�3��33S�3��4'd�3�|�3 �3�$�3�֭3��k3��3��3���3
W�3
f24��3���2f3�s�3u��2�߸2/i�2��2��2s��2��3�$X2ح2#�
3TG3��63���2��3H�2e�2���2�_3e�2���2�73Y38�3��3P�3�`3���2J��2E�J3v%3��2�F3 �2v�3mj3.]3*�3��2K�E3�(3k��2�3�$�2��3��25 W3��3h`�2 �2�9�3 ��2��63�Z3�E3�m�2Ն3��3�3���2w�(3�(3V��2���2f�3�73��2�P3Y$�2l 3郲2&'3�2�2w�#3���2W�L3t��2��(3��3�Y23�2�G3!��2��2�q3� @3�;3Mr�2B"�2�#�2τ^3�3 ��2��2�Jf3��2��3�r�2H~ 3��2ys�3\�3+�2�2,3���2s��2��43O��2�j	3�z�3�/3'E�22��2��@3�W�2d��2��43=��2���2>��2tN3���2X��2���2��L3��3�-!3T�33�y3�A3O��2��f3Z[�2��33���3�Q3�V�2L|�2Ŋ�2�]�2�#�2���26/�2[�73�2ʺ3>�43UZ�2Um�2Q�3\��2R��2�J�2}�3r��2�:3�x3bZ2~W�2?�3An3��2 �2���2F�3�:�2��3�1�2z3 �2=J3ͤ�2�#�2/�2'6I3���2YU�2� 3Iԫ2#g�2>�2�g3 3�3 �M3gTI3��3�L�2��V3�3b#�2�" 3,��2<<�2+�e2�V3O1�2uk�2ۨ2��t3�2G;53S�{3As�2'��2��2�H#3>�2�D�3��-3o�23�*3���2�/�2�6D3s�2R�3�3�2T93mv�2$�%3��3mX�2`�^2c��3"$)3}Hv2�I�2�`�2��2�B�2'��2��2��2��-3(�3��2�P�2�Z23gJ�2�K�2� H3EN�2zU3�N�2Q��3g��2���3*��2���3'��3�v3���2)�<3,��2{��3��p3�3ʢ 3�]3�R3�P�3�P3y˵3L�3�%3PI3N��3㑅3e��2�ӑ3�f23
:3ľ_34��3�H�3�r�3��<3�vZ3��z33�3�^k3�0�3�3�K�3�:u3!��3�R�2,�E3o 63�X3к�3_�3�{"3P]�2R��3�23�e`3a�@3�[4!�+3=3>3�AJ3E�2�#53��}3n!3��	3��35��3��a3h3�
�3A��3J:�2�On3��'3T�,3�!�2Q�3ػ!3��3�	3���3*�N3cc3@��3��o3��3��W3moZ35�3F�f3|$�3�g3��!3��43��3�3��^32H53s3�%�3n3��3��|3�73Q�3\Ѻ3~�~3)��2{sE3��X3rG3c��3��3Y5.3oA3`%�3QRc3
�3W�3}��3>�i3��l3�,�3Z�S3l�3H8D3���3�&�3g3o-�3�	4RK�2^Ɨ3��u3@3+3;&F3�X3�#C3(3z�(3UX�3\��3�3�.63L�N3��.3�&'3��&3��3�t^39Ox3�<G3��3i�3�r3^ה3}^F3
�3/y�3	E03M�+32A3�c|3��Y3+�3T\�3	�|3m��3��37�Y3�E3n3b_3G�+3��Y3���2y�k3Tvq34�?3ٺ3���3�rT3�L	3�r3ʹ3�8!3BB3�B^3~3�\3�l�3�c3�X�3��2�o�3O3>3�V3�^3'�>3ڈ�2F#�3��?3��83ٟ�2��v3��[3��3�Z�3:�3O*3d�x3��3��3ƣ�3;�o3ge3��q3<�2x7w3�3*�+3{=�3�+�2�Й3S��2��U3,q�3���2���2��(42��2�Ŋ3��/3�I3A�2�̓3F�3�S�2�/�3�xw3��k3��3���2}�r3'z=36��2jf>3^~3L��3%x93803��O3���3�%A3"�3*^/3�TM3mH53��
3c�3�F3L��3a�H3.�3!}4;��3���3Q|31]^3���3���2��3HW3VL}3���2�J�3~�3�ʹ3n�n3�d�33_3��(3��3S�3�2A3��"3?o3 31�Y3��3j)z3o��3>3JZF3Ȍ=3��2v�3*&3\]�3ڗ�3ƒ�3�G*3K�3 �3h�3b�K3��~3��=3��3f-3373^�b3Zg35PW3�6�3F1�3��_3�.�2�ߖ3�o3�f53��R3�Y(3wI36f:3s`3s3��3z��3k��3	r*3oht3w�P3� 3�o:3��\3�n�3�KH3z3���3I��3-\-3iw�2�xr3F�2n�-3x�'3��13�YQ3�3M�~3qTK3W�3B��2�A�3F��3�gB3&��2�k,3+�c3���3��3ƞK3���3k�3R�c3��2�~�2���3�|�3D�3��v3u>/3|>=3�+3�r�3r�\3vuX3�P�2�,�3^a�2h7B3� �3�_3��.3�3y�Y3�F3�
�3���3{%�3��3�_ 3='s3k�3�hP3��3:�.3$ud3x03ȏ3�~43�T^3�`.3�3v[G3u{3r�3�ދ3�he3��33��3���2��)3�3n�3CB3���2��y3�3�3�#3���2��v3��23�"�3n�>3��z3is(3�1�3�X3��(3�53��M3�;13f�L3}͎3�43>�03���3#�o3Mp3S@�2�`3K4G3cEg3�
R3�5 3���3�A
3�T�3�m3?3�l/3B<-4I�3;�.3e��3�M.3�n3]3D�e3z�J3ˌ�3 ��39�3I8V3LMH3<X3�ُ3s�D3,
23s٥2裑3���2ڊ�3.<A3��3�<�2k�4p3�JE3a3V3`	Z3�e3��=3�2PjX3lNv3��3�F3���2�Es3Z�G3)��2-�3���2�1;3��3�}A3Ù�3_`�3���3�X�3��*3�	3=��3t��3/�3I��3��3��
3�<3��3j��3#F�3�9c3�4���3�3�ԛ3�	�3a�3��]3��3Z��3q�3ͱ�3�P4��s3��f3v��3,}L3�؎3���3?�3H�13�3��*4Ć�3��3�S3M�3v��3
��3!{a3�k3I��3+��3v�39��3	��3��y3�4�3�-x3�U\3M3�3� �3J#3wW3/a�3"3Xӏ3+��3���3Q,_3��93�]�3{b�3�H3N��3$�e3u֨3Jn�3G�4���3f�3KwV3�J�3چ[3�ħ3E��3��3,��3��~3j�?3�@�2�'t3+��3x
�3�X3޴
3k�3�w3ި3o�3f�F3��&4��3��3"]�2vo?3� �3�s�3�w3:Cl3u#�3�G�3!��3l[63�,�3�y3g�3��3Kث3��3Ut3�[�39X3\��3?l3�7�3��z3��3{U�3�P�3\��3mmk3@�3��37�F3�e�36q�3!�n3N�3�d�3�3/߆3�3�3�$�3ӫ�3�P31�S3���3��3���33�ֹ3��-3Dӓ3X�e3��+3ŠF3=4�ݳ3��3��63]|C3V<3b�r3���3�Y+3JC�3O4�d�3��h3�P#3A�	4�5m3FB 3��3���2|*�3�`3cl�3J��3�J3�4'3��(4⮗3���3��t3�63� 73�H�3ѥC36�3� �3L�3�޶3W�3g�+3yp�3*?E3�A�3��3.3*-�3]�3&04�z�3�Ub3+3R1�3�Nt3 �3kt30/w373خ,3X�3���21α3���3N�3
�3��,3<c�3��~3��)3#��3��|3tW�3�%
3�P�3#�Q3Q�*3�"3|�Y4��h3��f3L�3a�w3a]_3�Xr39��3 �83H{�3x�3���3�LT3���2�֬3>�N3}h*3���3�D3�/�3S�3�|3oA63�e3��(34��3<�+3%l'3Ǩ.3U܌3���2̉z3��53
K�2e&(3��31�$3i3�XD3�d�3'ǆ3�hC3
�^3�x�3��3�d3I��3V�34�*3�.H3�u�3�^/3�&�3hQ3��u3h�I3�@3{S�3�,3�؀3��3��3�}3*93�&{3h��2�QE3_34�f3V3T�F3p�3��d3tRD3Le%3�Q�3� 3�y3	�F3g�^3=��2�,�2��?3jv83u�G3	s4_^3ʤ3��2�U3JW3I�3buO3*I%3nj3�(�2%��3�3:83��f3�Y�33�(3^'�2�AD3�23�I�2��A3��3r�3�"/3z~�3?�w3��3��2E��3{s@3���2��W3�3(-3a�3��3��z3��,37�3ξ�3��E3h�3ڿ33�X�2��>3e:b3@��2�KE3�;�3�Ŋ3�Ä3`��2�Y3�4�3V0 3�P*3�w3t�36P/3���3�=�3��=3Ӊ�2���3�3��q3��"3���3��A3���3�{�3W�3!�3�b�3��3$J3��3��3x�3�~3U��3�&3{�3yO/3��3z��2j�>3�rZ3��4�73�3|3Jv�3A�3!�`3?m�3�3��93s��34=�3�3^�3��c3�(f3��%3-g�3W�2�aI3�`83���3�)3�NW3���2b�c3lM�3j�P3_m�3��Z3�1Y3��P34�m3��M3���3��3L��3��53
w63l;33k�3.�3m=t3r�3V�#3ӫ%3p�4�3,��2��"3d"�3�BT3�h3]''3%m132&I3��2=/Y3�N3���3���3�r�3]Z�3���2,	,34y�3�/73Ռ-3�p3��3�j 3���3/�(3F�3��z3+n�3��2�v3!-3��43 �R3�%30�/3��3J�w3�ӹ3�B3�RS3�{�2R�83�L�2�#3�	3���2��b3�}3�Ō3B�N3��33k��2��3C��2�0I3r��2�(T3�L�2��43I�E3���2�3��3\��3Pq38��2Xm33N03�G�2�853�#3a�A3��2�fp3F�=3�`3�L3�N�3��M3ý>3��V37Gt3�5�2��&3�ʱ3'�-3n��3��z3�^33ـ3���2F�D3�	3p��2�<�2��`3�>p3��3D��3�?"3J�3i!3d�3Zz3�� 3��i31DA3Ο3=��28{B3��$3�s_3Dʹ3ݿ�3l��2�3|53]"3s��2D�<3&�3�Y�3g�13�\g3��3��d3��13:�3`�m3-3��X3�^�3���3��Q3��g3���2�e�3;l3��3��[3�I�2�J�3�h�3Ŀ?3�|3�>�2��m3�']3��3��J33zÛ2h��3[�3�	3��Y3j�2�KL3��3Y5k3���2��X3�A�3N�3��Q3���2�33�;!3��!3�_3��2� �2Ĵ13�C�339-3�
3��@3���3;�~3�C)3�l3'�!3�!3QyF3��3�3�R3+�3x:�3��@3��	3�w3��3.c?3��q3�*3(^W3�03QC3��G3
�53��2,� 4
��2Ш"3��3'�V3j�A3~3�Ξ3`+3��3��4��3�3��,3�q'3�13r1�2�*3�2wNU3�93�fC3��23�%3s3M4�D13N&3�C�3L��2�_i3��3��Q3�3;R�3.��3@n3FVG3t=�2��83��3�3G�n3�\�2ݏU3�&3���3.;�2�}d3��3E��3A3��[3o9Q3 Y3�(3]$3H�O3{3�@�3�P�3�~3[?3�
3[3%�S3�"3jB3���2j�35��2*�'3�'_3W23�v�2 �3��3+�~3�Ѕ3pZ�2zc303�N3[J�2�63���3Q��3E�3�	3B'?3�^3�o�22�3��2���26��2�d3x83��o3��v3P]r3�s�2�3�3F2�3��T3��3��U3�h33a�,3�w�3�S�3i�3�t\3��3�a�3�q"3[�;3|#�3�p3�
3�/�3�3�C3�E�30��3t�33&�b3��3�ǆ3ُ3^SR3�!3Ub3"i3�R�3͂u3l��3+Q�2O:X3��3���3]3,��3��73�[3��d3��Y3�j3�r�2ڻ�3H�3۾�30��2���2�'3).03�y�3�23��]33T�4{f23́�2�X|3��32�+3d�3δ3t�3�3]��3�sw3p�d3u|
3^ߧ32��2� �2agB3���3b�2�F3�g�3��!3���3�4�3�/�3���2�F�2Iz�3��L3��2��F3�#�2BՈ3�t3���3�C3Y�3<� 3��3\-3KT3�'?3���3|l3t��3o�3��P3��^3�3q�G3�63�4	3���3i�\3���2t{Y3�+3�zd3��83g��3A03iGH3�3��3n��3��-3Ӽg3�M�3�L�3ވ3���3a�;3 Z3�{3�IQ39� 3��3��3�:3ҁ2��B3�\�2��Q3�=�2N�3zS�3!�2C�30�3r O3~�!3Ֆ3��#35��2�=j3D�G3�i�2��;3�9�3=kJ3��Z3�V�2�3g<@3,E3u�~3/L�2�s�30w3Mă3�4[3Q�^3�(3�2�3&e3�d3;s>3��>3�R36A3�\3���25'3(�3�9�3�>F3��2�b3��p3Z�2�N&3*��2+P�3I�2��|3F�3Uv3�Y3�T*4��3e�H3%b�3n��2���2T9|3�
A3D�2ء�3�r3#S�3��q37�3���2�ތ3W�3�<3��3��3Q3�@a3_�}3��3��#3���34��2�[3�3��I3`*H3K�<3Y��3�� 3P�;3�(\3�+;3_��2�;3�9�3V	3��'3'M�3IrO3��13@%i3BM<3�T[3���3o�13w4��3�<3�BA3�w:3�3��3�2F3��93�[�34	]3���3��3F�N3�J�3树3�-?3�e3
�3�Y�3i�2���3�.p3��3
�x3���3#�I3�J�37F3��.3)��2��j3��3Y�O3ƙ\3��3��3�?�3v�3=e3^�3櫴3��33�n36�;3�Z3��T3�r�3rL�3Z8g3��3���2RD�33�M3��3�fL3Ma3��3:~_3S�<3
�4���37�p3x3￁3kX�3s3 8�3�s&3o�3k�3��3�d3\��3���3��3΃�3S�3�M�30Ҋ3�aR3)�g3ou\3�}3re�3�q�3?��3�q�3��S3���3Y�3�[;3��3�ʇ3�3t2�3rn�3�>t3r��3�U3��4�3��>3��w3�;3'U3C��3���3�3�O3�
�3��3Z��3c}u3�)r3�Ü3a�3��k3�c3d�3��r3��3�pF3!j�3��3&��3�>o3��3�ih3��63]t(3��3��|3k�2eޓ3�'�3g�3� x3�3�\A3|ǂ3G�q3�Z38�22�z3�F/3�<�3�13�Ө3�RL3!4��=3퍔3:݌3�ή3�	p3�Lv3�Tt3I33,�%3q�4��3�93�Hy3A�J3��Z3��x3`d�3	�3C8�3�4 3�
�3��V3~��3���3l
34�*3?b`3�F3+�k3��63�TQ3��3�/�2�^Z3
��3���39�*3X��2ם3��)3�Vg3�.]3�3�z�3q>3(��373lB3U3#�3Y^13� G3�L^3���3��)3�sv3��3��d3d�|3�X�3E^�3��f3]�3�O�3]3�-3���3G��3�r3X>I3ӓp3��$3]s3j3�p%4J�83�t�3�V�36nC3�:E34"�3�t�3�y3�r�3���3��3j�3��3@�3Ț�3��%3	��3��,3���3��j3 p�3�<3yo�3>xZ3K0�3��3F��3�O3�34�3�3�3��3<?�3z��3P3ϲ�3�s3BN�3 �{3�Q�2&^=3���3P�3?53^��3�F�3J�`3m�Y3U��3k J3��3�W{3�
h3�|U3u�3�r�3ő�3d�39��3,��3Da�3�3��3Q��3�/�3v�H3��>3��3���2��3���3jD�3a�3�x48�3"�3J�}3ۃ�3�y3�Z�3�,�3��#3�N�3��3
4�3��3�w3Yث3	��3�J3�+�30eY37P�3�_^3��35��3�Tq3+yz3���3'�c3Op=3y�t3V�13a�z3�Մ3��3V� 3���3��3�3R3��2c��3�v�3��x3O�3.�I3�0�32}t3H�3�N3.13؂�3�
�34g�3=��3(2�3і~3A�3�Qf3qo�3N�3P/D3�P�3*�3�ZP3�@�24�K3x��3��3�W�3���3�Nh3��#3�3�3��I3n��3��37��3���3��J3}bl3֣3� 3ome31��3
37�H3D�3��3M�3HuZ3��3)��3Y/U3�%�3!��3� �3��23l��3#�3��A3�S3��L4��-3 n3l3�h3͏L3h�33~u3��3B73f��3dM�3��G3�3�Q3g73���3��X3S�F3���3�\3�3�QJ3W3ԍ�3�#4a�^3���3�32PS3�FG3'_�3K��36.�2��3�2z3P�3x��3N��2���3!�s3T�3��4��2�^�3L�[3�$�3\�%3yɩ3)�3M)M4S��3Ͻ�3n��3Zυ3F�t3n��3�q3�%63�q�3�@�3��u3l��3�I,3��z3�!4�_m30}3�ܛ3��4�3O3Ϩ�3��3(�f3s�*3��3�x^3�M~3
�K3Bv�3��13.V%3!�3L3E��3���3��3�^�3$�2���3p�3%+A3���3��3�N�3y�m3�r�3,q�3&C3��	3F1_3�)�2	373r�t3���2��*3�rA3��3A�G3���3��m3
�3]�3�I3)m(3�?3v��3��3�3��2���3��33�P-3�;3���3-!3_�A3��2�(3��!3af@3�:3.�3/�W3��@39Q3Bf3�Y�2x�@3%��2���2� 3/0 3)�A3��3��"35J&3��m3(T3��E3� 3��3�2�3��2ޚ3�35�
3AN�2�<�3C�:3� 3Mex2�E3nD03˱2"3v�w3��53c�2H\R3S>3��=32�3`t�3�(�2C3�nv3ǏQ3�2��3Sh3\��2�s3�hC3�#f3i�S3�3�=3�j3j�2�M�27�o2��53��2��+39a3�n�24�<3�r�34]3�'Y3�2���2�R/3�3m�O3���2З�2�[3I�y3�|�2���2��03�h�2��28�3$��2eq:3H'�2P�Z3�];3�jJ3�(F3���3R�$3��3S73>3��13`3�73b��2��	3��3�Χ3[53(3�N3>�3�f3:�2�pG3}03���2�F�3�3V6�2z{!3BO�3z�3�N23qr)3V�37�3�t�2��z3|�73��2��3��@3��2��2U�;3�,&3�n<3J�3��2P"3H3N��3�{
3=}3��2u��3��2T�I3@��2�8!3���2�K>3���3q��2f�3�G^3n�T3��T3P�2;bM3� X3" �21X3N�B3l.3�C�2-�l3qa�2m��2�DO3��3_53�&3�U$3!�23��'37�`3	1�2��D3pi�3q�]3�Z�3W�2X�73|W*3ms3�l:3w3�73&�3�%3���2�=�2��2�u�3V�3UM;3���2B3���2�3��3���2_Y33v"�3<�13� 3���2��*3�X�2�ͷ2Rxl39��2m��2`c�2���3Qo$3��v3�%23���3`�3x-N3��3Q�!3��33�N`3�ږ3	��3��3�p�3�j4q�3�o3�93n��3Th�2��13Cu�3�3�63�K�30{|3/��2�N3��3L"�3s�3���3�?3H3P83 :�3��E3}�N3;��3�38�3��
3��\3�yE3]�2E�k3Xq3q�c3G�'3"�3LD3��Y3�>&3ۨ�3�lF3�P43�h�2ւ�3��3�!J3��n3;��2��3$`�3���3uMb3���2�zC3��i3��2�|�3K?E3���3\Q�2��3�O3�G�3$
O3�b�3�(O3��e3��/3h�K3��\3<y�3�2�3�8@38h35�33�3`�3L�2�Z3wn�3�s�2E:<3S3>}3R|(3�<�3�Fi3L�;3=�2��3�G�2qt�3�3f�3��3��\3�]%3^03N�*3�M3��3��83#��2)G�3o�23I�3Bi3ZS�2��53v�3nS�3na�2{~D3kԎ3z�3$�3��o3�8D3�`3M�;3�43H�3�"�2��\3ҫx3�3�#�3U�$3�U�3n	3��3�y�3��2Y&=3A@3��J3��Q3&�3&�93�4��3�w 3��m3c�3Su�2Nh�3SfM3�3AQ3��|3���3��2q�3�d3v43�U`3��M3JC3?�,3ur�2o|3�>�2;��2]�3Z�3�3�3��3^<3�dV3�Or3n%R3��A3��f3�3kK{3P3�Q 3��3t�3C��2�E3�-3�|!3� K3�VH3s�3�3�SW3��3��3,\3m{3�p�3��3�l3s�l3�i3{��3�ۏ3)��3�=C3�* 3�63<�3(�k3D33�?:37`a3	�Z3jQ�3!q53�m�2�3�2���3�35w3W�93�3�%$3
3$93߁2;�J3J�3�k3�i3��3��3��I3Wk�2��A3k��2���3B�2_�3q83�4獌3FO4���3`ğ3@¢3�p�3�q3�q�3�U�3�'H3���3�T4�;�3��4�ѫ3gm�3m�n3�43^��3W�3��
4��k3�u4�Y�3\`�3,d�3��94��3���37��3!y�3��3*�3�d�3u��3�Ѯ3�v4�#4��4��@3��
4"�4t�3���3�i�3fF�3���3��4�v�3!m�3�M3,4ΐ�3���3g�3qc�3�:�3	�4�4Rü3��3)$4u�"4+��3g�3o��3�P�3�w<3�t�3O��3���3ĥ�3�14���3]	4o,�3{49y4T��39b.4ca�3�&�3�	�3s�3�i|3+��3�W4c"�3���3�5�34��3�Ĩ3|�3獿3gp�3�)4,��3La*4%ז37�3�km3�*i4�3�]�3�3�P�3�_�34-B4��3��4��R4S�847�3��&3#�3lN"45bN3�X�3�3�U�3�@�3_7
4�h�3	9�3~��3-�4@��3�#�3��3��4�3�3��384`+�3y6O3��l4�R4��3~�.3���3z�4D�3L��3X�4P�4h�3h��3�փ3�Դ3uU�3�[�4��3��3Ww�3���3�X�3�y}3]!4��m3�S�3)@G4�=4��q3��g34�j3���3�B�3�s�39�3���3 ��3�j:4ZV�3�U�34��3=B54�p�35Jw3(�3�$�3�=�3�Y�3Bv4d�i3���3U�4�"4��3�D�3�r�3��3
�/3�J4���3�r�3ك30v�3��3$�s3~J�3�ld4>dJ3���3��3��3�d�3�3��3&�i3'�3<�4���3f3�3_��3u�3���3�n3��3'�3��3u)�35Z4e!�3)(�3(�3�4���3���3q�4�o�3��3��3��3��3r�4��4ĭ�3�=4���3d&�3�w�3C�3eM�3��r3d"54h�C3H�4�<4P��3NN3hD�3}�Z3�L�3�&3�03�M�3I�3�3�3>.�3m�e3���3��3�m�3f:�3ȗ�3�k63��3o�+3�e�35�
42�43��4���3��3��3r�38&(37�3ɍa3�=v3b�3l�|3i}3��E3GF�3���3���3���3P�3�ޠ3��3��Y3�{�3�3_�K3�@�3 W�3�^z3�ir3H�3��3��3I��3Q΄3wX�3���2'@:3��3��w3H��3~-�3\��3aO3R�&3�q3Om3�I33�k�3l~�3׿�3���2�U�3�P�3��3�'?3��a4�ڀ3ۯ]3�ٟ3"��3,N3wB�3� �3�n?3�?�3��4���3 �3��'3�3m�g3���3�؃3�9�3��3��73[�3Kԛ3�j3�A3{�4���3O��3�͈3��$3�23�w�3�W�3��s3H-j3��3¬�3
/�3U3��3�E�3jn3P�3i�s3w�3�Z3Á�3�^�3���3�J&3��*4s�x34��3��Y3){M3r@/3�L�3�4�3��!3s3S��3��3~��3�	23|��3�c4���2yHk3npM3`��3��3��3Y�t3�d�3[�i3^�p4}�3�3�]�3�QY3й3Z՞3m�4�e�3o9s3��
4��3}R�3
n3�J�3y 3̦"3�z3^�U3���3���3�k�3���3���3�UV3�74X8n3��Q3�zS3f>3�3�v�34��3=�U3P-�3��	4,�3CD(3�ǋ3`��3�6�3�x83���3q�3d�3��Y3�W�3P�3ɋ3�ql3a�(4c��3<�O3=�3���3�vr3F�3aT3	�33߶�3b�3��3o��3�J3�6`3!�$4çb3o�3���3�c�3�u3��4�:�3��3�T"3�74�a3�73@��3Fyl3�9�3h�=3��3PF3�~4�0�3���3�#�3(͓3�[�3��3RA3N�3ϲ;3���3��t3y�4���31�3�|t3N�4|�O3x;�3�2�3��4��3D�3��3|�|3i��3n��3W�3���3X��3��3jg3�v�3��3�ݴ3��`3Gu31V�3[�3��O3R��3��4��!3\�3,R�3��3�>�3���3�ѐ3��3!h�3��4��64`�3g!3�G3�7�3z�3�^�3|�C3�˾3���3('�32��3x43p�3|u�3:c3DĆ3���3A�3P33���2���3O3[ו3��4K&4vf3C�3e6�3��3���3�W�3E=J3��3�II3 U�3u��3/ˋ3��o3r�M4A�3V��3z73�Vl3�
�3��31i�3I$3�3=�34l^�3�`3X�<3��3�Ĕ3��43�
(3��l3+��3��P3z%�3+[g3><>3�>3N��3�8�3�23��3Rs3ZLP3C/�3���3�O�3��3eS4�4��3�� 38�d3ٔ3V�a3���3��e3�Զ3�j
3�@�3��_3��4��	4�:4�M�3 ^3�3��3�2`3�E�3a��3��X3T��3��#4	$�3��33��3}R�3x7�3��P3�8�3{p�3���3qZh3�1�3��3���3�{�3p�\4#HI3��3��,3�vk3�K23_�R3���3�:�3[ڦ3���3c7�3� t3��a3B0~33GBO3��3i163�Z�335�3��4}��34�3oI�3Z�+4�U3D�3�:�3od33��N3'z�3w�3Z h3'��34��3 <�3[�3P�63>��3HH�3�Q34:�3�XW3PU�3�E�3�4�-�3�+�3��23gc(4�?k3�`3;h-4~E�3�ݒ3Z.�3��3	�3 �3�4/��3�g3�rk3��q32��3豕3c�3��83 ��3*��3�<�3�W�3ڭl3q+h3�\�3��z3��4�iS3�#3>{�3�IV3�o3�;;3���3�K�34{/4��3J� 3��3.�I3_�3���3Y�3�g�3�?3:�3�&�3�y3�}K34��3�:3��&3Qm3���3ݩ33y�3Z�{3��3�j3���36_�3yMi3:39036h3M{�2�@93r�3�Қ3Y��25�3B�3�_3nX3�
�3���3h�3#��3;�Q3��r3��\3�d�3D�3�/�3a�3�E�3`��3�]3��3�,�31��3���3/03�Ϝ3<�F3L�3i+�3u��3��M3��3�53٫�3�O73��3*3Ls�3���3�;�2q=3*	4Ѱ�3_�j349�2�C�3���3k�2H��3)"Y3XW�3��3��3$w~3��532�3���3�E3�e�3�t�3��3��93�b3d�533�[3c��3�*�3��3I��3ݎ531$j3.��3
%13%e3�3�3�3�i3n̝3S�(3PȒ3>3u�4�Wv3�E�3���2h{�3�J;3�؏3lm3Z3��R3*24�|�3=P3��G3��3�Y(3E 73� �3y�	3T`�3t�3A+�3v:3Bsn3���3���3^�b3�RD3��u3��3�S�3뎪3�h�3��53�3fM�3p��3�M3`23��3��83�I3���3D`'3Zy3
&/3��3� )3z3T3�L3 ��3���3��b3L63�Fr3?��3ϣI3��3�.n3ZQ�3q�34��3X��3Z�&3+Ef3�$�3�fF3���3X�23�pi3'/H3�3?��3�3p�I3 �4%�63��3���3ZC=3��'3��3��m3�"%3��f3=�3a�3�S23�n3��3��]3b�a3d`�3��R3j7�3E'K3Z��3H�3�os3�}3�04�23l:?3�N)37�3��3YpI3-K�3�D3�xK3Ь3��3���3�73CQ3!)�3iR3^E�3�+3'��3?1�2�p�3��n3�hX3�),3] 4��2DЇ3O3�/3_~3GB3�T�3U[�2��#3c��3�2�3�k�3�3�3�)3;�)3U��3�^�2T�,3�l3�.�37~3+�~3�AT3`�3V�J3�Ȅ3T�13�L�3�3�Ut3��3�n3ג3�v�3�V�3���3�Bn3�4"��3�g3��n3�}3l�3"u,3���3�˙3V�3��3�I4%Z3F�t3��3���35R3�I�3�V�3�}G3a��3�m�3�j�3E�C3k�J3x\�3H�[3�3��3�43��3W�33���3��3�V3�B.3�44��P3�\3;�_3V��3�*�2rq�3{>}3��I3G�W3�i�3�@3T03�@3��|3��p3�$3�"�38[3��w3n�3��3�J3�a�3�P	3�04��3�s;3�|�3FdH3ٙ33�V3�Hp3��3��w3D��3���3�]3uK�2��e3yMt3�r�2�5N3�k3�M�3��%3Un�3a�;3�E39�u3��
4��3�bB3��13�m3GX3�R;3:83h©2��3.l3��w3�Y�2�h`3�D43.@k3�M�21U3#�3�M�3_o23PJ�3��3��>3�VI3�h�3�y~3��w3��U3�ud34,&3g�^3�z3S�$3�R35ZZ3��3�^3CI3ݱ3��3��@3���3+�3/�3� 3���3yA3!�3�3R3149��3�2g3��3�U�3�� 4��T3%E�3�� 3^&�3S��33��3T�d36T3�{�3a.U3�z�3�n�39�b36̺34��3���3�A23*33��03�54k3��{3�nP3��3�|D3R�M3n��3�\3�3�3 �3j��3���2 �3�[�35T13Ü�3��3�Ġ3�03f�3�ܚ3�`3梁3�i�3��~3lH3<|3;�M3�93�3��3�J%3Ş�3�3�#�3x;3D��2%�3ò13��3~��3�,3�]3�x33��3Lr�2�l3��?4<`�2[X3��3(��2(S�3{a#3E�3��J3'?�3 5�3�3��3b��2�h�3�7�3��3��.3��2�
�3[�-3��3,��3��3��	3��c3��53=3��3��3��233U23+s�2���2^\�3�>�3�	Y3�31s�37�3��3�p�2��c3��3�f;3�U3��o3�vp3�t3��k3�3]�3��O3�3��93Q;b3���3 4�2/�3�xq3�th3��2��2R5 3��3z�V3�[.3O3h)$3O�e3��.3�=u3��3,]3�g�3C�3�}3��F3=�b3�43��43#3� �3ߛ93�3E�73�3M�2�O�3tI�2֖�2s�3�2�z3��3jl;3̂3$q�2���3�j4}�3�E�3�$f3?{ 3�s�3h�3�gB3;83	z'3JG�3�֡3�&3�j�2�EH3-�3�B!3�f3��3�o<3��2��)3=��2��2�3���3��3�O�2�m13�"3f�3Z)93��E3_G3&#�2��>3{�3�u3�t�2��K3 )�3�s!3w0�2��i3�-V3�g3q	�3H��2��29A,3��3�a3�l3��R3��43�g3�}53L�3�r3��G3�4��p3��*3p"�2m�u3��
3� 3>�3�%�2�G�3���2}�3�=3� 3���2\-�3�\�2��3�e3��*3�I3��?3��43��3�^3_��3O#�3��33���2�[63�73���2{+�3e=�2��-3��3&�I3<�3�L!3��)3V�3H�3���2�43�x�2s03h;�38�S3���2@�u3��I3�<73#.3�7�2��>3c��2H��2��3�%23"j3pk�2��3�GK3j�3�$3a!<4x�3d:J3Jk 3QA3v�2�)3��3�=�2�O3���3��E3�n�2�o�2��	3���3p83�hV3aq�2��3T��2+�3sV3T')36�2���3�P3AP32�3��63lC3Lm33�F3i�3�T3�aE3�5�3� 3<��2��#3M�L3�:�2]�3<iG3��L3�v
3��_36�/3���3Zh3T �3@��3HI�3w'�3a��3dy3s�}3�Ս3�R3�D3�4�F�3U�3��r3e
�3\��3c@p3�<?3^��3JTP3��p3��3d�3�k3�,3K|(4�*�3��K3���3	\�3��@3�<y3,�3.�c3Ú�3�U3�d�3��4�3��K3�>�3s�p3���3��W37��3�C73���3�f�3ᓞ3��;3�#�3��[3�e�3�O�3ᐈ30�W3Z�d3qh�3�'3�v>32�3O�4�#�3?03d��3�z�3��E3�ճ3l�=3���3�D3��3��3C�3�q�3�44�Ȝ3��3�P3�3B�O3��3���3s\23�Q�3~?4��3?��32l73`��3���3O03 sN3��3W��3��C3�a�3O-�3>�v3�'3�E�3�j3��~3�|&3X�3�T3FN�3�=V3@pD3��3��4.��3*�3��22��3�A�3hj'3Ci�3̓@3��3�}�2k��3�ae3*4�3H,w3�
4�{3�H*3C��3�G�3~N3 ��34ܖ3B�u3}S[3���3�@�3xJ43ÿ43AG�37,�3�I!3�Sl3i�3�g3��2�m�3_�s3�7�3�3��4a�,3�-y3�*J3E�S3��3]�i3}��3�oa3�� 4�r�3���3D%'3{�&3W�3��3[/C3���3�/X3E?�3>h3GU4ܠ�3��
3��83�:4�3e3�/�3���3zч3�)3-��3t_�3���2��93j��3}P�3�4�3�$3縒3[�T3�NK3*��3ݸ�2�Ӑ3��3+�3؄�3*�_3H N3I��3�׉3�e�3`��3є3S�V3'S3c�3�v3�qt3}��3�z3�g�32Ȣ3 ��3�E3�0�3��3F�)3�+�3��.3���3!\g3U+�3���2i04
��2
G�30�U3�a[3�"R3Y�R3£�3�83YZ�3�w3Vc�3�3�%43�S�3JH�33�J�3��?3H5|3�<\3"�3�Ё3з�30+�3��4Ga3�M�3�ne3h�3��Q3.��3y��3X:�3J�3��3 �3Ā3P�%3�b4��3�`I3h)r3��3w�3�m�3r��3�a�3y��3�1�39�
4�Z|3\��3d�s3�ݫ3!�O3���3 ��3�'�3�޳3ee�3���3͂�3�3fɥ3�i�3�Q�3��3��}3F�3\6�3cu4"�T3�C�3��3��)4���3a�A3�`3aK�3z�K3`�3&}�3�}53��3���3fn�3K�3a,13�W�3C��3�E�3���3Jb�3C��3�UM3���3���3>�3m��3�v4�>�3Lu3A3�N�3��:3�$�3�W�3��L3�&�3�L�3-��3w˃3�C3��3�$g3���3�|3M�3k��3��r3(}�3�ڎ3���3�;_3���3���3I̮3Q�3�ۆ3�Q^3n��3��3��3fE�3D��3�3X�p3Ș*3��3#�3��Q3�3�3��3,03��37?3{<�3��3�y4��M3|؎3�@3Q�3r�X3Z�3�X�3=�3aǙ3��3���3��w3��]3�a�3S�3f"y3���3�>3�'�3/��3��3Deo3���3���3��(4�U�3�Z3�ML3ls3@ߝ3@"�3��3}��3!{3�t4�3׋+3�-�2���3�2|3~�3�,�3u�3�y�3I~g3Y-�3�k3i"�3�D�3��4��e3�S�3���3Ѣ�3(F3��3�X�3�!31��3��3<@�3�[�3/�2}u�3��3�r�3��3+|3�L3|�A3�K4eO�3�C�3}Z�3S!4�ō3%l�3}��3��3%�f3b7�3�3C`Z3��3xӝ3���3_3�3Zj�3���3��3^��3�Ϊ3BRy3���3��}3�~�3��]3Rp3���3Bc�3��3#��3� �3G�l3I\�3͒3�vp3�;l3B2�3�	4�D�3�Ї3,�2|�P3&_�3؈�3ěk3k�c3�&�3��3;��3�A�3
{�3sr�2��3�-3�~^3��93<��3�63��i3���3�z�3��A3=�(4��3'�/3��3x1x3;�53���2��u3�uP3���3�&�2_#�3�D^3�"�3���3��3�^3^yd3ۦ43��3,3�3}��3�y�3C=$3c�30�3�7�3?y3��3i+F3�6�3��3�G3;;}3�<D3�}�2騜3e+3>d�3݋3@p�3J03�ӈ3pU�3�T�3�b�2�*3�593�D3�Z3$��3e^�3�XP3���2��*3n�.3[�M3�B�3z�93Z�3:3Eʞ3oH34p�3644��2ON3&�3C�3��3]U%3���3l�e3]Z3&�3�PI3'�'3=�13P��3�=3�-X3��3kDQ3v�3��3�_3@�3�3y�3�"4B�:3�83��36��2�")3;�j3��E3�3Q��30��3�<�3c�v3���28[�3��V3��3[��3T�3�QU3�Nj3n�3�E3$i�2O#^3��3��(3�.�2u�3�ތ3�h3E�H3�HE3Uj$3�D3��3K�3�g73#��2�d�3�z3y�j3��{3�(3֪~3YQ3�}�3彩3�"3�� 3�@-4?g3��k3c?G3)�3[13��^39��3�AS3@��3,��3��3�3���2#@3B�33�3��313M<�3��3���3�3xGB3���2�X�3��H3(	3ι03��3P�#3�Z�3��3:�Q3�Ʌ3*��3�z�3:�:3�"3kZ�3U�I3H�"3��3t+%3d'�3�"3(��3L,3K33��3x�3�+t3�g3�_*3Bb43X�3Ol)3�*�3=�+3l}�3��#46�3��s3�=93��f3;��3�mb3(X�3S�F3T)u3�E3���33�V3<�@3
�[3���3գ3�g3���3sv3�Yy3�s3�(T3��2?ü3]�4�3p��3�#3���3�63K�.3��3B3_,�3A�3�4Tf3R��3��2�c3
G[3��/3mfp3��3�k-3���2�3)z�2��3Q�|3�f�3R�V3V�3�uw3�=3�U�2 �T3ry3��V3L�3��3CL�3�x3��k3Xk�3��3�x�3��h3��3)�~3���3t�`3�ZX3G}B3H��3�h�3)A`3���2vI%3ӑ\3�H3lA&3<*3�	�3�Q+3M�?3�33�j�3ُ�2Yψ3���2�K3�qz30�l3��13h�3��3!Z%3��"3��3�xg3�33�,�2wS�3AaM3Ӈ�2(
�37,34��3d3� n3Ʉ3�n�3��23Qx3�C<3��\3Z2C3��A3�'�2��M3��v37Y*3��3N��31�3�E3n�3��03�a3�.3�g3��33wy=35(33o�3Z&3��k3��X3`�3��33/QU3-��3��3l�?3ΞT3x�h3���2 ʂ3�0�3��3qx3n�30w3��3��!3��3�53{|30�3�Xz35,Q3�D3���2���3�l&3�+3�`e3V�38�3e�)3	lR38�2��n3q6�3��3Si�3���2�d3��33eA3V�i3���3���2E�~3ǧZ3D3�3�,3R�35N3[�,3G63��e3<3Zu3Qu3�V�2��3h��3Fq�3���2S��2��#3��83��3�	�3�@�2,yY3u3�a�3�%Z3�Ҕ3G�13���3I�>3?#a3��G3U' 3�3�3��3E�2�&3�NY3�JP3�;�3��Y3�\�3�mw3�O3Z�3l�
3�[3�2�2Ŝ3AZ3F4G3-H3_��3^�l3�3�MM3;��2ЧX3��V3�;�3��2�0z3���3�3�39��3�430�L3�Ҟ3sG3��#3��3���3}�28/O3�~3�%3|��2ʕ�3�d"3SN3i�B3ү3�E73[g93��R35K3��3�"�3牸3쏆3҅�2��3��e3_��2;�Y3��03ԕ33�31�3�\/33}D3M3��3a�`3i 3p�N3BG3z�~3�Î3>�o3��3b3{��3��3�|�3,�,3 �/3�~b3a`:3V3��i3%`G3M�3�<�3��U3Ç�3D�3If�3+۞3�5Q3C�y3 �3�%�2*;y3á3�,3�S@3G�v3!Y�3FGa3G3�R[3�<3���3k�-3k
f3eх3=�g3�l3�v�3i�S3��	3��3{�3�x�21X�2<
�2s�3���3�p�3��k3�5�3�׍3�hu3�x'3�e?3��3֜^3�P�2��A3�k3ό�3�P3��3a8i3���3�ώ38F�34�334�w3M�93Oz3Y�h3!S�3��k3�RE38?23�i+4�K#3��U3s��2�	�3X�g3�q3�T53�3���3X�e3�2�3cK3M�3��3�Z3�B3�>�3 �,323P�3~UG3c�D3��	32mF3@��3���3�53� �2J�3��3Z]3 �;3P�33��3H3��^3�	A3��b3��2���3�n"3ĭe3��f3�,<3��2o�>3��l3��2M�3�V�3�<�3��@3A2�2���3G?�3�K3��3�B�2�3"*3p�%3TB73�a3S1[3ӆ 4ׄR3�l3H,3j�3@3�63+W03v3�:l3�5�3a�3�[33;�2鿊3|K#3�#
3u>3�3�H�3�%3�G03&o�3hR�3D�2���3�3�z3��3�F^3M43Y�3b��34 �2�s�3f�3�Y�3���3D)�27X3��3��3^�31;'3ꤠ3?�)3�;�3���3�zh3գ3���341"3U�3b�}3~�(3��A3��3��K3)o:3:i�3J��3OY3�H�3i*3y�U3�L3�� 3��3[3�Ĕ3j8&3j��3��3 e3e��2R�4e}H3!�3�^�3׮�3��3�ƪ34dk3���2��3v�z3��3��N3y%�2���3c}.3.E3�f�3��2u�3�C\3-��3���2��37գ3�!4 `3��3w$h3��3��3$��3OR~3g3C�J3(S�3�7�3��3s�*3�ؽ3ă�3Ƈ�3�М3%w�3�M�3�X3꛺3�3�VK3�A3U�4��83�?v3�_F3�'y3d�M3�_�3r��3�ʂ3]��3��3 ��3_�3�[�2eX�32°3ӝ�3��Q3��a3�.�33t��3"6�3��4�_3^�/4,�3�b�3��N3o�[3�,3�ր3�k�3 �3u�3�[�3���3��m3U&3Ȋ3_
|3v�3d��3�ښ32z3|��2n��3i�\3��3|\3|�4�J3��d32t3�M3�3�-3N��3ơW3�H�3O��3F��3�3i3���39��3F�H3b��3� �3S�3�p\3���3 t3]"3gC3�4i]�3^l�3lw�3��3(�q3T-3�T�3h 32ݴ3�"4�Ѹ3�ޠ3{�<3Jw�3#�3*�d3�?�3e$.3i��3+�W3���3T+�3�Nv3�+�3���3�f3��H3LH�3�0�3_�_3ݾ�3]]�3��Q3�yr3��3�"�3eQi3x��3y��3�1�3�,36�3�C(3+�4V.3�-�3�*�3��3m�\3��4��t3���3pF�3�eu3(3�3�v�3>��3v�S3�&�3�(�3���3w�V3�	X3�{�3�@H3�5�3���3r  3� y3��3��3�O�3⫲3�4G3�4�3�^�3�Y3�s3���3}8�36�3��-3i�b3��64R��3*��3�#"3���3/��3��3r�3�J3S��3_0c3���3��Y3�3ݽ�3���3/�M3:%�3W7�3HPR3���3��3퍸3@<A3�+�3�$	4uu�3�G�3]a�3��3J�3��d3��3~.*3�!�3R6�3-�34~T3�4�3��3��
4��`3��3�Wx3V�,3p�3�{3���3@H�3���3D]�3L��3T��3l�53z��3��3�>3���3A3y�3,�32��3�x�3�,�3��3�޽333*3�3?3{�l3jc3�#3���3p�j3K2X3�S
3���3H��3蔚3ēU3�»3�D3�k 3�Lq3��r3'|�3��3?��3=�%3�|3op�3�D�39A3��3��e3rg3}3��|3xƉ3�=�2��
3��3�Dy3Nʌ3E&�2oA�3���3H`03y@3��k3��
3v�2�R�3�O/3 �"3��3i֚3�3CV3�f`3���3� i3�he3DT�3��3*�P3U!�3�Z�3�:3E��2ی3��M3E�3�3�<3��]3��3�H�3�&�2W^K3Y��3��B4<	�3���2\`,3|��3$�m3��t3���3�4?3��3��3s3n
C3B�!3�3L�u3�p3X�3Z;\3c��38K�3v��3�K3�PI3�'3_k�3�|�3.�3W53sZ43��N3wED3<ǘ3��"3|mv3G�3}|�3�g}3��L3���3v�F3 c|3Q��3~�.3e4m�k3�n�3̒p3mU83@�$3�4*gE3'�v3p�3���3��c3���3��3ڗ3N��3N��39��3��@3�>3o�p3L��3�ʐ31?3�3i��3&�b3�ܵ3���3g~3��d3(
�3���3F#Y3��3g"23���3��3�w�3�E�3�o�3��3�,�3'pL3�a3q߼3s^3��G3�%�3�3��3F�03�g�3���3�fJ3&^o33�4�T83I?h3ԕ3+�-3c.D3�EX3Wi3ë93���3G�3H��3cn�3��3�۔3i�h3�vz3�گ3�]3�\�3��!3d�s3%�x3d�e3D�3��,4���3帖3�s3ʪ"3\�2��3���3Q�3\��3���3z
�3�oF3��.3�X3�$w3�+�3;��3 �3�Dd3x�K3�Z�3�oo3�\3�e?3�&�3PF�3��3Ϻ�3�!�3 �<3�M\3)%�3�S3V*u3Nާ3��3�[�3��t3_�^3�^�3;`3�B3�3���3��@3lR�3�ik3��3"��3O	�39(3�^/3e3Z3i~�3G��3�Ay3��S3r3�Ի3��[3e��3=E)3y��3L�3G�3�@3
t3�~L3�>3}k�3�0�3�G3��q3���3q�J3a�z3��s3��g3��33qj3�h3kH)3+�M3Ԕ�3VB�3G؄3�3���3�f3���2���3Һ3l��3ԍ3ҳ�3)��3ݡ�3 �!3�׽3�W3�rb3$yE3r�3�93�u�3h�"3B8^3�|O3��4�C3�h�3Q��2�AU3!j[3��3�n3��3��3��'3V�3}|n3C�^3b</3�;�3A)n3�863��E3��3��3!WN3va�3H�"3��!3�w�3pF}3�[3j�[3�3�i�3�ܳ2f�3���3��[3�:3宁3�E(3�343С�3P?3�&J3�#3;�39q3�M�3���3,�3��I3�j�3�x�3H��3�e43���3kb3}V�2cjj3�3HU�3Q�3�g�3	�#3���3�jN34��3o�`3��&3G%�3�=3(�\3�Ѻ3v-�20��3Q'�3_�3�IG3�3��m3�"�3/o3)?3�B3H��3q�M3^ݘ3ii:3o��3K3Z3!�4�H3b�3G,Y3�X3l .3d�&3G�h3U��2sE�3X��3�4�3HCk3+�2�;3ڌ�34B3�
-3�2�F]3Ӌ_3Jv�3�h�3]�?3 �y3s�3e)P3�<�3�D`3�\3�$<3�$3.W3��M3�o�3�* 4$:�3��Y3�/)3u34^3Q(�3o|�3$��2�k3(--3� K3�`3��43��&3��<4Էw3h��3j`3��D3"3l3ہV3��!3 
�3�9�3T`�3|W�3�2�R�2$��3@/3�3�"!3QF\3ȷA3y�3MM>3O�=3.<&3��3�i3�S23� u3q�h3qtF393:V�3@.�2R%�3c*�3�1�37,Q3�S3��3�M3�0k3��3v3��3'#�3��]3��3���3��32��3O�3��O3A�$3�l�3o=;3�3��e3(p3'sQ3��3���3�wx3�g3݂�3l�3,3%�F3W�3�̐3��2�*�3��*3��3�͔3�3T�3iN3q�3�$3�A3��3-2�3Of3�m�3u�3z+�3C�\3t
33�5�3��i3�0�3�ۚ3X�G3 u�3��C36��3}��36�3	�L34h�3��O3��j3�׏3Ԅ3*=/35ߝ3�z3�H3�3�o]3�#'3t�3�ؠ3��}3�A3�ڶ3��)3QCG3�K3�3�393��3� a3���3��\3��x3Wj{3�n3��63��c3�(|3ͼ$36]`3�3�ڽ37td3��/3�ٙ3�aQ3Wr�2��3A<36�3��Q3 �i3m�X3s�73���3�=�3�-83*(3��N3`�3��F3߈3�h�3�yN3rY3��3|M�3�dV3�f(3lr�3T�@36BY3yae3:G3
��3�(3U�3aG31.I3�'*3b��3'�3��t3��36q�3H�|3��U3.z�3�n2B�3& 4*�3
Wg3�}\3pEm3 *?3s�53Eec3l�3�3=t3�ˌ3�TZ35i]3��3n�4W053�#3x^I3�mF3J�?3��-3�y3��#3��3�e�3i��3N|:3Z�&3��3��U3��3s�a3%M�2��3��93���3ͼJ3�E�3�/73�g!4C�Y3�)Q3��y3�2�3�83ꢂ33�s3LD"3�j�3�Ҭ38Mr3��3��2�'�3Pe-31�3���3k�3Q��3d�3ų3�h�3n�N33u8`4{ڍ3H�H3���3!�V3W.33ve3�k/3�3<363� �3��3\��3U�_38�63mL�3;�p3�x�3ы73$��3�b3,aj3pS�2�'3S;3&84�3�{L323R�K3:d3h�m3�s3P&�2� b3<C�3uЫ3��.3[�&3��b33J��2 F=3w�2ʎ�3u��3R�4e�Z3��3\��3�E4ޜ�3	�83��$3���3h��3X�3l��3}'3ej3ƈ�3��3wx�3�A�3>��3�S�3n@,3��3Ԗ�3ݮ3~�r3ũ4$�~3A��3J�l3�A4��3��3��e3�2�3¡?3���3E��3�3��3�W�3˧�3'�u3��63�	4�Z�3C$Y3�5�3��3�c�3��E3��4?r�3Q:4��3\�4�}3�y�3�V�3��4�B�3<D�3	>4�g|3Dc�35d	4��3�~�3:��3�� 4�Eu3�g13&��3�h�3bB"4y��3�4�=�3�n�3~^(3I]�4)G�3t0u3+?	4|��3�@3���35~�3��$3KA4߷4W�3ӕ'4��L3}�3:k�3u�53	y�3g�3���3�G3��#4���3F�4{��3��4O�3Cu�3rڑ3���3˰�3�|'4д3ьu34��3��/4O��3-WT3�U3p�4ZN�3m�v3��3~�n3�&k3�#�3�!4_�l3�Q�3z�3�(Y4�5�3垓3���3�?�3J�3���3��3�A3¢�3	�4|+�3���3<��3�3�4Z��3��4�r�3��4 F�3Ć�3��3�ʧ3P �3y�h4���3=��3���3��3���3���3�#�37$i3"�3��4"�!4�]�3}�3��4��3�?3��3��(3��3�߻3��4dă3�"�3k��3�e�3ȶ�3̔3䜳3�V�3��3)D�3'��3���3�mi3�2�3_�4i��3��b3���3�3}�_3F��3�O3�'�3m�39Z�3i4��3>�|3��A4�w3:��3		�330m3�hx3���3dx�3,";3t��3K!4�4ܜ�3�Ci3�3�:�31d�3V9 4C483ك�3.�/3d�3���3�"�3}��3XD34dJ3�h�38�3I.k3�N�3�^z3&�|3"�3�w4��4`�4���3���3�ޭ329�3E�?3o��3O3<`�3�t|3��3%�32��3�K3֫*4�3[G�3�#�3p��3��3�X�3��{3��63��3.�4y9�3���3��K3�r�3��+37z3\�3_(�3�u�3��338�35Ӑ3X�3��3X��3Sz3��r3u��3�}�3���3B�3I�3���3i��3�}�3[4��3�RW3[>�3�ۨ3ڕ\3Ч�3���3JԳ3��p31S�3��3�F�3qN�3�1f4T��3�4x3���3k��3�M�3<�3�o�3J�]3�	�3)�4��3�<�3��3+�d3��4���3ז3q�3�[�3艁3<64���3�"�3��3��P4�}�3��3=�Q3[C�3D�~3���3���3�AT3*t�3��4���3���3�lH35��3rG3㰅3WA�3|��3��4p҃3V��3�l�3�f�3���3Q'4Am�3%}�3^3n��3fl�3�&�36�3�ֱ3~?�3�R�3X��3�HY3}�3�?�3${|3���3*��3��[3��3֥�3P�4?��33�3\�3g|F4��<3��3��3���3h�53���3J��3�ll3;��3kN4��3'�3P\p3'�3��3!;m3�v�3��3���3�e�3N��3��3x�3�N3�S4�v|3(��3���3�˙3�	�3f$x3M�3))F32e3P��3���3��3<�C3~A�3J��3U��3\nq3".M3c�3��36�4�ژ3�-�3��3�H4�Y3�=�3��3-d�3a��3(��3���3�$C3(I�3N��3O�3�C�3�,f3&v�3���3�n(3�z�3�У3AI�3p�q3�3�yJ3!�3o�W3�+4w�3>V�3�v�3a�I3��3; D3�_�3�ҟ3k��3n��3�1�3�E�3��93i��3"X�33��3��3�@#3< �3��3]�3��^3gKI3�?@3+��3g\X3��53ɿ3Ӿ�3�{3�7l3y.�3�23�6�3�=�3�3O��3�s30=�3���3��-3NL�3�*�2ؑ3�y3��3ͭ�3��3F�3���3ԕ3�633���3��3�L3v�3=P3��]3:��3}��3���3�#�3�w3���3�:�3e1O3��e3�ݤ3PtU3/�A3d4�3�3sc93�C�3؇�3H��3��J3��3$�3l6C3{�w3���3�j3��W3G�3.��3O��3M�d3��l3*�3�d�3b1�3�n%3�Q63
��3���3*��3�*�3k�3_��3:WM3G q32R�3���3�rP3��s3ꮑ3�3��l3rG�3A�3Wi&3��b3�*s3S<3�33�`�3ls;34���2XO�3��p3��V3��H3�)�3��*3e�B3<o�3�i3Tyn3'�34�3F�3Ŀ�3��3��3b�3��2��4I��3"�)38@03��3���3CI�3�x�3�[�3�'�3��3S��3�z�3��}3h}3���3f^3I��3x�3�X3��3�L 4Jh3��R3\3|S�3�;43��K3�@�3�X3G��3��3��3~TZ3J"�3>>\3J�3[��3^4�3z��3\V�3�`3ӗ;3?�3�IP3?m?3 |�3W¿3�ţ3+bw3߾�3:�3pK3q��3X&3�T�3)�i3�5�3a=3��31��2/�4v<3�R�3,l3�3W�X3� s3Q��3oB�3ۍ�3�f�3&C�3l��37H�2x��3Э�3���3U4�3��|3��3�V�3�[�3z�g3�̎3���3mw.4#m�3)=�3J#o3Ie@3m�w3xU�3�3�^33�S�3ʅ4�W�3�h�3��"3E'k3C�V3�rQ3T��3٫73f�3oXC3�y4䭔3���3�%\3�L�3�o�3�B;3���3Ah�3�l63Y�3	n�3�{�2P�3��4�"�3D�y3!�'3�;�31n�3S�:3�r�3a�q3�4Q�63�v�3y[m3��3h'3�|4��j3���3M�3�9S3���2Ђ3��l39��2�)�3�4i*Y3�I�3��	3��a3��3�vh3�A3�g!3���3b�.3w�4�%*3�'�3�`a3bO�33�13�{c3�Q�3�lw3��3���3Wk�3�"3V��3}O4��3���3�j�3;��3��3|��2�q3�>3b?�3y"3~��3��3�U�3�m3_a�3!�83C1Y3��t3V��3�Ղ3�}�3�N"3�Dk3��3�l�3�R�3:Y\3��!36V�3t63:7u3��x3(0]3��3f�3Q��3:�~3S��3�<?3a��3�<m3�3�pu3���3j�3Aӏ3n�3�?3��3f�3�@�3�G3�UD3oX�3�w�3�M�2�3�3n�3R�U3F�3$�Y3�]w31�3�353Is-4lp�3�'3wH3��}3�^Y3�T3DQ�3|k�3��]3�B�3���3aN3q��2�p3���3�|r3_��3ړ�2�1f3�ϝ3mV�3�E[3��3]�3n@�3��$3P��3�CR3^��3��,3M?�3��3X�3+�j3�t3�(�3 "3�i3��p3��H3��23\�3�
&3��|3�Y|3�U�3l�	3���3Yb�3��3�5c3x�3UF{3U�{3�o3ŋ3G*�3Wt
3`/U3���3�y�3��3ǌ�3{`�3ͱ3�"3�͏3�H33�3qQ33`43��W3$�83T�/3���3w�k3�943��,3��3L�B3<�3i�3ʍ+3#w�3��3o]f3^�D3��(3���3%�93v13��3.�3`�3%�_3 �3p�3�or3⡑3PT�3$�
3�K|3�\O3C3[t]3�x3u��3��>3VrU3~/	4B=�3y/�3�*S3��3��3�3Q�'3�3�F{3v�b3�^4�my3D�83QXy3	�*4�Ii3=�,3:�Z3R�3[̂3��3K63][?3��x3Hv�3���3�}3/�$3�݉3�(�3�:3��3Ԩ3t,~3t�>3C;�3`V=37�X3��f3�4	��3&#�3t�3�i�3m�S3Z�S3o̦3r�3_�3ν�3�n�3���3u}�2{I3 �73#�3f��3�2�2�!�3�Ln3&e�3�x�3�)}3���3�3x30�S3��m3��3���2�T�3�AZ32S3��Y3�"�3{xC3_�13q�3�B�3�?3��+3DL�3�,3&�33�p3%;�3:w/3��+3�ZU3���3w	�3#�O3!EX3�ޡ30�P3|VM3�;Q3���2�O3Lb�3(�3FX�3�cm3�Q3�r3��3 93,��3k֥3�;3�v3|3��3���2�^�3��3.�H3=�C3�ӗ3X�3gu\3K�#3�	-3[%=3^{�3Z��3���2=Ƚ2m�3ֽK3sX23k3��3�Xz3�1'3%��3��>3�@3�_v3T��3_�33 3}
Y3�lB3za38h�37mu3'�2�+a3$�3~w�3��H32��2OԠ3�H3 D[3}ē3'YQ3.;O3�g�2U��33�t3D	3�[�3� 3c]C3X�D3[?X3�63:r3�73�	�27R3]�q3VՏ3u�a3��2V�3U+3���2N�j3*�2A��3L�03ֺ�3`�	3��43)A3I�D4�3s�D3e~�3��*3�*�2��U3�ɒ3�v�2��~3�x�3���3&�3���2_w03��Q3�W�2�{h3�3�Ј3�3���3�kk3Zj3�7�2Y�4bg3>I3��3�(83�U3U�3�<�3R,3��$3[x4ڳ<36�3���2�5o3o8#3�Y/3aTT3���2��3oi3�X�3$�F3g�;3��R3e`�3P'23�/3Ր�2~��2�^(3qo\3)��3��-3�g=3`��3�QH3�I#36813|�w3.f3��73e�~3=Y�2̠�3Y�3��&3�:3+3�ir3�:4gb-3�ɉ34T13E�*3_w�3>�~3zyT3�c�23�Q3��3���37�3ܶ�2H��3��3AE3Fk3�
�2턡3�3�3伛3 -3W�2f�2��3�w"3�=3iX3r��253<)3�b3��Z33��3���3��Z3l<`3��2[�35c@3��3sM3FXJ3�YX3E3���3a'[3�̛3�y3"$4���3d �3=��3߮3�,�3���3�'r3;�c3�t3�Y�3�x�3�<4��]3��3���3~�|3R�3�1�3���3��3���3.e�3sӝ3	��3%)�3��W3��3��3�B�3�5�3k4O�3Ʊ�3*�3·�3}p�3='�32iO3�@�3-�3�s�3M��3�xF3���3�34m4+��3�#�3��3P��3�¢3*�3f��39�3��3=x�3A԰3
�43tO3���3���3�#�3�x{3��3�\�3�{%3N�3��3b3	4$t�3�x4�S:3���3$}�3k	M4�+�3�ܭ3FԌ3���3���3φ�3~2�3�sI3A4P��3b)�3�d3�bA3��3scp3�3�Z�3N�3v�3��3��3�N�3Â�3y�23V�3�к3��3oU�3c��3��n3R��3O"4(x�3�3�:�3Zj�3���3��@3�M4�2�3��M3Z �3Mٵ3��3�׊3��4c��3�c|3�-13K#�3�l3���3���3|�3�z�3�<3�3e�G3T�3x4$�3\pX3X�]3�
4�yg3f_C3��3OK3�74i��3���3�I�3h#�3iOA3�.4�n�3��3�J�3�,�3��p3��3�st3R��3U��3�"4ld�3�V�3cM�3R��3���3��3��3ƻv3"h�3��3C\�36��3���3cO�3k�i4�<�3��3�7�3��3p�m3%#4EQ�3=U�3��34��3c��3�æ3>c�3u�38��3��3��=3'D�3��u3�5�3a��3�B�3��3w�-4���3�+�3y��3}Z3�+�3᫒39.�3�^83��E3��4@�3�2�3��>3�W73��34��31�3�:�3Kw�3�O3��4o/�3�u~3�13,�4�%�3���3��3���3X_3/I�3��3���2~��3}Y4u��3�@�3z�23ƴ3�&�3�03	��3]3U��3�8?3Om�3�>3o�u3
J�3�S�3���3Q�3���3\��3�Ab3���3��3 ]�3�:3>	4�;y3�y�3�3���3g��3'k,3|'V3�7w3���3�3�j�3���3S��3���38lL4��D3|w�3���3-��3%C�3�D�3�>�3J�t3[	3;k�3���3�n�3�jq3p�3T��3^��3��3qe�3�y�3��}3��%4/{3��3��x3��405�3�Χ3Y3 ��3��P3WL�3���3��73�\�3��4m��3�r�3�P3���3d z3�*�33�3�Lo3�3�:3a#4�D�3S�3J��3��4^-�3��3z�f3��3��3�3z%�3�g03W��3y
4�6�3~��3�cQ3��3��3�3B3 ��3�q3w�4S��3�4C�3��3n��3�	4GD�3nG�3&'i3r�3%��3a��3�,�3,�s3�d�3<R
4rF�3l_�3n�L3`�3���3���3��3��3堥3�/3&L4�D�3sw�3���3)�4��3�%�36��3�ُ3��3��3樬3�[H3�g�3&�4g	4�4�3��v3J��3�sv3�c�3ZĈ3{$3�a�3zx�3Ԫ�3v�`3�1�3*NE3rm4v�-3��3��3!Ҋ3z'3��3���3���3���3�-�3�)�3��3�Ё3��3h��3��3;ǜ3ƅ�3�n�3��2G4;4�3+@^3�3�4���3�K�3�^�3Vt3p_�3��3��3��43�t�3��3"b4\\�3��+3;*4ӈ3/�73�4�i3�8�3Q�2304 �4MZ�3|V�3�;4ޔS3�	�3#��3�J|3Y�`3���32H�3�z3�<�3���3��3���3*�3��3U�3w�3.�3m��3"��3�ɺ3|/�3s:�3�w�3��s3�3�3�p�3��3� �3�G�3�n>3�w�3���3�?3s)�3M�3�m4�?�3�d=34�S�3���3���3��3 �3"o3ed�3r��3�C3��13���3�.3+'3ؑ=3133�,�2��]3��]3ޤ@3H�J3k��39�,3ل�2�G83�3:��2���2�&3�� 3�Ȃ3!�2ө�3/�3&�p3VID30�3�Fl3vo:31�%3�!�2��+3�3�33��2�T3�4�3�b3UQJ3�e 3{�3�N3n�3!!j3��%3n-:3/	(3���3-�3�m83�TG3G��3��53�43�!3��&3���2:t3���3��u3�C�3X�3�=3��836I�2 �q3�q(3_3�U3�[D3�=3��23(�X3��N3v�N3��22z�3mi�2'3$�<3�fb3��53~3�!�3�=�2�=3�{Z3,M3��M3 ��2�AT3Y�33ߥ[3�y3}`3�3Q3��o3�QE3�^>3J�e3��g3�!+3�3��2��3��,3��t3n$3/=N3e��3ey3��2�3i�33�G3��)3Ì3��2��93`�k3�43�83:�+3kK73""�3\n�2,D	3Q}Q3E�&3��3��!3
&�3�8�2�:3T�3�QW3�Q 3M�P3��;3��J3{��2|q<3K�3{�3���2|H^3�3�1�2�T�2w�32-3��c3�B3�K3P��2���3RtJ3�3�@3��n3	393v��2H�2
�3�2[%3�G3��2(�2�53_o]3�/3jA�2]�/3v�3O
�2W63�"�2�je3"�3xaP3{xX3�ɼ2t�3ad3T�y3�T3���2��V3b�!3���2Y�D3\�2��c3�3�y;3*3r	3.�*3L��3ڧ3k13�I3ؕP3x�;3�@3�Z3��2)�?3}h3�iD3t+93��2*Y3L�2!&W3���2�X=3�q3Z�'3|�3d(�2Z��2cL�2�̖3>43 t.3C293}�-3�.>3N�,3��'3|G�2
3��+3}_�39;434�%3n<-3��3��3T�z3�8�2�E3�J�2�x3I�3�ը3XoP3e�3�s�3� /3��3��e3���2F8f3��m3M!3��3�9�3��[33Б3S93�,�3��03�?3�*3
��3�D3Z��2�Ǐ3�l�3W�3�S�3��4�jz3P3�ҟ3r�3M�T3��3�g�3�C13��M3���3>Y�3���3�3d��3^A36az3�Q3[Q3'�3=�T3��3fV83H�/3��O3��;4U�3X��3w�V3 R3O|3�;3��,3�93Q�E3T 4~�3��C3�1�2�132Zq3��3eU�3�;�2{uS3$`�2�?�3��G3�u_3&�83���37uQ3���3��S3�Ʒ3z��3�٘31�3��a3۞�3p��3
�3���2�:�2x)�36�3��d3�^�3G3��D30}23؜36V3J�R33H3`��3T�$3`H3��3#�3��M3Ic�3e�|3�F%3��p3dq�3j�h3ۤ�3G5D3d�}37m3��63Qq�3i�_3֒�3�H3xӆ3�[Q3���3Pb3*e�3�,	3[L�3�3>�3q[3���3T3S63�|3:��3f��3Fـ3��T3��3��?3֫(3��r3,�3U�3�8;3+?�3O�03��3o��2�ɥ3��'3��03Ok3��V3o�_34A3jY�3��3�b�3���3��^3��:3ϧS3k¤3d�3�v�2E23��3���3�03Cz�3�o3n�3�w3-o�3��O3�L3'�`3JG43R�R39V(3u�3A)3`e�3��44O�3�6�3�S.3Dk�36)�3�\3��3�H3�T�3g33^��3�k{3m�3oQ#3s04i�T3	HM3��3e�=3$�J3ڶ�3�y�3�<3�]�3`��3�[�3���3�|#3+p.3�w�3{�]3]ۥ3��^3}Y�3��$3|��3��3v��2o�3�A4��	3gpR3̍X3g�-3�G3�U3�o�3Be�3 /�3��3mԒ3+�W3�/�2@Ÿ3�sX3�F3�83�E39͛3Ik53���3��~3ɟ�3m��3�.�3�}03��b3F($3}5h3�F'3H!l3�JE3c\�2��&3�u�3Z��37]�3��73�f3�O3�83>�:3܁3�1x3��/3j��3��c3%i3^�\3l�3��3��93�\93l03ϡ�2xZ|3�7P3��2��I34��3�3BC�3��
3V�3�Am3��Y3|N3FP3Oqc3���2�~�3�P>3�/�36o-3�~4jnQ3���3B]�3��I3]~3U �3�J�3�g3cA�3/�3�Az3	F343T{�3��g3f�3y�\3��H3�R�3B�3 �~3��3z��3�3�5�3���3�83:U\3��3*3�-�3��-3��3`�3ak
4� �3ޞ`3�F�2@�3'��3�>g3��3>�73X�3ܕ]3-3+V3ڵH3F��3��(4Y 3��u3x|V3�"Z3��B3�Z3�l3�3�iD3/��3���3!�*33�>3��3��#3�\"3IV�3�B3�E�3�{J3D��3�3��c3y�N3���3�Hy3�X#3S2�3���3G3b�~3�٫3�s3Sǁ3O�3�%v3��3ͤ-3m��3�"�3��^3f�3�3�Ş3��,3��3�3(343�3-s�3D N3<�3[b3+�2(3(�3[�n3�y3��s3A�4�ߡ3u�S3�r3���3��73�TL3�A3�3Oׇ3�M3��3	f,3��s3CeK3s�.4��n3�
d3|�X3z�r36w@3eB3"ʋ3$532�3֙3G@�3␄3u��2V�G3#o3Д3��3��13&ea3�� 3L3�3��'3)�A3<h3Ο�3��W3�GS3�Ԏ3��`3��3��3���3ux33�h23؞�3E�H3c�a3�E/3o�3�X�3�X3��3%3�݂3�3�ւ38 Y3@PV3���2�ѽ33��W3��3�#3��$3yҔ3�4�3��2Q6q3���3 �o3�H�3y3��3 �P3�f3�ׂ3O��2RN�3��53Q��3��93hg�3���3��3�?r31cJ3N�33YB3��N3�'Z3So{3�"�3��3[��3�Մ3t-�3O:3�_�3f��3Y�,3�z(3Y�%3B�3mf 3�c�3��38&�3g\v3;�3���3;�3m�3��3i/U3�@3��3Օ�3V]D3��b3l��3��L3�@3;K3���3ցT3�3F��2��3Y�P3tn�3c��3���3�P;3���3nM�3��+3�$�3>Q�3�qf3��3�Z�3e#3wa�3��3g��3�:	3��3�_j3���3�v�2���3�<63LI�3�ǃ3�Ԓ3� /3�sh3��3�i�3��3p�q3���3�Ӫ3D\W3��3�q�3mr33�>?3�<�3<��3��d3�
#3���3��3��Y3�l35
b3��{3�<&3���3�Io3�{63"��2��4�bn3q˄3z2w3��3᳂3�Ɠ3-Æ3�3]Ɯ3�]�3Ũ3`#3W��2��3�	�3�{34Q�3��&3G�731�!3$R�3_�3(�3䲀3�4��3��t3�iW3�\�3�"�3�y�3�2A3��2\�L3U6�3$v�3�R�3�'3�T�3qv�3�w30V3�hL3Ax3��B3q�3=�c3�^3.3�'14u�
3�83��x3�y&3�<�377�3�i|3��3��=3g�4N��3��p3:y(3'��3!35� 3��3��g3o�3�gP3om�3�A3wb3U5�3n�4H�L3,�3%��3K5�3fƉ3L��3�3�[3�O�35/4�'�3ı�3l83ۋ�3�E�3N�23�޷3�w�3���33��3�d4Qo�3��x3t�m3PB4`�33f��3�Ϛ3utF31b|3�V�3_�3H�q3�%<3� �3�P3�6i3q�>3vTo3Ш�3#8�3�y@3/*I3���3z*3��3�1�3K�*3�]k3�J�3m�D3���39�'3qcZ3 �<3���3���3t�2��U3nγ3(��3A�13�@3�g�3kXf3	/C3��3k�e3ꃙ3T�3x�3�3�c�3�,f3T2�3?A3
Z�3:c3A�'3�>/3���3�l�3�;3Z��3�{�3@]�3�UL3YB3R�h3�CA3e�3|�T3/3U�3�934f�3��Z3�a3N|Z3Qm4ԭ�3�]>3���3'��3�N�3!'�33��%3(��3n��3��34�3��*3t�3:LX3��3�ߦ3�3zw�3��?3>�3��3���3�sA3j&�3D�3�<@35Y�3��D3�d3|[3]y�3d!3vP�3gR4]a�3��3�J�2G\�3+�3G�3	��3_M73's�3ز3t�3�'3N�h3+s�2���3�.e3*K3��3�@�32�3�`<3��3��3��3���3�~�3h��3M#3��3xU,3ko�2��f3�hH3d��3�x3?�3	�b3zZw3�43���3c��2�<I3�D3 OC3p�N3�J;37tf3�p3B8�3���3=��3�TO3���2��j3�w3-��20=X3�3��3̈A3K&�3ф03�Z
3;$d3O	�3�?t3�>m3d2B3.��3Ѓ3-3�Q�3��&3Լ/3��4q��3�!n3�(�2m�{3�{b3�&3�}43��3D��3/�3:�3�Z3�L�34�2�54mم3fv3-�3��}3,%�3iT�3��3
�3�V�3�Ӵ3�+�3��3/3h4�3�M/3C&31�M3�j�2!m�3�α3A��3Ž�37�h3!&�3�m4�e3d�!3 �F3\O3�b3�r3ǹ�3C|3͝�3�E�3�\�3��L3�P&3��H3�}`3�U3	��3`q!3ą�3z�3wĵ3�n3�B83^�n3��4!S3Ҙ[3y�!3�$93��`3*�03���3P]3*�x30@�3�W�3F�!3l�	3��l3d�X3�3OɊ39��2՛�3�3�1�3��43���2�^*3�3	^3erp3S�36(*3Ki3ƹE3��3�k?3Q�3��%4���3�z�3E"�2���3{�{3�U63n�43�3�A3�vL3Q��3��23z�4���3��4{��3�~�3�A�3
ě3��3੪3���3��3�B�3��84N��3G4���37�3n��3���3InQ3�ì3���3���3��3*�3.�3X�364B��3�4��3�34$��3�3i3)��38��3���3'D
4�.�3j��3�/�3��3ۨ�32��3�ͣ3�;o3rȨ3i;�3���3��3�^�3F:<3V��3v�3z3��3��3.�y3\�4��3�F3Wޗ3[4�@4x��3�Б3x2�3g��3Y=3�.�3o�3)�/4�r�3m@�3�k�3��3l�3k4��3U �3��	4���3���3�t4�R4�;\3�*�3��44� �3L�3N�)3�}�3�Uw3D��3Î�3���3x/�3>`�3m6�3'
4\E�3BQ�3�r4��3�N_3O��3�3�y�3��3� �3'}3�u�3��q4b�4)i�3S�3��3{��3lH�3���3���3��3v,a3��/4T�3��i3͞�3�54m�S3#��3�-�3g��3L+�3��3�>�3j�N3{S�3N��3ݮ*4|��3�bp3��
4��3dd�3���3�`3��3���3H�^3B��3��3�.�3�4�[�3��3m,�3��34��3��3��M3YXx3��3��3���36��3���3>\3�(�3p)#4i*-3�ؙ3;��3\�3��3i4SF�3g�K4.ʘ3�!�3�=�35�x33a3���3e/�3��k3D�3�t?4cu�34);3���3��3M`3���3�YS3 ۦ3m�3g�U4�v�3�[�3w��3pd4�a�3�U�3���3�l�3��3�*�3���3�n�3j�4��&4��3/%�3D�3���3a\
4<�3[�3ak�3I��3�g3�4�4�3�&�3sSf3-��4P/�3��3�!4jj3���3Y�43�\�3�}|3J�-4l-4�(4R��30G3�A�3u��3�m�3���3N�]3IU4�n3�"4LF�3��$3�v#3�X3zM"3:3֞-3C3�^3�B�2/�3�/3Cb3Vbb3�g3N�3+��2_�V3
�3��2��3/�2�39s3��C3�/3t�3;3x�r3�3��3u�2,�	3��3��3�)3$��2=6�2ya�3�P3K�g3)��2�H3mm43�M�2��3��2�I3�-3ʲk3�e!3OE3]�3>��3�l�2�D,3q�]3�5[3��2_�3H7W3ru�2 �D3���3�q%3<�3�h�2*3�_3�m�2�F39N�2��[3��3�T3޲3&n#3Y�2�V3�83�	3g�,3�7�2	m�2}n�2�3�y�2l�L3�x�3�*3�K3*�2���3�'3��3�V_3�3Vq�3O�3UW3�q�27n3�2�2��n3���2��'3WUr3K��2���2d�3��_3�)�2?3]�3;A3�c3��2;�,3̘3��2���2a��2�I3�2�2[3m3��2�T3f%�2���3k2L3ԏ.3�3s��2��2CpU3H��3?�26O3��3k�3�p�3���2T��3��2�D�2�%+3R��2#$)3�3��_3�w3U�2M��2T��3�X3�M03I7�273M�3h�3*g!3�X�2�nU3�\�3[_3f31~�2��83��'3;;�2ȳ2s��2�i3��2@&3��<3|�/3@�2:��37�%3�;	3φ3�:3�<�2^_G3��W3���2z�L3g�3P�2M�$3)�2�ґ31�43Y��21�^3k��2t3��2�>�33�-3�
�2���2��3:3x	3u�93@�3�H�2F=3b33��2��73A�~3ͻ�3��J39�2�3�au3Z��2�a33m��2��m3���2F�3�� 3�3nO3{wx3)��2�3�m3Ę2��2��3�vT3*��2��32&D3O3L�3� 3M��2K�13���2�y3$��2�I53�&3���3U�!3w/3��3��Q3P5-3� 3�ځ3��3�2��3�kK3O�"3�m3���3��32�<3^3h�3S�93��2��"3��v3�*�2�3�y�3�w�3��2K�a3��3էM3(�3��3�D3't�2�R3��3�4:3��H3��{3m�q3D�{3/�3��~3���3i3��3��i3���3Z��2VĚ3M�3د;3�Ab3�h�3��3�F38�3��3�5�2I�3��Y3�{3�O3!��3��i3A�3��D3��3`��2�@
3��]34�D3�r3FN�2��3�}<36?3�3n?�3M 3U�-3�w.3a(x3=�T3!��34Z3T$3k�>3'�u3J�S3)<-3��2�O3�3�63�O�3��3j�L3��2��\33�)3q��3�iF3��13�O-3m;:3A['3�Ժ2Xm?3��C3t�2x�3�ҙ3xJ3��a30k63y�23�*3���3�q�3��"3Ҹ�3Ǿ�2��t3I3�L"3u��33�3�k3҉3d�)3<Q;3>��3�)d3�n�23^3�(�3��k3A�3�u�2R�`3��3�CO3��>3���2���2�3qf�3� 3N��2:j�2"8�3��p3e\3y�v3?�^3rQ%3��!3;�L3+�2�cV3���30,�3��'3D��20��3.aY3��Y3�5s3�	�2���2�L@3�E�3��2��2�K3}��3�Ӌ3`��3Yx3-�>3"�q3�J^3��3���2�5E3�2�3���3���3b�2-��38�F33z+93go
3�r�3s~43)��3�2Q3Գ
3�Q3j�3(m3�R3�
�3�0"3O(%3x3Y3��3�M�2	 �31�4]�3qR�3�3�;3�*�3e��2P3/;#3M�3��2�3�3S>3�3CH43"QB3���2[8u3�T.3<�#3�د2uS+3̅>3�p3�E3���3sR�3 �/3n*3~�3�=\3�k3��v3h�2.'k3�N�23@3�@-3��a3S8W3Z�3�13�eW3��73�3���2&�z3��$3í3�>3��3R`43`�3�3��}3�?3� 3=݃3+�&3IHt3��3��3�$3t�N3ͪk3`�3��T3�=3�y�2�3���3�+`3캦3Yh93e�38�3�?�3�-3��20v3�g63i�;3;M-3m(Y3d�{3w�33U��3�:z3���3FO63ۙ4��03lq�2��m3A�(3�=3R�W3�h3ؓ2�P3���30!�3|�S3�3�3{�N3��3Rh3��]3��p3��W3y}T3]$s3�Nv3�3I�4���2y1.3�\3�^�2pb3�|3��3j3 �24|TM3��+3��
3Pr3��a3jn3#&3�3�ے3C��2j��3�^3�3յ�2Q��3��
3b��23|3��X3<3]=3�/3z��2Y|3+B�3:��3�W3t��2��G3��A3�3 ��3Nb�2�̡3:�&3t�3
� 3{!3��,3��3��)3b6Y3D=3uT3p�3@e:3;�=3`��2�53�_�3�o�3�i�3V��2�Wa3dBZ3Ea3InJ3�3/tF3$3���3��T3=V3)��2�^�3��39�63�T3��N3� 3ʶ3�`3��2��P3oG�3�>�3��3�X�2(��3_�	3R3���3�	3�<3�S+3�Ճ3�=�2^h%3�#r3?��3�w3e�3�h$3��?3� 3���3s�l3r��2�[&3e��3�cK3q%^3g`�2�T�3;&3��839�3(��2�aL3�a�2�	�3,��2�3G�53���3}3�o3�i3.,3+s53lA3�^3ƨ�2���2q2�3��j3�S3-�2�M3���3[223��I3��3$�3���2��M3K-e3Գ�2X��2��3��/3G%3:�3w'3&s3f�63��3��3uI�3۠73�P�3>�3ޒ�2�5�3uAH3�Y�2L�R3�*�2�G|3>�13�L3/��3�,�3͑N3�A�3b�+3R*?3��3@��3�"�3�3�}�3�+�3�\-3܌�3Z�3��3	>3���3��3[��2�w�3�2�3�[�3J�"3�ݟ3�Ũ3~�>3x�/3u�3�O3Qt�3�v3��t3D�J3�c�3�0�3�;3�Ij3(�d3���3�FP3��2�	�3�,e3"�2�π3e��2{-I3*�>3���3��33�v�3y�n3з?4�tf3u�3��P3��@3�
3�:c3��3�e3?*c3�3:��3��3:�2�5f3�3*3���2[Ȋ3o3^��3C�3�r_3��l3Q�3OW3� 4��*3Tb(3i�2f�_3(�;3m0�3�0[3y?3&��3hɲ3�#�3�G�2FS�2��r3���30�-3��3's_3�ȑ3>!37m�3��2��3��V3y�3{a33�4}3\��3��3��3jD;3���3I�3�F3�b�3�� 4Fw3�� 3��3�3pm+3��3�z,3���3V�33�4�g}3�
C3�r3�4��`3�g�2�l�3@�}3q4.3�q%3#�3P��2��r3��}3��3��u3�,,3�C3���3�!�2t�q3w�3��3��A3r�_3MS3��?3(�K3)�3$�n3�e3dzu3��G3[V`3���3��V3~�V3@zU3���3�WP3�Z3��N3��F3<� 3{��3G�p3ӌ3��J3��c3])�3K�3�=*3(�'3s�"4iT3���3�w3�]V3�~3�w3��l3>�2ڙ�3V��3�3��3"{�2��3%��3(3�1�3���2(�o3�63�"�3�>@3�B3��3O�4�s�3y�3mKg3���2~�y3��3��13j� 3�W3���3_M93�	�3?�3�J3�c3,��3�"3<�b3���3���2�˃3
�3���2�_<3�@�3�q3XR:3�_�2.�2�-Q3�33�@�3hn3�2S3� �3���3��3V�3���3��!3��2u��3�Բ2�%�3dנ3�/�3	 W3�1�3���3�E4c�3�4�3���3q�(4"��3���3^�3-�3�֜3P�4t��3z$�3��R3��>4���3�k43�(�3Ӿ3p,�3��P3��3}��3��3��3n��3YD3�f�3�F�3��3�ߥ3���3��3#��3Z�3K�,4|#�3p2�3���3�2�3�Nu3�4v3��3�y�3��|3"�3s%"4�E�3!�3_��3�4���3�a�3S��3�o�3��3W�J3
d�3�S3�ض3{�4�M�3��x3�~3"�3�5�3�o�33���3�H�3���3��3���3�S�3:�3�-�3c��3��3�y�3��3o"_3��W3?�X3�-3��3Y4JY�3O��3�]3+�3�s�3U�3�{�3��3
=�3��d3}�3�j3�uQ3m��3(o40��3���3|��3�=3�w�3Z�3/3���3mȻ3��47J4�3�*�3�j4^;4mٕ3>��3cVt3��3~�3�ð3��3�3'�4���3e��3�^�3��3��3�3�O�3^�3LP3V��3XkI4Ӌ4�L�3�x3gֲ3�4���3U�\3���3Rv4��3rt�3$W�3!�D3�^3Z4�y�3F��34�v3��y3�J�3Fs�3���3k&3x��3�� 4���3��3Z3�Dp3g��3 O�3��
4g�@3:�3��3_au3�0{3c3¿3�C4�/�3Y��3�u3�3)�3_�4��3H�m3�Ϯ3Gk�3_��3���3��#35K�3��3�y�3�ա3Z�H3�3�9�3\I4�ա3.��3P�3��74�q[3W7�3LR�3�x�3�OU3�`�3���3���3���3qZ*4�i3��3sgs3��3�3 ��3�A�3�y�3} �3-i3���3&�3�J3(_z3�Nf4ջ�3ٹ�3��3u�3)�e3�H,3:&t3�V?3>6�3�4���3rZ�373��3���3v�3��3��^3� 4�ފ3��
4)�33 �3C84|�4ki�3Y�3�a]3��=3��P3��3q{3\��3@��3F��3�g�3J�3,ә3��3a
X3�OB3�ؘ3¥�3�q�3�R�3P�4�4���3�Y3��4AS�3S�>3�A�3�=�3�m3;�y3֎�3��f3���3C�4�"�3�C�3%83D�3�t3�KA3Qk�3*43�3�i�3�#�3�-�3��O3K6�34	��3Z|�3��3/N4�!T3��4�̤3eD�3z�3o��3J�40
4FI�3�3>4�}�3���3yɲ3��4X��3���3>9p3X�l3hS�3s� 4Ma3�:�3�¢33)�>3���3�%�3B��3VD�3� 4�k4��3q�F3���3�έ3Fԏ3Õ�3�aU3��4[��3V|�3��o3�{o3D7c3�H�3}�M3���3˗3�O�3=p�3Ժ�3
X�3�O3�3�3��3~�3�g3�T
4j�3TtO3 `�3��r3nX�3��V3�9�3u��3��3iu3�1\4J.�3��3�(�3 ��3���3���3��3\�53/�m3a��3�x4{��3m�3Z��3�K�3���3��4ͼ43��4���3*��3R�3��3�3�T$4(�3�;�3��V3��)3�~�3�L4��3[�3�a�3��O46C4���3��X3�4E<�3��38�3�F�3� �3x�x34�4���3�[�3Q�3b��3H�^3[0�3�f3$wr3Ϲ3�ͽ3��3��3g�3P��3�4��w3j�T3�8�3��3��3.4�3���3j��3<Ҽ3�@�3܍�3nΡ3

�3�D<4A�3�D�3�6�3���3�̙3ͱ3�x�3D�_3B��3��4Fʉ3��3C�#3���3?|�3��3�033���3�T�3�)4���3�3�Z�3ßB4u�K3�j3�!�3y]�3�(>3&�p3���3�s&3�o3��4�ԍ3_>�3h�)3O��3�S�3�3M�3Nk3h��3�3�3�3|3he3y�2��3J[3��3��2f�e3$c�2/_Y3���2"�3V��2�&43Hf 3I�D3��2�S@3�  3}�2&��2�TE3�"3�835�3�B3Y>�2�$L3��[3��22�3��3���2��!3$*3iH=3[Q"3�j$3^�#3t"3��3xE�2D	&3�[�2sE�2�%3���2��2��2�k63V:�253ai�2�i3O3$�"3�k�2�*3�ޜ2M��2{ 3oߓ2��2�ڗ3��v3��3;��2�s3��R3h3��3:��2�33E�2VG3=��2=�Y3�W3�^�3l�3/��2�%B3<w�2e�3ǀ�2e�y3�H3K��3kHw3ј2*��2t�2�O�3�j�2���2/ 3��2�O3r�3�3Z �2D��2d�	3w"`3zV�2�� 3RH�2vT�2��*3��N3
�2�!�2&��2�33��]3��2��2Z'm3Z�%3���2�T3<%3�h&3/� 3v�13��2�35� 3��3�b�2�03�*3�5�2B�3��35�2m�2��3 d�3eǑ3b��2I{�2F]3�Qg3~Q�203v�2dKI3'=:3 �3@93j�3���2�CN3D��2�{�2n:
3��2JD3�='3L�s3�3Ȧ#3�l�3�g3���2݅3�y 33K�2n(�2f�!3=q�2W(30�2\9I3���2^m
3=؅2�ݮ3>�3�]�2�~ 3C�2?��2o�3�h�3���2u��2��c3�=3��A3��2<#3y��2Tb�2�Y3\�2v7I3�@�2z[;3a%3}3Z��2��3zH�2|�A3��83T�2i�2�[3��-3�%r2�^"3?5�3W3�(33��2o�+3t�
3�!3e3>�3�>3
��2�)�39��2՛�2�ӆ2] �3�3�2��2n�k3��20
�2̸�2�l<3�k�2��/3��'38P53Go3��2��3_3�H�2q�|3��2��3��23�3%J3UU�3J/e3S�3zI?3C�!3��n3���3%��2=�Y3�Y[3���2�Z�3�u4�Z�3�_m3��2[�3��y3ο�2�k3��`3��3kv�2�vX3PY>3'R3R�*3�o�3l0�3ξU3�Yy3	g,3S3�\$3��c3*=&3D�S3��3?�o3��2��2��3�OR3��3 �3�W#3�Yo3䠯2��g3�M�2��3�e3�3�)^302x3d�p38H�3>��2i��2:�3�3�&�3�
�3��[3��3v3md3��<3S��2���3%��2�b3��3�@�3&�3!�38�63���3o�N3�;3��3��2M�3@<3$�-3v�K3�d^3��39��3�/3"��2���3�%43�2�,C3���2ef3U"3s��3�D3]3ږ�2��4���3(/43�<�3�'3�:3�Us3hU3��3��L3�a�3��3;2�3�]3�V�3��"3��2���3�v3{��3�~�3l�3&�93p<~3��3���3w�+3'Z�3��13�dq3A��3b~P3�f<3n�3ƻK34�%4vG�3q�g3���2~8\3�S�3�R:3��$3�cT3���3�33�_�3 h�3��3�3�N4�\382;3(��3MPN3��2`{V3�?G3��3�w3�53wΉ3pt3��2��)3�N�3]7t3Z�u3;�3^�y3��2_G(3�c+3��F3���2�4� 34�3~�3y@+33��2��3[V�3'��2��3�h�3�H3T^3'�3&ƞ3`�2��3dn�34�*3���3 g�2t^�3��:3!\3�3f0�3(�'3j��3�Oe3��'31Z3�)j3��33��A3n<^3.�3_y�3�d3�C3\��34â3��:3�_�3�3��U3��%3��N3o��2j�3�y�2է4ڕ3ZE39uR3P�i3W3�3�9@3��T3�30_4�+�3���2@��2��3�c�2[13W��3�,3�?y3M�93�+�3���2��p3PR3�*�3�I&3��3U�O3Ht3[F�2�uZ3h3	 (3�i�36ʡ3nT_3aRP3:� 3�3��3M��2���2�F;3r3�b<3Y��3��a3<�j3Տ�3��3y�73g�t3p�O3�s3>�'3��3�h3	�A3�cC3D�3�7�3���3}4�2N&F3=�K3�%3�À3b�d3�^_3��3Y�a3��R3`r�3K�<3<��3�]3a3�Rj3��_3���2z{3';3�R3��3��3�[3n3x�13)ΰ3���3�NL3�*j3��3z	J3ϻo31C�3xGM3��*3[�+3�d4d|�2��K3��?3;Lu3a43��3�ζ3/q3t	13��3*r�3��3��2��A3ӷ|3�Q	3�Bf33�3XU<3\�4�m+3�so3a�h3���3$
+3�q3�Z3�3NR3s�W3E}�3Ő!3A޳3X��3O�`3/"3E�3���3(�T3�gJ3�b&3�-)3Q�3E�$3G2x3��3��3�܇3���3ьS3�3�S{3��3��J3<�.3�'�3�,3��3�=�3{�y3E	�3�7Q3jv�3��3Fa!3�5^3{�13<I�333��3'�J3�a3d�U3w��3[R3���3��3�J3d�U3�3�Y�3� 3A*}3�#�3!{23�9�3} 3U6�3�)3�3�v3�33�Q3��N3���3�R3`w|3IW�3��4��3��3z}3�o3>J3b�j3-s33C��3��73��3?�3Dɚ3���2�63�83<e�3�p�3�S�2�)3%�J3~�3_3#3갍3���38P63�T3�N3�ނ3��/3� �3�ap3ҴL3	��3���3�ӯ3i�v3�&3ڶh3��Z3x+j3y$�3�63=5�3�3�3c(a3y+,3�>*3�oK4�O[3z�3-l{3��G3�,37�3ʂ3�;�2?��3;��3_�3���3ם�2���3�Ed3�j13	}S3��2�k�3�[3E�3F��3�V'4�E3w
�3eE�3���3{�3
�
4�JA3��3#�Y3���38r�3{6n4s�3~�B3bO*3��4�4SL3��3\A�3�_�31._3?�3%��3�>4DF�3��W4��3嗇3���3�F/4�Z�3Ҫ�3��4��39�3��"4Xr4$�%4"LI3�z�38�3��3��4�v3$��3[`4q4�#�3��3�f>3ˠ�3�^�34P>44U3V�3jr�3��S3CR�3S��3)�3N�}4���3�f�3�R3s�3���3��3�
�3��3-�3�k�3J4ꓚ3��4i��3h�4ߑM3�	=3�3�3yf�3�V�3��Z3X²3�3�e3�.N4���33*bH3��4��3��3�b�3�3Q �3�4$3G<�3 53�?�31�63�c�3�V4%��3�g�3,,�3��3���4�o�3ߨ3qY�3B�4�0�35��3��y3m�3ɱ4�\�3�@4��3���3��3H�144ۮ3��3"�53�v4	z�3���3!�;4r��3�ϫ3��3��p3ɸ�3�*54AV�4�R�3OH�3h�J3<�3�J�3ުB35��3i�3��3[�,4��R4���39��3*Ч3�+�4~2�3���3�G�3_�3�7�3�	4���3���3k4%G4���3�x�3��`3��!4�d4�8�3!�3xj�3��3iz�3%�33C�3��S4�3
�3<�o3��3[(�3�}`3V@>3���3�#!4igB3�J�3$v4y��3*� 4�<}3*�3�B4�;�3X˟3*�I3M�4��3&�4w�k3p��322�3 �$4�V�3��;3O%�3�&�3Vz�3��3&&4$#63 R�35�'4��3c�3;�3� �3��3F��3S�o34�T32�4��3T4b_�3X�u3�<h3�yn4��3�g�3��3dGf3���35Ŭ3��3s3���3\�3�G=4�"�3�73��35P3�S�21��3s�K3�A�3Wb�3�H�3�I�3y��3�3��3�z3OJH3y�3�z36�&3n�x3��F3�"�3p�a3c��3%�_3d�^3�;3��L3��3��3u!*35W�3��v3��+3���3�%�3�h23��3�ˬ3�?3*=�3;\�3��d3�"p3Kg�3n|3��=3]2o3*(4�zO3q �3$!�2�fZ3Z3�6%3�-�3V�^3
T3�(3�X�3��13�@3I�F3Nt�3W΀3��g3<Rv3��J3��*3�3�nz3f783��3{��3a�`3D�:3m�.3�|�3�9h3�`3��3:%3=�X3��'3�˵37��3ox�3l �3�Z�3}R3no638�:3�q3�x3R�3���3��u3� �3�34�b�3A)j3[3��d3���3̼.3��3,o3���3��*3�'=38f
3I�i3��P3#��3$e3!�K3�\�3rL�2�53�~�3�+�3P9i3w�3�6�3ٿ�3��
3��@3�Q�3�K~3ʊ3�Z3�73k��3%&3\��3=�;3|f�3{p3��4|��3�d3�-O3��3��3ːW37@�3��3��}3TV�3�D�3w��3xF�3�3���3u*3�,�3��3��n3��3aO3K1X3�~83e�2��3=�23���3�zI3�rk3D�3*�3� O3��U34�O3�]�3�1�3��3�823jQ�3��%3�t3D-M3UE3�׍3ĺM3C	q3گ13S�!3��3�d�33��Y3�e3'Ad3�3�m83g�3�%3�s3j� 4�j36�3WL*3�(�3ct�3k��21fU3I�3޼P3>��2��3��3�=3�rx3|�-4u�L3��3啁3:S3(\3D�*3!�R3�
I3�-�3� 46�3��3@��2��<3��3��3ʰa3�s3�`�3{��2iH�3Ђ 3�u�2�$3�B4{�3'�P3fh�3a��3�3�i?3�x3��37��3�Y�3�h3�.3��&3*�D3��]32�o32�`3���2s�j3J3�Z�3�3�3�Q|3l�3��3t39�o3:[�3��03C�3 �3&�3�:'3[�3�?�36��3��-3��3�ʏ3�u�2(a�2e4�3m�@3�#�2Q�3o��3�e3.~V3X*4{�)3Z�a3���3�]34�3���3"D�3k%?3�n73d�3� �3�xy3��
3O*�3��;3�63!)\3�[/3̣N3d��2bu�3AO�38�~3�C39B|3��#3�P3�3b�3��28�y3��38)Q3��T3jd�3���3:��3s��2xG3k��37�	3E�3�<N3��^3*�]38�83��w3��o3��2���3~�~3�Z3S�3`3� 3,'3�8�3�&3A�q3�Z4�53��P3�D�2n�3�m53��2vE�3�M$3#9�3���2�&�3G23�(�2���3�T4XV�3��	3��Q3�͞3��;3�3�3F�:3lj.3ھ`3I;4)C�3�3}�	3s�3:A�3�'T3�y3��E3�%h3�F34Õ3��z3��E3l.w3A��3�ԉ3w�*3�3�9G3:�M3̛_3��3c�3���3�}3-�3�S�2 {B3ڥ�3M�3`�33:3��"3��x3�\3V��3��|3�L3���3�G4�893.�3EQ'3 ��3��"3uף3�3TA�3ֵ�3��3Aֱ3�H'3�83�=H3Y��3+0�3k�3AB3n��3�?�2	�3m��3��N3�%�2Th$4$�X3�Oh3��3f'3^�\3�wp3�U�3J�3�e�3��3�3w�c3gi
39��3�Y3h�3��a3�W3���3v��2��3�83�I'3�x3_44K�3zV�3[&53+pA3�Q 3�r�3t�3��$3:m3��3�_v3�V�3k7�2d|-3t��32�3��3��	3,��3R��3��3�wA3���33�!3���3�s3*�3�^3W3_�o3�u�3��3�3k�3��3h�3�U�3�3�io3Aa]3`%3F�3�KC3[��3W��3�l�38��3 ͘3��x3�.�3�^43�^�3s)�34�^S3�v�3^��3�ۉ3,|�3i��3N+�3ˍd3_u3�p�3ư73�093mɇ3s�(3�_�3:33�.�3��3���3J~3�$4Zb3�o3���3�h�3Y�3 ˊ3�Z�3�X3gG�3�/$4��3c��3I�3��3���3gk�3���3G�3�n�3�(3��3D;`3�V�3�O�3�"4��'3R�3<�3�\�3=3 ��3�m�3��3t�s3���3U��3�AG3�13(��3�Ǖ3뽇3�M�3��^3<W�3�k3�^4���3��|3m�g3�k4��*3��3sݺ38`�3��3���3&�4mq-3qx4�34Z{�3ZP�3�`�3~i34b�3�>'3���3�E�3���3 �d3wr4�O�3	^3!D�3��	4�A3��3z�3U�&3�`u3���3��3w�M3^�3�3��3��3	_�3<��3��3K+=3TF�3�-�3��3"]3~�3�.�3� |3���3��&4H�a3�nm3��3�jc3�GP3�e�3 ��3��3�[�3Y
�3�7�3�X�3@o3}4E44i%3yj�3��3�s3�RF3�\�3Qe�3-X3+~R3��4}}�3YRp3��3�L�3�a�3���3X�3=TD3V)�3A��3-~�3��3"�3	��3�s3�Z�39��3�O3���3`*!3�T4�r�3[dB3�`�3��	4��?3M�H3��k3��3�U3`5�32-�3م�3���3��4�p�3�ل3��2.�3��3��3.��3	�j3�W3We3)�4�8�3,"�3v��3��A4᝕3yhy3��4a�83�$�3e�3�ܲ3�W`3��3B��3yJ�3�f�3%:[33��3�3N�3C
�3�43A��3W�3�Jd3ZZ�3��3EQ3c� 44�[3oG�3���3���3g�t3X�3�?3C�K3�a�3�ȫ3`Db3�/
4h�P3���3�Ԍ3��-3�;�3��%3���3�bI3���3e3d�3Y@3�Դ3w�3��t3��35�V3	B>3��36}3�3v�3B�4�i�3� �3^�p3C��3�>�3>�M3��X3�|�3�Sv3NO13|ь3z��3F[s3D��3��3שL3X��3? �3[0Z3b3~�q3�,�3�0e3��3�:�3��3��3c��2��3��3麄2%�3�`�30ʳ3��(3���3�O�3�Sk3�H�2a�3s3T֧3�n3%�3�0�2&g3I��3�+3|S[3���3ayc3z]?3�M�2�oF3��;3��3&�v3a9u3=��37�
3�3t�I3n�q3��g3m��3�_3���3/c�3ź�3[s$3��%3��3FԎ3��3�ܩ3A#�3&�G3�a�2�X�3U53;2<3A�^3\|M3��c3=j3��K3�x�3�F)3�z�2cQ4�݂3�N-3�/3|Ƀ3S!13�#_3~6b3�3�qY3��F3�u�3{��3g�3���3A�f3��2���3A�c3rY�3��28��3�3If�3��3�o4�gV3�*�3㴗3aBF3���2��3S>K3t113N-3��3{)�3�M,3��	3�Jl3�\�3�9�3K�F3 ^F3a�:3'Z:3���3"43�73G3��3�83�^3��93+�Q3�4�3V�3O�d3D�]33��4bK�3��3�83̡3%�D3�y93M҉3���2e�P3��3�3�3�3��*3E��3#fE3E�T3���3�(�3�	�2�_i3��3��;3�R�3�?74�f3�GI3n 3%HX3j�3���2��$3]S#3�.�3��D3R��3/B^3�X3ņ3�'�3a30�3�I�3lU�3r E3;+c3��13Ot3�*3з4��i3��+3fe�2��2�63�.�3D�3kP3��h3V7�2L��3fO34o3���2�&�3�*3�zG3;`�3��N3J�,3+e�3��g3$�
3�ah3�7�3�˄3,�q3�qE3!K�36�G3��32�3o�3��3׀�2�3�3j3:� 3Ѵ3$0�3k�N3r 38��3C�b3���3�G>3v}43x�d37�3��e3�s3FW�3,�k30�3�M
3�v"3�L3oq3<M3��2��3��W3��C3Ӭ43��4h�(3~O3�Ӟ3�3��3-��3"U3<3�t�2�+�3c�3b<3!h3y )3<+3�3� �3��3��=3^T33�R�3 rx3 ,3��/3���3Ri3��3�&3��}3	p3��d3fb;3��3�@3vȌ3ɝE3j4~3B(3D��3��`3D�A3�a3��3�!+3�c�3
 �3��T34��3@ 53���33*�2XtD3�~�3�{3|;3��O3J3�H�2{�v3��3j�j3��E3��93��3�W/3~"3�M3�m�2,�3�2O[�3ta�2�2/3H�+3���3�_r3"�J3[2�3գ3��@3�d3o�{3��2��3ח�3�ox36N3�Ĩ2�3�:x3���2�ԉ3�=Y3ϯ?3�W&3�O~3E�#3��3��Q3犵3dHs3)C�2p�3��>3�"3�3�PO3��(3b~3&4���3�\33X�83�,[3@f�3��3p73+JC3S��3�hD39h�3v��2�!W3��>34��3��3PU:3r�3w@t3."3�83ڹm3�3��3?��3#f�3��$3,�2���3�3h5-3�Ԝ3��2��:3�3�bQ3�,Q39F3
.F3dH�3a�(3y�F3W#3��'3�H3z�&3��3�� 3��;3�x�3��t3puH3y�q3�N<3��3k3s�l3G�+3��3F,3��"3�.�3$L3�8I3�%�3\3��332�3���2��3�;3��h3��3�#3u�3P�3��,3�	3��g3ױ�3yg3�sW3`�?3��3޲�2�:�3
�C3�i�2m
3l 4�6e3ڍ3z9�3v��3�d3�L3(�30�3��q3��3"��3��73/G�2T1X3� 3�2\33z�2^Ut3l*3I�3x�23RW303-�F36J�2�3���2�3.d�2� �2�A3lVC3�u�2Bc�3��j3�jj3k�+3v��3�8"3��2 ��2�F	3C34��2�j3��203Ɇ3j`�3�3��2ۛ�2"��2c�"3��q3�[3�um3L|*3�}�383��P3C9�2$�;3Q 3;px2��2-DG3�3�53��#3K�/3��=3{53��3�U3A�3�a30(V3��2�3f�<3� 3��2�Fy3y� 3�93V;�2E�2��:3���2�Y3��93�G3�e�26�.3�433�39�3C/�3�3L�'3��,33 ^3��2f�3 ��2�3�3�_3TZ]3��2���2:�3]wB3|�3�,'3�s/3���2K�^3J)3�^�2i�3�E�3�d:3m2&3;H3ͮ2C�20��3d�3�+�2~[	3�93�u3'�#3F�2V�D3T�2�3:�n3:�3�D3�}�2�+3�C�2p�3S3?��3Cu3w�3��.3�u3��3�<�3���2�L13�A3��3��-3\�3^��2�3*3��c3�=3��2�gI3��3H��2j�2{/W3�3�,�3�y)3��3�?,3��3<�3&�V3P/3��2�53���3Gwd3�l33�?�2��j3!�G3���2�g3l�2�3`�3(r23��%3�3�7�2�k�3���2��A3���2�,�2)�,3�N3T`3��3�3�!X3-�3�A?3��2;P33�2��2D�3C��2�F�3�3Ճ 3�i,3���2��3<��3܂m3Hr�2�s�2:W3�_�2��a35�:3g�2&�3�ׄ3vvE3��3��]2���2�~�2߃u3�m35C�2�(3^p3΂�3���2z�2lm�2)�|3���2�&�2.1�3��:3?3�6!3v�.3���2�P3Q�3|s39s3�J)3h�(3�;3(c3�s3\�2L,�3Ew3*�53��&3%�3�iC3��3�Sc3]�3�K�3���38�3C�3�<�3� 3�J3G��3z�3�!�3*�_3jh�3��3�.3��l37v�3��O3,3Gݜ3�3k��3:]�3��36�q3��3(�3Q�3 ��3� �36�3�ol3�`�3|��3-��3��3N'_3j��3��C3m�3��3TZ�3�A�3�?�3wW�33���3�3��,4ҙm3�Gi3�A73-�3��3�^3ag3up�2q�3�3'U�305�2��3��3���3*535��3�3�3a�3�S3���3�KX3_�i31_�3M�4��)3���3�7�3U�z3ֈ�3,J�3IS3��3���3ݘ4ED�3�;\3G3Ⲙ3��3p$3��3��3�-B3�&�20��3� 3�`�3���2/��3�743��3��2{P�3�:P3�Ff3$ݼ3�$�2&�3+�'4��3��D3��(3���3	{�3�'3S��3ʰR3��3�4L3:5�3�E3�30�3H�3��
4C�3H{�32t�3o �3�q�3J��3�)H3�N@3w4[�3'�3-r3�^�3�V4�S3�9�3�#3�Q�3rX3^��3"	4�jq3%Z3l�-4�'�31C�3�]w3��$3_OG3@�r3�=�3�?K3�ϐ3���3��3�ԙ30i3w�3v@�3O03w�3��(3Nz�3�f3;��3g�3��3с�3�]�3�x3�S�3��L3 a�3�v�3$��3���3�?3)��3�64��	4��3�
C3���3�~3��3��3v�3wq�3��3b�3D��3B?36A|3�.C4��3�U3�o3�z�3���3dl�3o�3S�>3+��3���3���3���3�03��<3pK3߹,3%��3�]�2�R48�U3u�J3"҇3�	�2c��3pt4��2�P�3:�73,!v3�B3�vM3hD�3�P3��3O��3�,�31ׇ3��3נ�3�3�3�و3��3�v35�63��3�:t3�|3e��3�I�3���3�C3�I<3m|z3�:�2H�3qR�3%k3�JG3-�3��~3"=�3�V�32��3m�"3�m�3�K93er3���2ӭ�2��3�yd3B�3�V^3��3�f�3�/�3`f73t�d3�&+33�~q3�F�3c�^3��3��3�[C3��#3���3J�_3�ߦ336�E34��3!�a3�&�3� X3��3��3ߐ�3�3k��2n�h3F�3�W32�/3͙�3�u�2��w3r�-4}`�3�3h!a3~��3
g�2��3[�3;�3��q3n�53/V�36w3!�d3;�2���3s�k3*�3`��3��3x@13)�3׬3��3sgZ3]��3��3މ�3d�3�ex3�wR3��3��i3n�&3�I�3[�$3�s�3��z3^�"3��3'�3WD3�3�}E3vo3��3�u3|M3�>G3��73aN�3Ye�3��93'3�7�3NT3��*3Y�4�Dx3��m3���3[�3=�X3�Ŧ3��*3�|4=6v3t^�3��:3獢3�v3{)L3m��3�3��3]8�3P��3���3��;3vf3�1z3��Q3���3��[3���3Ć)3Rkw3�v)3+\�3��E3��4]lx3�*�3<�3�Wx3�*3���3��3:�(3�r�3���3�R�3;iR3��03��3�e3x#3sۣ3� :3<��3�w3��3P��3IL3;^�3;J�3�Fy3��H3�޻3}3&�83��3�G3��13��3��3��3�[�3��_3�~�3;�o3�^3Է�3�[`3�p�3q+I3���3'�3�C$3��/3}0:4p��3�p|3 J�3�u�3��c3�+�3�ʣ3�j3vH�3\��3`�3��N3��3��Z3v�t3�*3�m�3��.3��3e��3�	�3V�p3k��3��26�14F�"3�`3�DS3;tF3�C%3Mq3���3��2xa�3F�3׆�3Qo13�=3H��3�*�3�63���3�u>3�f�3�,"3T#�3Y�m3)7�3x�3��h3�f83�u3�z�3���36�;3/`�3�x23�b3�=W3�8�33�3+�F33�W3,�3�k�3��*3a݄3!�"3+�p3�93�\�3Hw3�0�3U�3�غ3��W3o�l3t�3�=U3�y3B%@3�$�3��&3�C3�3Tk�3��c3w)�2	f�3H~�3��3�S30��3�ɟ3��,3\}�3I|3T�c3$�3���36�3��3�a\3M	�3]�j3��p3��3S��3W�3���3�ݑ3���3Z13��3��P3��3�ݙ3Y�(3\j36X3v��3	?�3��a3��p3}2�3#�e3w�r31T3�Z3|��2��O3�W�3p�3r+B3�=�3ë�3K,3�'3�3Kb3g93?��3wV3���3��+3�3oq3-W3Ū?3AϜ3ݐ�3Q�P3�d3�Lg3�+Z3�֎3{6�3_!&3��&3ϟ�3��3��A3�MS3~V3Uc�3�L-3�V�3A�3��23:53�wI3��k3��U3���3�D$4�Bz3�Gr3機3n�e3)�J3��y3
�3��3
�S3!:�3c�3NF�30R3䢠3Y��3�� 3��63?pI3/@�3@S3��3�%H3%ڄ3U�2���3�^3e@b3��,3eRI3�3�{g3�h�3NA3PZ�3g�38�3b�3�03Ё3So3�Q3�{3�]63�}j3-:"3�5�3�k3�8i3Ia<3�h44�l3��3�73p.3��d3j��3�s3_�3�G3ɹ�3&�3��a3��3��3�Dr3d�3D>�3���2�̗3�G�3���3OeF3A�63��~3�G4��i3��"3E�3��/3��a3��36i3�` 3���3
`�3�3�3Y�3k�D3���3�٥3�'c3HK;3F43��3?>[3�ն3#9+3��3�'^3�K�3�#3��3'�3��03��+3t�X3�՚3�3k�3���3Ͷ�3eX13]d93%׃3|�n3���2�'39E�2��3Tv34��3~O3^[�3�Ev3�4�31�3�rn3˦?3QA3k��2��31�h3^T$3���3`��3r�m36:�3��D3mk�3E�630�3�+q3ޢt3.�s3]nF3o��3��o3B9�3Iʾ3���3���3gӘ3J�_3�/�3�
�3��r3:3�3�M~3�QW3�0�3A��3��3��3�3C��3��B3�l�3[g3��n3��3��3u�D3#�f33T43�k�3M�N3�L]3�c31�;3Y3R�p3�~�3��3]y�3?"�3TA�3C}�3�Z#32��3���3Z�3$>p3��[3a�3G3�3&&.3!�v3���3��4L�L3'�3��3��<3�J<32Di33�3��3yI�3�B�3E�3�[�3��3(c3��3Ʌ�212K3�\^3r*e3�x3co;3�C23��3(�Z3���3�30B3�\53��3�Qt3��3�m[3�.3�3T�-411�3wY3~��2ue�3k�~3�*�2�z�3Z�3r��3	��3��4�}3�u3�$3�3`�3)�833};�3��M3f"h3�4�3���2�^3ɭ3��O3��K3��2�=�3�P�3d�3z�2k�-3ׯv3Hd�2Ӎ�3�zy3C1�2"��2��3�� 3�τ3��3
�/3�
3^3z?33�B3oz3���3ǘ}3�3re3�O3��J3�2�dZ3��2���3�63��B3�Gb3���3ɇ3|�3yT3�l%3^a3��D3�_3��P3p�3�@!3�63='�3=X�3��	3�h#383�3w=�3��3���3�	;3A��3tQ3�3�m3�3 w3W�4Rw3G�3GP93��M3-93ݰ"3�Ԑ3�s3��3���3���3a�j3�e�2K�E3�|�3�H3�OZ3ߥ�2�ҟ3�!3�3��3(b93�f�2��4*36�G3��3�,3�/3��M3�X�3a34�3.�32_�3�^f3�(:36q�3H1Y3%l3�u3S	3L�63�g3E��3��53��u3s� 3FR�3���2]U3���3⪅3b�.3|�Q3L�B3;t&3�-3$)73m��3��H3+�3�F�3|y63M�3��J3�;3�2p3Mr�2�/�3{�$3�GC3��&3��3͍�2{�3�j3*3ñ%3���3i[3D��3;K3�3jD�3T`�3f��2���3}�3oRg3X/3��2��3��3��>3�33�m3hV"3�*�3��2zl3���2H!�3�c�2��3*S3E��2��3���3��/3A;3��2?�k3�3Y�2�f3�:�2 *3�9�2�2�3�_3��Q3E 3�sk3�h3/HS3��}3�[�3��=3��03x��30�	3]�Q3��3��a3��j3��63�a3Gz�3�x�2��Z3�2h��3!}�2TZl3&�13�C]3��3+ti3S3�D3��3���2�U�3爲3Ʊ�3�m�22�:3=�3�۶3��33��G3�m�35763��3�$�3ְ3	�3C�<3[/y3̖)3-3���3���3כ�3
E73;�W3�d�3�#y3��
3�8�3=��2�23���3�I�33>`3�3��X36So3�!3��:3Jջ2xMm3�!&3�F3T�-3ǰ+3���3Dd�3ȴ\3^O3��J3h�3�:3٘23��73��-3vT3�ѹ3t�3d_3�"�2c��36�{3gk
3�l/3�)43�CC3�iZ3Љ�3�L3���3=�\3�g�3�x3N�]3�
:3��x3%X	3~3=4`3> 3�L3I��3bu3�Q�3��3+��3�F�3 ��2/�3�H3���3�i�2*n3�[�37�2�J3~E�3���2w�J3CVI3 83�G3�#�3�A3Q=3�n�3$_�3�R�3�z3��3:>3P�D3�}?3�93�LL3c�a3�&3:�&3Z�S3{Q�2ˬ3���3���2�q)3��<3Wu3'J�2�:3_�j3���2.3dM�3���3 �(32��2 �t3P�e3�E3(4�2��3+�Q32�2z��3��v3n��3`�{3�2�3l�&33�83ׂ3Ae33i��2�.�3��C3皉3)x\3v!�30�I3T��3�R	3�Y�3�3y�34�3� �3��\3�F3V	�3��g3�WP3��y3��3OI.3�ZT3|�K3*V�3T��3&�x32~�3�B%3@��3�/�3_}�3|W43��3�wJ3�l3��T3ׁN3�Y3��3?.3P��3�sr3��C3H2e3N�3c�/3��83�>h3w:R3�38�3|Wu3�BM3��^3�l�3۱�3n�G3gj%3�q3_�N3ag3�3 �g3eۻ3R�3���3!j3���3��>3v�4}I334�$3d�Y3�*3�/3'�3wA3�9�2ր�3�#4�r�3>�3x�I3��r3rm3[ٍ3u��3i-j3�Ħ3�\N3�E�3筍3d�M3�_3W,�3�u3�Uj3IQ�3l�s3ȁb3CV`3�3�&3��3��3�*w3�Y13	7J3q|M3I�d3��63��f3h�R3�o�3(�t30ג3���3��3�߬3��3zO43��3��.3�zg3oj3��c3��3��2,�3w��3�I�3�g3639e3~�3�e3��3K3�2s3v��2�Gh3s�M3R�23d��2�{O4��V3wr3�~Z3�$�3b�s32/�3_��3��3h:�3j�3��3{�d3�R�3-J3�3Zo3��3��3|J�3�o3s; 4�H�3��432�<3}��3��}3wMz3;�33'K3�c3ʵ�3�ܝ33 �2n�B3!��3���3D�S3�3�g�3C�m32�631̋3[�V3�'t3��:3q�3o��3�؈3�X3[`�3��3O@637�Z3?�L3�WK3%"t3&V]3�a�2�E�3��3��3i�3�L3΄3L��3��30�38�P3mS3wВ3��3��23eJ73�}/3&��3�?3���3��Z3$�t3�3w�73�/�3e��2 �3\�3���3���3{��2^f3��83c�.3��{3s�2�"�3v>3�Կ3��p3��3�H3AE45�3�o3ɋ�3KG�3��3l��3�Wk3/�3eWr3�J�3�l�3��31h3�14�w3 k3�|�3�D3�R�3�43u}�3���3��3���3C�!4��33K�3�^�3�Lg3[��3)��3��3G�z30�3z	4Xf�3N�3��H3�͎3�y3�f3�s�3���2a+�3cF�2@��3^�3���3
Dt3��3�'[37�3F?�3��4^��3��3�<�3� �26o�3Y�243��3v%�3�|3�l3��i3xZn3$�3�`@3uQ�3��3��4�3萦3�yk3�$�3R�_3^/�38��37�3�e�33�k3�.D3�_3M��3�\ 4�U3&�4:U83�3��3ø+3���3qA�3!4�/3�ڡ37F'3:)|3�qN3�42)�3��q3k�3��3��2�Qq3�r�3��3�g�3w!4Ǎ�3�İ3�K^3��3<�4��	3��3�?3���3]3�\�3�3-X�3�nU3�4Bt�3�$�3���39�3ʀ�3��O3II�3�A3��p3#4��4mr�3�xv3U��3�`�3Wζ3A9�3�A3
��3=�3��4Y��3�{3;�.3��H42J3�v�3��q3 �O3DSQ3�;U3!bu3���3XA�3{b45}�3�"83ը:3Ŕ�30X�3Pg�2�R3ʠ�3E��3ۧm3l�3z�3�X3�/�3�Z�3��[3���3�>K3W)3{�I3t��3���3�G73d�^3�a�3�M�3���3�@3c�3)��3z�c3|��3�k3T��3��T3��3���3d3��3��a4<�n3�32�3&�<3��3)�e3�Ǭ3`�J3:��3��4�^4y��3|�<3~�I3T��3�Ʋ3鋇3
�&3��3Jk3�.�3��o3��83@%=3q(4/�B3[:�3o;3m4�3��93�:�3�3]\^3�G�3�4K�3��p33ې3��3o��3�V3�3�3&��3�34׋3���3��G3��3��2���3��V3��g3��X3\SL3�R�2
�v3wK3���3��3r�3�GC3acx3¸039�3&|H3�3/63d6�2v�F3~�2���3��S31�p3��3S� 4�,3��k31�|3��3U$3>J3*�3�fO3l�c3�>�3�c3��r3�ʸ2l��3�3��%3��F3N83��3�s<3�m3�b3�A�3m�B3�)4��"3m�M3�s_3:c@3�:3!��2e��3�i�2�r33��3�6�3��3��2�c3�+s3��2*g83���2�]3ET3���3y+3=�3��H3�4_!�3��v3�4�31�93w�L3W�\3��3��3�ˢ3�4�k�3A�P3#D%3�6r3/�E3��,3�V3B�3"�3���2��3+�3�=3f��3�U�3��&3�-x3(mM37�2mX3F3勀3�p�2�P3a4���3�r3��C3"@S3�ŋ3"�>3�3��3��63E�3���3xQe3�|�3)]3`��3���2��l3�C�3/�j3"�3�s3�F3�o3K/d3 f�3�ɐ3X�3��3,��3��l3q3�l�3��H3�^3,�3GR�3`�P3�զ33Z3�3*513�T3(�23��3���3mn�3ȅ�3ƸK3ѥ�3�I�3xў3=W'3�*�2�Jx3ǽK3z,3��G3���2�Ɨ3� 3��3G-03d$3���3T$�3UPR3�s(3���3S�3\o	3o�3�v;3�3rYT3"ݷ3���3r(g3c�B3G�3~H�3p3�U3��"3�
=3!�2���3��3|b3��31�4y3PM�3�'�3W��3��z3x�=3�n]3��
3L��3��387}3|��3ѯ3�&3��3�W_3�=3�u�2Yю3�:3��3q@�3���2�3YǙ3�/3��-3��73�S�3��33�Z�3D�3r�2�PO3��3�'�3�>3�3�T%3�+E3��3�F�3��3�6W3Z��2ڃ�3��D3��_3�ˑ3�җ3��3OvX3I~;3O��36�63<3�3��P3�$Q3�X23�� 4@��3{��33N��3��)3��:3��3ca3�~3� <3��S3�[-34��3��3�A�3�13w;93D/�3n%t3eI�3��3��3���3�c35��3G(�3�.�3% 3ݫ3�NW3p�3,Յ3Mj?3�4�3�a]3\�3J@�3e��39K3|�4:3C �3��
3,�e3��93��T3Ko3*K!3�G�394� q3��93c�2z9|3��3"�2�L3��3�[3�y3u@4�%&3�;3�]3���3�P3�6031.�3���3�R3��(32ԇ3lE�2��f3^k�3KQ�3�ђ3��3'K�3�Z3*�2��P3J�2y7�3áp3��S3�So3z\3^�G3ږ�3NN3T�/3��13��3�~3���3�h3_��2�.&3.��3Py.3��D3�]3��3�.3���2,.	4���2�c3��3���3��2��[3|+3?�j3؊p3�y3�3�3T-�3��e3�ٛ3�VM3m��3aЖ3[��3�tL3�43��Q34�3�C�3�Τ3�3�c�3��&3�L�3�@3Q�)3��32 �3��P3$X3�lr3*��3�
�3���2�D3#�3�Z_3�Q�3�WI3M.73�5�2߳�3�y363P3�t93��3��~39j�3�e3�}h3��31�3Zzc3�lq3<?�3�f3[~C3�ZP3JR3o�3!V3��x3�^�3�~3���3�3�N�3V�3�L*32��33㶡33�X3�H3��Q3�PD3���2k��3$+�2��&32֗3 �G3e{&3�zR3ѣu3ڥ�2� �3j��3�j3���3eD�2CH^3w�s3�<%33*3�93s�3��-3��N3���3��2�3m��3ͨ=3&Va3�<3&3�/3�?3J�%3�7>3ܾ�33�3(��3��H3�q�2sV_3N"�3��3.�3�M/3B�S3ȂM3ǀ�3��3��83ƕI3	��3�p3}�3ey3��2U��2�[�3�a�3��3s�:3�҆3W�33�83���3wo�3���2~!3	�3�6g3z�3l�3��3�83��3DM�3jg)3�L3p�)3�y3tW_3��Q3��F3�q3�.3���3eap3��<3x3<?�33s> 3���2�
F3��3�lD3`@�3T3��+3��~3,�3�L�2�<3��(3��83e�-36�\3�'b3��3�+3
��3zg�30�3��3��?3�w43ܤ�2&r�3�v3k�3ؗ3��3ݎ-3��3�gi3=�4�B�3�]3���3Jq3hn�3H�L3�\3*a3��Z3.XO3Iv�3Q�|3��<39&3H[s3z�23	�r3�w�2�U3䝇3ܷ�3`3�3��R3�y3:��3��3��b3���2�Sg3,{I3�w3���2&��2p��3T�3.�!3��2H�l3X�s3Fh�2MEI3Yo@3i3�Iv329�3�#3�3�9$3O��3~)3�903��3Y�2��*3)~63M
�3�)3��3�-�3F�a3�U13,�#3��o3$�:3&�P3��B3C�3F�93���2�M3�43�+3���2M#4w?�3�|3\&<3�3SU�2Gٴ34t�3��O3��3���3q�X3��I3H�#31�e3�3�3"3�[13he3�3 3�t�3��3؅s3'v3=�3��A3<(3g�&3s�@3)~F3��43t?3���2A�J3�ں3�ob3���3�� 3f�3�l�36ǫ2
3�:3`�@3��(3�[�3��3zˀ3�3��3��X3a=�2��M3ހd3x�36m3�m3n�
3^^3a3�Z}3?+3�FJ3
�3�"n3s�;3{=m3�}
3�t3i�$3�'3�23h3N�3�v4ф:3��R3�b3�֡3p�2���3�/y3�v3|�C36\=3�(�3�UP3���2ަ53g�"3��'3�v-3v�r2�ҏ3<�	3- �3��3�Z�3d�q3�5�3��3�i3^d3C��3�U3]c�3M�3joH3o8k3-�3���3�_3�M?3v��3���3��3蠇3{�e3 "3�g3��4�;�3��3��g3^�4)�3ɣ{3�=@3	1�3�׼3GA�3��3��o3ũ�3��n3� �3�'�3qS�3ɕ3��w3��3/��3���3�.u3��63�u�3��3Z�|3��~3Л4Lp03ˬ�3�Z 3��3j.03^��3���3�'3܉�3~��3�,h3`S+30H�3��m33�3Sc3�U�3�(�3P$�3/�'3�33�3Y�3Pj3\?"4�[.37�V3��o3�F3�vy3��3�|�3�%�2��3@��3�_3!X�3�[43~Ü3�:t3�j63X�3�3
`�3yLm3�D 4E+�3��N3&\�3�J4"��2���3�g:3�2�3�'q3��h3��V3ɀ3�zF3�4�G�3N{�3��h3a�3Zj37�.3kt�3�q63���3`A3��3r%�3��3:�E32x74�pe3I>*3�(F3}�3p-�3.��3+�3@3�"�3��3���3:j3��\3i��3�/�3�`3��3�3V�3�0E3ER�3��.3s�j3g��3��3�~W3���3Bp]3�q3Vo3�Z�3�Q�3ʗ63�a�3vY�3��3_8�3ZI/3�~�3)�n3�R3�3��L3^�3�3��3���3�ژ3r�?3�G4�739F�3��!3ú�3c�~3�T{3i)�30L�3�4u3���3oD�3�h�3:��2��3^�4,�3�o�3��n3�?�3��[3�!�3b��3�?3k�C3!�3��V3��3?�3�Q3�Y3�u3ө3�3��3L�3[%�3v%�3q#3�	=3���3��<3f�30�3�,�3׳#3$�3�!�3E�
3pa3��4���2+Z�3��23 �A32�X3K�W3��v3Y�3��3YK�3t��3!	o3D� 39��3��L3�jF3��e3�3�ɠ3�C)3Lۨ3w�3N�2At�2�:3�lt2���2�}'2f1�2�;�2Y��2e��2c��2��15�3�Z�2ƹ�2*Ɔ2U�3B&�2�zS2��2��2_:�2n��2��2�ŷ2��y2�"^2�33���2/��2�T�2�M�2(��2s��2y�2W�E2��2;��2�3���2��p2��2
b�2�<�2�?�2z�2r��22.R2���2���2v�2��K25�j3Hxn2�s26BY21x2\�2��g2���2��&2�=�2�
�2z�2�C52��82��M2oZ�2��~2�[�2K�72�щ2,@2���2��2Y�[2�s2:qI3��"2�"�2[w2���2��k2��2F^�2�w2��d2��033��2\s�2i�2¯�2]�a2�I2&\�2p02�$�2�L�2t3¹�2�/T2���25�3b��2(��2U�23U�2��2�2�΅2�?2�Π2��.3�f2硿2a9�1�Lj2��3���2C>x2[u�2���2�J2�k�2P�Q2���29�B2;�3���2���29�2��2��2B�2u?�2� �2G��2�m"3�2���2��D2�r�2�x�2�%I2��2��g2Tϧ2,�1`�2���2Ԩ\2H�t2l>3z7z2Ο�2�R2�U�2'`p2�4�2��2x�M2%�_2���2��2�J�2�@d20�2�Nb2�/2���2�{ 2G,I2�`�2r�2!#�2��2��C2]f�2s>q2�O�2K��2p�2��N2$��2n�2U�42 	�2�Y3^��2���2hM29j�2k��2E�2- �2
�F2�k3��(2l3X�-24r2�!2��R3�}�2(}�2�#�2�d2ǁA2�4�2��~2%��2�2���2�Q�2�8�2xrd2���2�7�2��2{�&2.��2o��2��q25W 3�1e2s�k2��2��3�2ñ�2%�2%��2Y�72b�2��S28Y'2���2S�(3|��2C��2`*2��3���2r52f��2�Rt2#H�2�Hd2���2=�2m�3nd�3}[v33��E3I)3��'3��L3�Ǖ3r�-3!o%3t�?3��i3�^3FW�3{=3p��30L63ޞ!3r>L3�73<e3`�X3O�3
A3�z�3�y�3��3BԚ3��3qC3��33�n3�5�3�3��L3'��3g��3
�a3©63t,�3���3g'�3
�3?&[3<�3r%3�3b�F3�a#39*3f!�3{N*3E33�i3���3��2G�30�i3V393��S3j�3�N^3��<3/Fg3��_3�Hb3�J�2�3�"C3l�l3��93EО3��63� �3��K3�3N33B>3^xa3^&�3_�x32%3j�23Tt33��k3��3/RV3��?3v��2�D]3&%W3���2���3	w�2I��3�43�/#3\��2��2gq3�¾3�l�2�V%3�]W38�+3��>3C�s3�CU34p'3�E<3�6�3*;�3�m3���2Ӭ�3�B73���2ĎI3��2��3_x�2"�j3 �D3���3 �(3�m�3�F/38{�3�G3a3n�3G�3Ņ3�b3�P3���3z��3�zD3�M,3���3qW�3���2�@3��3lL3��3uY�3+3Z#�3�\3N��3CsJ3C"b3�c3��2h3�k3�I3r�3�l�3y�3K+�3[3��C3��3؄3��E3'̃35j13� �3[		3���3�'@3�y3\�;3��3u��3��O3�a�3��3�>L3R�k3!_�3�x3+�c3ƀ�3uC�3^`B3M�33@m3L�3�:33���3I@-3Ó35:3ǔ�3��G3A�]3HJ3��C4�hl3�=�3V�^3�P�2�@J3��J3R�?36w�2��W3���3�o�3�R�3.F3�R3z.�3A�3��c3��3��3r63M�3]�:3۝3�m�2��36��2^&3g�33�y3`��2|�3�3f�e3���3�1�3pSg3@i�2��3Lk�2G�2޼�3��3�d733A?3���3�5c3Β3��N3�s�3�N3]�B3b�+3��^3z`+3^��3�*�3�3��.3/�3LY�3d?w3@��2.3p3��3�q.3	�(3�Xf3�҄3�YY3�]�3�3,��3U��3��3��]3��R3衅3��3��3973@��3��x3�G3۸3v��3bxY3"W3�.�3]0�3/%=3��3H�P3�<{3AR3�(�3�{3E+�3�d35˯3��X3z=k3��3
�^3�ϐ3\�Z3BB{3���2��53���3�9�3�_3'3{��3Na�3��3��k3>�i3 1~34�K3Ld�3Q�[3�^�3Z\x3��4��t3��3��d31�z35:G3&͌3?��3bt+3�'3�y�3Ǝ�3j�13�s3���3K�3
?3ZZe3�`�3Cd�3�w.3��3��s3vee3Q�z3C�3�z*3
��3B�3��>3ۡ�3�^U3o,`3tq�2U3\v�3�*�3I<3&��2d��3���3S�Q3��m3a�53���3�j3Td�3��x36��3���3���3��|3of3��3�kv3�:q3Q��3�S�3f��2c�73���3=��3��32�K3/	�3�D3�N3�]�3��N3�E�30�s3	��3�Ì32j(3$gP3��4�yS3�Д3���3�9|3M)3���3r�3���3!ܓ3�Ӟ3\
4��p3��3Y�3b�W3��3��3t)�3�\q3C�z3���3ir3���3�.3
L4u-�3$"�3�	�3.�S3�%�3˔3䲁3Z6Q3k��3��3�{�3=ٝ3&3�3��39V�3�;�3�RZ3���3)E3�5�3=3F3%/>3��'3�N4��3���3�^�3y�.3D�Y3��H3-?�3��J3�ݧ3���3z&43	�3:B3Zi3��3�23�3]3�В3�tN3���3��p3�1�2��3(<�3��=3Ct3��3O�?3ud3��@3�Rw3�3���3j��3�g�3�qC3��2��3�7_3�W$3��32p3�}s3��53/&�3�FN3g��33;e3�o�3B�w3�$�3��3҄�3c}]3���3ka�3�#?3��<3���3��}3��4�t�3#[�3Y�d3��3�G�3��3�x3�>3-�3�Fq3��,3&�3}�<4�W�3���3=�/3
��3]&3���3o/�3K�T3^4�3j��3�m�3*��3D83��~3
jA3.�3�2#3�/\3�=�3�+3 ��3U�l3o��3�}:33+�3�8"3�i\3v�=3�w�3�ԉ3�3��37�3�dt3s:N4���3���3��q3��3ц�3a|�3�y3��g3} 4A�3��3E@�3R��3��U3�r�4�,43`Z`3z�3�NX3(R73�p�3�d�3�H3��3�4���3MUZ3ԙ�2��3��]3rd3��3�>3C=�3��]3�4v�O3	��3��2('�3装3�"�3�e�3ق^3�e3��3f�3��3�%�3?�4�?�3!��3��3~�3�c�3 �:3���3F�[3E��3���3�ڐ3�t3�i3�-Y3`��3?GZ3 s3�rm3�9(3��%3��3ڵ3��3d�3WT�3�ς3�C�36U3���3fߍ3�YD3�`�3j�3�/�3�K,3�e�3+�3:�G3�G3�4~.@3Co3G�^3u�3�Bf3`$�31�3m~3!�3P�3#��3z�H3$�>3�f�3��w3w�m3&�3(��2�v�3�J�3R��3�l�3��A35��3�R�3�p�3{�m3�h3��3�3���3r��3�v�3�#�3�6-4>��3��V3?�2��3���3�?3�3o0*3o�3F�3�B�3hV�3�:e3еp3?3e4�53� f3�*�3�ͦ3S��3�r3$S�3�FZ3��3p�3�84�̅3tD*32*�3�nG3��c3H/f3�
3b��3�M�36��3�@L3���3@�t3�%;4�37D�3�y�3��3�� 3��3���3G[3M��3v!�3�ɢ3��3�13�Y3��3��C3v�3��+3�+�3�d3yd�3�3��m36f�3�{&4�3�#3^#3��A3R�03)�38~3>��3sK^3��3X�p3ϙ�3�'3���3UA�3� E3Lf�3U0x3J�63��3�E�3��3�%�3��3��3�B3���3*�3�,�3��3��3Ln�3w"Q3Cg�3�k�3A��3U��3/�3Ҟ3q�3�� 3hp3?��3��g3ԗV3d��3�
V3A�3�pg3�P4��Y3Ͷ3�i�3��}3�GM3D��3���3��W3N��3�4�_�3�!X3S>3W�3rA�3�)3��Z3��X3���3�o3��3��3/�3�35�>4-�3/ߛ3�W3���2b�l3;��3�.�3�9Y3&%�36�'4�ɫ3$y35�'3`T�3��3\8:3U�H3�/3��3U`364�3��G36�/3R4A38��3M�(3��[3W.X3b?3��333��3>ԗ3̂�2y�Q3Jn�3&�3�F@3��2G6�3/��3��@3;�K3JE3��3g��2p�^3!A3��M3�Et3AI�3�|3�Q�3�/I3��3��U3�D3k�3�Q+3��k3 4���3�8`3wg 3'n�3|��30��3f��3�V3a��3�H3���3��>3>UK3�3�
:4Қ3Wom3P�93dL_3���3K�3�t�3��~3?f�3�ޤ3nl3Őp3��63s�Z3��3ΒB3��c3"�3~�N3��Q3}|�3�3��?3ځ3r�4c e3�h�3��3Wo134�l3�+�3�P�3�-k3�S3 �3y޾3%	a3��2x�}3��3F.f3=��3��3��3?}3UO�3��'3�!3�U33@4R�73,��3n��3�{j3I�{3�&�3B��3U{�3��3%��3ѓ�3p�3��2给3y�3^\O3�13!�Q3���3���3zu3�h�3*�2CS3K��3׹3��K3���2��e3-o(35kJ3��3�W�2�ʔ32��3�J�3مX32�:3B�3��3	�<3iZS3�>3B�33�� 3g-�3k�3\t.3
�[3��m3:23�\M3t�2�!l3���2U�63�o3�:s3.*w3��3���2��\3�$3��O3��3Ԙ3F�2��3%F3I¸2�/d3��)3��v3��/3>��3K�3#��24(�2��63EP3 %=3K�63N�3��03�FE31�b3XG3��)3\O>3*;�2Ve3;�_3q
3L�03/3��3M�3s��2	�2F��3P�G3*a�2���2��3�'3��J3_Vr3M23��23��3�3m��2�\3��<3��a3J&�2��3��#3}�R3HJ3r�U3�53y�3]�2;�3��21Z43VxC3U�2;�73�8m3�^3���2��53�W�3X�73@a3���2[33��(3�]�2v��20��2�NO3kh�2Q�|3 ��2��3~Z�2��3��I3��3)A3}�,3 �b3�E3�0;3Uy23$*3Z[�3�3j�3Lr�2��v3SP3�l3ڏr3�^43%n3�x93��N3Z313j?3�d,3�bl3;�3֘d3��3�A3��3V83��Q3.L�2)�2��O3��3sj93�2��/3eh�3���2�Y3��^3��3I��2��13X�L3�"3�>�2bZ3p�2�K3o�2�3h�U3H#m3�O�3�>3޹`3{p�3�[@3��53v}:3�)3���2؁�2��3���2s�3��3��k3��(3���2�F3�T�3n03"3�)3z}3���2��^3B�3���2�pI3�>�3"+83�d�2}��2�<83��2=��2ba38�2��3�β2�A3K!�2-�f3w�
3�o�3�Q�2�9%3�
*3�M)3u�2�j3Y�\3�*�2Y�23uq�3՝�3�73���2+�3�:3��2=K3���2ɠ�3�3��A3�3*�2�l�2���3�2$�3�CS3b$3+g)3�|<3��=35��2K?^3z0/3��e3�qT3��2�643V)33D&3+�!3N�2��3��2�Pb3�gP3C�3E^_3�[�3W�	3G�F36�=3FW�3��-3�Ǟ35�035Z3vAy3�z�3���3,)�3
�E3,ئ3a�A3��3S�D3��[3m��3΄3Ye�3A�53���3�~63�3�333�v3=��3��Y3g�93���3��q3.�j3� �3�Ғ3w�3��3�V3�H�3��G3K$T3�!B3��)3'fy3�t�3��3�ź3l}3��,3ꗟ3�QC3�~3� 3i13�!535��3��3c�!3ف�3x�4v3�13�/3���3*�w3p3�z�3�f3ַ�3�]�2���3��3�3�V�3��3y�B3��53N�N3�3�W�3�� 3��z3B�63�1�3>��3�3@t�3;J	3���3ēe3�#3�E+3,B|3��l3E3��3j�3��83��P3�14��3�q33O�3�+I3��3��3�~D3�93Y4�Kl3�co3_ 3V!4�-�3Ev3.Mg3�N33͘*3_&31�3�Z�3�3�Cd3n��36<�2�3��r3��;3or�3]d]3J|�3�1-3��3�S4ܗ�3�63N 3>��3P��3�,H3�L�3a3SF�3��d3��3��:3VD3H�)3Ut4�ԁ3��Z3���3Kw~3D3N3��N3�d3fӕ3��@3��3σ3=��2]-3�^�3Xc	3:�]3D�D3��u3<5�3�1�3&KH3t�3^�o3�.�3�&73`$A3C!3b�i3i�3n+`3\{�3��3�+V37X�3\��3��i3n&3��3��3#��2�:q3�53�v$3(�=3É�3L�[3@uD3ݟM3��4K�n3%HZ3��3c8�3zS3U�3	�3�)3���3���3T�33��3o�N3�p3$��3��B3���3�*>3���3�=D3_ٚ3ۢa3�$>3\��2j��3oe3Z	�3��{3��*3C��3��P3�n�3�:3��:3>�3�Ǥ3u13��2�y3�s3���2��3���2��3�{H3	l�3��.3\�3�3���3�<3���3��Y3���3��?3L9�3T[3��30s-3K��3)+z3`��39�a3���3�wL3���2��V3��_3��3�$"3���3�N�3+^3p=�2���3�g�2\L3�\3^�]3N�73\�3`�3<�P3��j3��3q3�3{��2���343�3��#3�^�3Z�'3a>F3B�O3]�R3��;3�^�3
��2R5�3��.3�3�13�=3X`I3!�E3�=�3���2��3q2�3H�3��J3�3�Z�3���3v�3(�W3���3�ߊ3À3\�Y3��f3�l3��J3�A4t�3SH�3n�Z3A;�3ve�3©R3���3��3��;3�l�3��3Cq&3�<3bh3��~3j$P3���3�0,3`h3�t73낫3�{-3m�h3�/3��4dQ3�5H3h�93+�Z3��	3��_3r��3i�3�gn3'�3��3<�3��>3ܟ3=�x3	1 3�e3c�93�uZ3�J13��3��V3��3R��2ZB4��.3rk3���3t3C03z��3�_3W�3�,�3,(	4⡋3q*3���2l�3�dn3M�3�/�3�"�2�ӓ3S3�{�3c\@3=�31�3�q3r�S3y'3��h3�
�3�+o3v�3�_3��@3(AJ3$�3�G3m�>3-83d&3��03��3�L�36L3.��3 3Q�3�j�3�13>k�3��4�Fn3�_�3�aA3���3��2w��3�֞3��3�f3I �3zه34¹3��3�9]3쒰3�$13H23�E3�W]3�j3#��3��03X�3�eL3��3�`3_��3��.3Df3T�|3u�-3�-_3C4P3��3���3�5�3J�{3ʓF3a�3i7�30�{3�=3ߓ�2�ea3U�v3uF�3���3"�3/�3ߵ3��O3+�3JX�3���3��f3�m!3�.3�!3� �3냆3I,�3i�3�y3���3�,�3��@3h%^3�3��J3u5.33(�3Mλ3�E[3W&�3)�z33�[�3B�?3a�b3��3�I3��<3�+83��-3p�3�9�3Pz.3I��2筇3,SG33��2-�`3y�83�}3,3�38WK3f�[3��2o{�3�̖3�F3,�@3�v3D}E3�AH34�_3+3QU3R�3�@�3N�3v�13��s3^PU3��73hNM3�u3���3+3\�L3��3�΄3�3�m|3�z�2OT3��63A�~3���2�B3Ḧ3,�2�=f3S��3�{�3�0�3�k�2)o3"uk3�T�2��R3��L3㉈3���2�}s3�� 3�t 3�+�2�Q	4��%3��2Z913�p3Z3��3�qN3�ɴ2 ��3���3M�-3#/-3k{�2�Ec3V�03�W�2�{V3�:3��l3X��2�u�33O"3Q$3�-33!!�3�-3	�U3C[3�M3ɔ63�o�3o�=3�3�2��B3ֻ�3���3�n3l�V3���3+z3���2���3̗03pD3��3PG�3,�2�K3/	3-,�3
1N3,�B3�*3nnC3 R3O�$3�m�3�|�2#
y3A��3 YY3!�K3Чg3Y�303/~"3���3Bq:3�gE3B�2�o�3{�73�Q.3���2���3X3���3�GR3��3*353a3e�3bp03prb3�1�3=E3�� 3&� 3�S3��@3�W3[PM3�C3��3GD�2*�3�;3jC�2��3���3�3B�t3#�!3
�D3�3`b43�~g35�53*+3(s3rc3��`3Mh�2}�\3�N3@�2V3�� 3=�E3oE3>x~3R��3��+3�!53us4��]3";33�V3p3�*3��3��>3���2�o!34�3���3��u3o4%3 �V3]Y3ў)3�3���2j�2׿.3z�u3�#�2Z(03�3ft~3�<�2k�Q3*a�2Q�?3��2��2ől3q!�2J0n3�ڴ3��3��@3���3p�?3~�u3r	�2_~3&�)3k~`3���2���3�o�39��3��3KD�3c��3Ĵ�3��K3SǊ3���2;�3�̃3O�3{3�� 4H��3��3�`3���3�`�3��J3xt�3��.3���3aB3�A�3�=�3s��3�X�3���3$�3���3�\3/�3�d3`H�3Cк3�:3?_3M��3���3w�93�03H�k3L�L3惩3C��3Pm�3��3�[�3���3C��3C�r3�3i_�3w�H3�{�3�)3��3c�53RMQ3��3�8-3�5�3���3}�3��3s'3���3�\-3��3��y3��;3��3�.3_�4Wzz3g�3�	�3�6	4��v3�}3�,�3��I3�܀3�_a3ǃ�3-Y3��3Wx�3��3Zk03�043+B�3��13��!3�f�3��E3�w�3�J^3�[�3�4E3�Ii3��03�]�3�r3^�3+�u3�8D3�f�3Z\3�%u39�V32��32,4�
h3k�{3�C3�K�3V[�31A3���3:�3]��3.V3�4yޚ3��:3xSR3"4�e3\(73��3�h�36i83S�F3�E�3��3�.Y36�j4ϲ�3��y3f��3N��3�g�3���2i{�3n�c3�3(��3�	�3�=3E֬3�	e3<��3���3�=l3�3g��3�s3���38<�3�p�3��3M4:��3�ѓ35D3�J�3fB�3��3��v3�3���3pT34^3OÇ3��O3�{@4�;h3m|32c3��a3X�b3(\3l.�3�5Q3�D�3$�94���3��N3��3��3�T�3��u3�+�3� 
3ğ�3�k3���3W"3[��3�Ʊ3��4�}�3�F�3�v�3�3Lqw3���3��:3��a3��3�y�3���3Y��3oI3�M�3�r 48��3�ج3W�w3AЕ3�|K3��3���3��{3��*3��3 n�3"��3��3���3�~�3jf)3^��3��3e�q3���3�tF3��n3��:3�2�3(�|3wI3Q��3(ă3})3�;)3}S�3S��3��3��F3+Y�3/�[3vX3�:3}�[3`�3z��3�N3-R3��_3���3��}3q)�3��3m�G3�73/L�2�?e3�^�3�y]3�t�2O�3n��3�J3�73��3�`	3҂V3*�k3�.�38�*3��&3��K3LD3�@(3�Ƣ3�D]3�_3�2	�3cf3�3�Q3��43�Kk3��2>�3a0/3n�3��43A9�3})3�x�3�q�3�Sm33i�2�j3֛F3�M<3��%3���3=�3�3�$3-�w3�p3���2;��3��"3$��3}�O3��M3L�E3̕M3_Ă3��3�$�2s�3{�3x�{3pv3�OQ3�5�3x��2Hx�3�I�3'��3�=%3�P�2tVj3-U�3a 3�B3�H�2�	�3оa3�)�3IXl3S�3C3�04�8[3\�3��y3�\3F3OΏ3��_3H�3��E3���3��3e�3z�2z�C3���3�h�2�B�3=�R3'CM3�3�g�3]�n3��%3�:3ZY�3�� 3Mfa3��3���3M�3��e3	M�3-<3GtO3��3=��3��'3���2���3@��3e�K3OC�37�2{R�3{�U3��b3Mφ3}�H3�3X3;X4�3��\3��3t}[3�,3R�N3�x3��3��3�ʂ3#��3�-3�3�m�3�D33�3��s30%�2��3�3�˂3PkC3���2���3$��3��Q3ÐM3l`3�A3��z3�h+3?�3-�r3�E3�c�3IA�3�SZ3��3���3�3��3
�3�	3\��3�2�,�3�X�3O�"3�Z3�H�3BQ�3Ƨ=3��`3�F�3*G3��3��b35�3�	�3[� 4֮3�bQ3�3��s3�x�3G3�2O3�hX3�J31	3hȹ3oc3l3�83���3�YL3�%�3�)D3=��3̳3��M3��o3C��2/�3���31r�3+��3�3��3p�B3{3_�`39�2��j3$_3�u{3H)@3�>3x63�'r3Ҩ83�z3��D3.=)3�d3���3��N3k�R3���2��m3fc93&�L3��2�L�3���3uX3��13��3mo�3g�3Z�=3��]3z��3)�3S"�3�FF3���2%�}3���3`�3M3t\M3)�2<M3ؓ�3"��3*�?3I�2U�3�^3��2��j3��?3!%�3���2�N3kjs3y=v3�}*3��3�Y*3��q3�x&3��R3�r3�.C3�[93��;3�+3��3��I3&3���2��3��e3�Cv2�/Z3�b3�T3�1�2���3l<;3�)$3��3�7�3�3�^3i,3C\X3)LA3%�3%[u3��2�� 3��3y�3��?3��2#�]3�@g3t��2Ēv3Ѥ!3�7�2n@3ƅ3f�3o 3^�2Ɣ3o�-3�j3 �a3��3J�3Yƥ3m�3
 �2P�V3��3�V;3�L'3Ff{2י�3It:3�\�2,N3]�3~�,3 �63��3f�?3�83"�3`�]3#>�2C�y3:�3H�
3�y3k�}3Gu~3x_3�m3ȁ�3C��3>��2��	3b>3Q,�3,M3�63. E3�]3��g3��3ǟB3���2?"�2�r�3ū73�63c�3�&3�%39id3�F3��(3��13��3�Ѯ34�(3ۄ3ȿ>3
`3`�"3��S3��3�Ke3^�M3�g3��32 3m�3�ǌ3��n3�YK3MF%3��]3T! 3�lc3fД3a�+3��_3���3>�3�&3F83�q�3CK�3�3$
�3��B3h�@3�3�-\3���3I�43UB3|��3�k3�3�mJ31T3��2b�i3}�Z3��
3\�|3e7�3x�Q3��3?3EA03��3�k83_Q3~L>3�n[3�}3�%;3�13�,3��2?5 4��3)S3?�$3�Z53=3��l3�^3-V�2��83@��3rߜ3�9P3��+3>t3�d=3�3C�39 3�%g3�k3j�3u3��3�_~3_<�3�83�3�3�ݓ3Fl�3�?3�p3]#�3j7�3�d3u��3�9�3�d�3uއ3�K�3;�f3�3("�3^c3�J3��03δq3d�3��;3��~3�4�?3/ 93臥3�l�3%��3U&�3ѱ3:_.3�7a3k�3��3�`b3�423�9x3Ԇ�3�83�.�3��2�^�3�e3��4��N3E�e3�#p3�"(4j�X3�X 3ɏ/3=��3�"[3ѓ�3�=�3L@L3�Rm3��3Z�34�23S 3�h�3đ�3P�k3���3�n�3��3ꅫ3�o�3�:3(<�3c�U3��K4"r3�C3��]3C�Z3��[3�/A3Υ�3�>3:�3�i�3�*�3OY3a(3��n3�ܦ3���2<��3�!I3jz�3Z�>3Yl3fwR3�\3�ڷ3A4��{3(ۛ3�Ε3��3J*t3��3��j3+�3�Ey3=	�3��3��3)M�3ݽ�3��3��E3��39�3ʮ�3��,3�3�o�3g'�30q�3��4Gz�3�a�3��i3�,`3���3l�^37i�3H�3�j�3p�3�1�3�=�3�3=�4�K�3
y�3[ɕ3�43�BG3��3,ȇ3��73��<3:�>3g^43#r3wσ3U�?3䇆3��3���3�L�3���3���3؎�3���3 �c3Z�%3є4��w3��b3
v�3��3Y��3��3�6�3<{�3^8�3]�@3n�3=��3K3�3�+�3=$.3Qw�3"�3@�3�8�3���3��4�ֳ3���3��13�d�3�v3���3�F�3ejy3���3�B3��	4J��3T� 3
2d3�+4fF�3]_�3f��3h�3@g�3�.{3�̐3��Z3�L�3���3p
&4�e�3��2Qj3���30�o3�vF3N$=3��3g�u3`bm3s~�3C�.3oYp3�]4��3���3��{3��@3b]03Dc�3�q3�3�g�3ܒ3�K�3r:�3�B3k~�3罔3w�3A�3{�3��3�Y�3��
4���3t�U3\�2�T3O�3�P3�Y3?Q.3�7 3��2%$3B-W3�:3���3��<3��3��_3��36h�33�I3�yv3�N[3��W3�ʀ3�;3�U 3��q3��@3]�3�]U3*��2��?3��:3�~]3��l3m�r3p�139]%3�.v3*P3��2��3�uG3[�3�:+3�AK3(�/34�3ל�3���3o-3͋3t�3Co3YFv3�J3� �3��3�+t3�m3P��2��/30s�3!K�3��J3�{03�F3�33-I�2��-34N�2^��3?	'3��V3�|>3�+p3c� 3�C�32$3k��2m|3�3�2r�;3h�3�3�2g�M3��3I�x3G�3���2��43f3<'�2��3�>-3��3"�53�V|3qY3Y35l3��3�
3�
33<�3U� 3�h�3j�C3�t�2NlV3�i�3�'3C3���2 ��3a��2�W�2��O3uM3�oO3w
;3��]3ΰ3!G3i&3+�3�f-3*
$3S�.3��K3.�P3�M3	HE3� 3\��3T��3I�E3v%O3i�3��]3/�:3�
�2��L3�Q3T=`3L�%3	�30�c3�23X73��3xb3¢e3�M3��2��3�13
W<3��2��}3�
c3�_3�{i3g�2��3O^3���2�C3J��2�	3>3��}3��/3w�3�7%3���3�b�2 \3��3�wd3���2��(3'nQ3��2�g3l$�3���3R�P3�Q+35��3Ӡ3�k�2#?3�,�2�A�3R3>bv3A>63�)3��*3�ˮ3 3j�.3�~3�3��27�J3�ha3�\�2hY�2C�3��3	�G3���2\�3W��3�3~v�3h y3O]3X�3��r3��D3*m�2"�(3��!4���2�'3��>3"1#3�n3�i3�(3>��2�%�3�ʒ3��3��43I7�2�im3�'3m~�2,��3���2�dW38/*3��3z�3Ț�3�u�39�4�d3�U 4��<3�F�3�O�3RJ�3�ُ3"�`3��o3H}�3V�3���3�63���3	 �3���36�o3�(�3���3 X32��3��u3�J�3R��3��4U��3&Y�3p �3UZ�3'I�3.�3hّ3�M�3���3���3��3B�3M�23��3,�3�l3{�]3�V3?M�3��v3�r�3Xǐ3n3�3Q�<3]�W4�W�2�KH3@��3���3.�93H�3�t�3�?�26E�36�3PƋ3�I�3�NA3���30e�3�3���31�33(W�3'J�3E�4]֖3q��3i��3o�4�0\3pT�3N�3ϡ37��3��3m�3d�39��3�54^��3'��3��f3#B+3�	�3wz03�z�3p�"3EE4RUg3��3�Uz3��l3�:e3e�42�@3<u�3ђ�3:�3�X3|M�3F��3l�Y3iE�3��>4ƞ�3��:3�'3dt�3^َ3�a�3���3o��3%��3��[3�F�3��3��A3H]v3w?4r%�3v��3'�%3�5-3��F35L�3�	[3�.3��3�@M33�3,D�3k;3�&+4���3Z '3!�43�_83�6�3�3 �3��3x&�3�@�2�TM4>">3'�=3�u3�A�3(��3b]�3��3��N3���3�s�3���3�0R3���3�3�h3�23;�3�@d3Ǩ3���3��4�3��3���3{iR4�ĭ3`V�3"��3Q	�3��3`�3���3q�3�8=3�tS4�}�3���3:�j3���3�4��73�$(4\��3N4�3��S3��3��:3a�A31��3X�s4�s3��3�3Xf�3���3�y3�ݱ35�L3!:y3{��3�3ϊ�3�|3�m�3F��3���39��3�3��3�l	3T@�3�K03�P3Ex)3?�4�jO3N��3W��3�t63%Q3���3,��3�a3k��3
[�3��	4*��3�`3���3�/3 �3�64n�|3�4�a�3=4��3U�_3}]]3\{�3D3=�Y3�3"�t34H>3�V�3��3^�I3K�R3�B�3T�_3���3-4 3�w�3���3f��2��$3Q O3�9�3�;3� �3)H�3W~u3��3�3&^3n@3�`.3��r3�3Ⱥu3L̇3�a43���2'�P3��L3`щ3��3%043a�z3��3�D3�nF3��3�}73�3�(w3i�<3�03r��3��3�j�3�u�3,�^3e1�2rp73@ȃ3�J37�3=մ3x]i3Kx]3w��2��'3���3��	3^�_3���2�3�q3�I�3��3Tχ3�m3���3dC3�63�aH3;r3`�2� 3!~m3&��2~�3B>�3;�'3613t��2��73��38��2U�W3�'3:�{3)�'3���3�s30Gh3�b�39��3K�3�I=3F�)3��I3*,3���3a��3��3�,j3�z�3���3�E�3���2���3��b34��2-T�3�dD3+��3�F3I�}3��33�R3�S.3M0�3�B3T��3;�3F�3�ST3��G31͖3n�`3�&32��3�ǔ3~Ql3�9�2Ï�3��`3�3#�N3�9f3�M�3�*3Df�3c�}3��<3���2�I�3��o3ڣ33eƘ3�$3�Qt3x�%3��o3}�3�I'3ma�3Kd�3=�3aw3q��3zn3AɁ3��3���2/�%3��23l��3q�3[63�o3���3�
p3�\O3�X3�$3&�3�G$3c3w��2�O�3O\�3SG3|�3193��33WG�3N�_3jV�3�Q�3p�!3��@3Q��3�^3�^63��3�;�3�&3�h�3��Z3�f63��&3�_"3H4�0^3j�83��3��3Y�i3�&S31A�3�38�3��v3�(3_�3�..3{��3aEE3h�2��2L;4��.3�Uc3�3W�3�13�G]3��y3�O�26�,3=�3�7�3EjX3Y�3`o3��g33i�2Q��3��2ݴD3X�53�0�3.�"3��/3Ȱ|3� �3�3R�<3�/3V3�2��32|�2	3F�3K+�3�|\3s�m3�r�2f�3<13���2#s!3`�"3�733���2v��3�I3��3&�2�!I3ɋ�2|�A3u�93�*>3�vH3�/3Mnm3xv�2=}53�a3+-3s��2��2VFs3�3ї�2�h3�h�2>b�2Ǚ�2��@3�{A3��O3"03�	�3D^%3�3�,@3�n�2Y��2�-]3~g3��3Zs\3�c�3ϽR3��2��2v�(3�h3�f�2�_ 3��!3p�'3 )3��,3�/�2��X3���2���3�'�2�`�2�$#3j3��73L|63@S&39S�21�E3̎�3\��2[3ΰ�2��53,(37	 3�3�PN3�$3��2��3�	3�3���2!�3�3X��2��3�2i	34�3� �2��2��B3Y-3�7t3��53�Y3�D3���30�/37�2�#37�Q3���2z��3�6l3��2޷3${�3̚3�A%3X^�2�q�2��3@?N3n�/3�;�2l�3��Y3��N3��3�3��3L�X3�>3y 3�k
3��Z3�4�2g}3n�03��53��$3��3�53sA3��2ɮ 3�:3��"3�&@3N�3��28V�3oK3�3�3Ԟw3fF&3E'3ֆ3m�2n��2oH,3���3_��2��'3e��2��T3��3���3��$3^�)3 ��2�J3Mev3[3Y3�(�3��S3a�63st�2lo3>3@�3�M3-�2�i-3���2XxB3�D�2�^�2F�F3t4�s3/�I3��N3$+�2�-3?R
3�=H3�*3��3��53�,i3��:3['3/wS3h�3��+3(�3��3�Au3���2t%z3z 3�q�2�3è�3�3y�^3+��3It 3�3��@3)-3�
�2.ڃ3��3��3'\3�e�2�93�2�39q3!(^3�\�2���3��73�<3�g3���3���3A��3(S�3�A�3Q�3���3G�+32b�3�RZ3�~M3�ް3��3>��3�]�3YX3�g�3�:�3ᖃ3.-!3�t�3r�q3g�o3B��3H�3�5^3��<3��	4l��3o�3��3�u�3�C3D�3P�3}�3s6�3|��3�:�3M��3&3G�r3���3��3*F3�-�3��N33���3[u�3}n�3F�3��,4�H�3 fI3�]Y3���3,$�3�i�394�3j�)3�n�3��4���3uF�3��U3n��38��3A��2q��3���3�p�3�ߟ3 >�3�}3H �3d�<3��4�^3�ψ35��3-�*3K3>��3]>�3{7L3��3��K4�@�3Y:�3.҆3���3�	3`-33L�n3���3�X3
V�3�Z"3�+�3/.:3%��36��3ߵ/3�?3<�3SՊ3K��3�F�3?{3��I3��4���3qgm3b:3���3��4Z�[3��3iB]3b/o3��B3q(o3��u3�3��3F�4'S3X��3���3㙠3u�m3��a3_�3��"3aD�3K��33�3!�Z3��3,J�3`�|3B9�3w�s3���2��3�$s3q#�3'2g3`��3&�2|��3�N3���3�l3Z@�3Uo�3���3CG�3��.3�o3�4P��3z8V3Sq3�=�3��33M�X3���3ݔ&3<��3"Q3D��3�xD3��p3�z}3�4��3�!�3��K3�N3�73�p>3���3�]3H?�3�-(4�Τ3ޚ�3tZ3E3C�3x3&3���3�B�3
�3��O37�3�+3�933�Y3�5J4v�3gh�3qޣ3�up3*�3E��3g��3��33r��3�Q�3HG�3�¹3c�3ۯ3&D�3��93��3��3���3U��3G(�3�s3��?3D863��4'3;��3��3=6@3�Q3}�3I�4؋(3Ik�3(�^3�H�3���3���2�m�3�Ӎ3�]t3T/�3R�3�4�G�3��x3:��3n�3��2dKU3�Z&3�e�2��3�$3�R�2�u3��3��w2\�	3�!c3V�3�"O3�2v�.3wt,3���2��(33Y3�83T��2|��3e�#3���2�9(3�'�3��2��2��.3��2���2B�=3��3��3�l�2ϑd3�3ۢ'3;+3M	3�3�I�2$�z3��3>��2	((3�43�3g83���2�!�3+ 3��2�q�2QxS3%�j2�2g3��;3�K�2D��2ln�3��2a��2�3�2�z3j�3�1�2�+3�\M2��2��3s13�� 3���2��3>��3ޔ�2n�2q�\3*a�2�:	3��2^g@3��2��
3>�v3�Q3�6�2]nW2�63�63vl�2�_3���2�'3F��2ҧ[3�_�2�މ2X�'3�3��2At�2x-3�0,3��2�53�g3s4�2�3��@3f�?3p��2l�c2z�n3y@32e�2sR�2�(�2��3V��2z�.3pȮ2,�3y�2㻮3�*�2�K39G�2w�3���2��
3P^3���2���2*h�2��)3�~.3�`�2x�3�53���2��2<u�2�3e�2>Q3-��2��
3	�2���3S>�2�3��3���2{g3�F3M�3x��2��3>s!3!C3�-83�w�2�t3J�3�3w�3�˺2ċ53�3�L3���2��2�x�2�3��2���2C�3�x�2�A�2)3�3�y�2�?	3l3�34H3��2T�	3��!3	�23
�2�03���2�vB3՛�2���2��*39��3S}3��%3�D,3h��2K�3�$63M��2=��2�]37�3�C3��3���2P��2�n 3�3���2%V�2�a/3�3��f3g�2��2!��2���3-��2t�2@4=3�{34�2�Z@2U3�)w2s.3�k.3Ȣ�3(�3N?A2�F^3��@3*�2���2 +�2�P�2�Ɉ2�&C3��3�I73�z3�}�3��3� �3�_�3�&k3D&w3qB�3rw3{�53��3CI�3�X�3~�3��&3c;�3h<�3��f3�4b3���3��`3n�.3!-�3׵�3N��3�у3��4 U3#�v3�̊3⟜3�o
3EƇ3,��33m�3�'E3�o�3%��3���3�a$3�N�3r��3�3�ݔ3�b53��3R�n3�Θ31�w3M0�3+��3�zS4\˂3I��33f�3��3"8�30�=3�3�B3�J�3� �3�Y4m�!3��2=3Ym�3��#3�i83�:3���3�TO3���3��!3s��3 �A3�G4K*}3=O�3�m�3�r3Mϗ3ǁ3��3�)�2�©3D 4��4���3��3���3T�3��$3�Jh3�=X3h��3+u
3�`�3A��3;�3S5"37�4u�I3��3���33�I3|;|3��3�D�3��3��3S�4��3lWS3o��2'��3���3\Be3�	�3�d�3�JI3��o3���3�EJ3%e�3�(U3���3�XB3�X�3
��3�n�3DZ3��3��3
	e3�N�3K-4���3᱓3�G3應3S��3�Y36�3_j3J��3�El3\v�3T��3ϣ3�z 3�$�3j��3��39G3��3GUd3�3\�^3��3XX[3��4ǭ�3qZF3?P'3�u�3%�3�N3�~�3�e�3PT�31�3���3�g'3���3Ѣ<3��3xh�2��~31�83�տ3ֺG3Yڿ3Q��3�E>3=��3bI�3+U�3+j�30435��38�{3�3'G�3�\3ST�3�UT3���3u�v3��/3��A3��3��3�7�3k��3��W3�Il3L��3�ξ3}*3���3���3���3���3.D3-^3V��3�L3(��3�3��4�(3��P3��3�C,3@�3�&44"�53�H�3;3�=B3h$\3�i63�ch3W��3?6�3g|p3��3O��3�j13��3J�Y3�M3�_�3��X3�[o3罠3��3��v3|�3�i%3p��2L�R3��3�K�36�3 �@3��<3��a3�Y�3��2�3�3�=Y3s`O3,.3+�B3m�$3�3��2�a3�sI3�Q53�2}3@�2�f<3��C3BՐ3���2��w3�V3YUp3^�33cU3�a3�I3^�g33ٰ3���3�u3"��2w�y3���3�;�2-��3�m
3�GQ3��2�e`3��3{W�3�7�2�s�3ޘ$3�d�3̀�3�!3$/3�9V3���3
b�2�%�3�T�3��3 3!=�2�_3�PR3}��2	�633N/J3I� 3>�3i�3�_�2��3�4��+3 oR3f� 3��23�J�3�mu3��E3�c�2++3{%�3���3��{3�3��3?��3>/3Lj�3c�G3
=53�x3�FV3<f\3	H3��3]��3�3���3-�Q3}�+3��3[�3�I3o#3zN3�Q3폹3�X3���2�:3D�.3!i3��C3�_3ˑ�3ce�3��.3�J�3���3��2��4R�2w�3=��3`3��2�]<3c�O3�o�2?T3�{�3�'3
%�3S�Q3�!3��b3�Ϟ2�3<3+u"3Gj63C�/3W��3��3�p3�3>��3S�3���3�)3K�*3T�:3�<<3�u3�v
3r{i3c4���3�3v��2�je3w�)32�3zQ63r�3)k�3)9�2���3I�Q3n�2��$3S��3s�13�3��N3�X3��-3 '�3��%3s]�2�#3��3�/�3�z3�>�2�SF3��63�lF3�,�3�k3A(/3�P{3ݨ�3��3�?43ޤ�31�3�3�+n3�T3P3g�_3tI3��3f��2&I'3��a3^%3��53�K�2��@3+��3P��3�ǈ3>��2�d�33�3!�3�d'3�&3-و3_��27�3��2�9.3�C 3�3�$�3j��2�*�3\$�3�RZ3a�,3Q��2sO3[�3t 3� }3P�23v�36��2�!�3`ZH3���3V��2���3��25�Q3���2yz3v��2��63�3�2G�3�?>3ư�3�kD3&rr3��2^�a3b03F(h2�m3p��2c�3��2���3�]3�#3?��2ک�3�3<�k3��3hj63lMk3֦3VB3َ03��>3�:�3�3E�2���2�3�lb3��2� 3��3��3�3g��3?x�2/q 3�M3�k�3��2�g3[�G3�}03�/�2�
$3��z3a�2�h3��31��3N3tn�2$�3	��2��2<�3���2u�|3��3?"3�.%3�#y3-H3Y+�3Ww�2�5P3��3�w3���2�?3�3R��2z~3 
�3[�p3��13�E�2�3M�P3_H�2X3�q3��3k1�2`�33C��2y9�2) 3煄3a�3�23Z��2z�3B��2wi�2�w3� �2���2c�`3��a3�&�2N�2�3�73ư3;�T3�p'3�E/3���2d��3�bz3{�3Oh�2R۽3��53H['3��3q��2�K�2
x3U�32X�2T�R3�	�3x%'3R�2���2��i3.\F3�w3l�$3}�3�y3��2O�c3]�*3s��2vH�2Ӗ�3�9�2��3��2�3]�3=8�2�13/�73�d3So�3.�3(3��2pX3��2��2l_%3�%3B3�L3�Ct3�J3�3��2���3�(^34�33`�F3'�3��3(S3�E38�2�|k3)V3� U3���2H��2��=3�|�2 �2�*_3�B�2��S3 ��2R��3�T�25�2G �2ڜ�3Q3�3%��23�2�۴2�34f3Ӄ�2g�Q3��33� �2���2%&83o h3S��2���3|Y3�'3���2݀�3�� 3&��2s��2�q43�3S3�t3��3�k=3o�3[0�2��2W�3�G3���3@V$3N"�2×3�� 3���2��^3z��2�3N3  3r.3�93��3��3X�3�E<3\:3/D3�f3TO�2#݇3��?3)�3�Z3��3Բa3��3#xW3f��3L�3�!�2��3��m3�XS3�O�2i��3��3LQ'3�[g3\��3gI3�|$3b�f3�Ve3>�3==�3c3�33͑�3���3Q[�3ټ43o'3���3d'k3�'l36�3�E3�h"3^�<3�C4)'G3<ig3��>3�Z4_O3��C3l˔3V�3��c3Z�-3ɵ�3��b3�M3�Ă3�r�3��d3��*32]3n�3�t 3 �a3��D3��Y3Xt3��3�*3S;E3�03��84e�2�hs3#�3��+3�-3�vL3�ܽ3��E3�1�3~ӻ3~Յ3�9 3�c�2(�)3���3���2RX�3"3Z!�3Jb3�>�3A$3"E@3�/3:4�!i3d�03�[3f(3�%3,m�3,��3�!3 +g3 =�3��Q3Im^3���2�w�3'Oh3Õ=3t�3.�2�ې3*�3�1�3�-33~�l3T�B3��3��q3�~3�c39F3{�^3"cS3�%�3G3�9!35B�3�3l4o3-�=3P�3�%�3�$3-�R3E 3�fg3z�32��3��_3�f43	T3)�3�[3�"3�3�3�"G3K��3~^w3��U3�!836m�3�	�3�x3���2�3愅3�F�2�@F3�!3�:3�"=3L��3�g53��3��3�6�3��%3�{3��F3���2�3��3�`�3}#3A�3�Ӳ3SlW3N��3�C�2�I3��3��53�&>3��>3]�v3�Ђ3�j�3*�*31��3�&3M��3�>K3l£3��3Ԑ�2!�<3oɒ3��m3+3�_r3�~�3,�`3.+�3 �D3��3g��3 �.3^�I3�k3���3��:3E�3@�;3��
3�13��4��3GT3�g3_.3(�2���2 43<� 3���3k��3+�34�3A�2�^z3�P3 �3Tr�3ʜI3!!�3d�?3��3���3���3�v�2�؎3��2�b3 �N3�c3ϫ-3��3KG�3��N3.�3��3���3��L3�b�2o��33�3N��3�I@3���3e| 3�@�3I�{3�s3���3��3��P3�=�3V��3b�j3�gw3ͫ3إi38wE3��3�І3�1|3�m�3Q��2�GI3˼p3Qy3&�E3<�3�G�3�23H��3ٟV3�1S3��2D��3�S.3�I3^�:3�#43�3`�93Bc�3\A3I�t3Gɺ3��d3�;�3�ɧ2���3�x�3�93%9>33f��3Sm3Tf�3vr37�3G�T3&��3@�3!�#3�l3�u|3cq�2��3��3Ī�2�҃3K��3j�t3`�U3�,%3�^3�T%3@D3o�k3�3��[3�}3�p3���3��
3��83��3�RN3g�i3F3�ew3��3�o3�A3q��2�_3,��3�z�3OB3���2��3�e3.�3�N�3��2y-/3�I3���3K�	3o�m3 �3���3�-3ޔ43�}s3���3�M3�P;3ja3��%3��Z3���3�vZ3*�2��3+w�2�3�{B3�/C3�3��63�[�2_@G3��3"�03N��2�g4F�I3�_+31�J3<Y3��J3�&3�d-3�{�2.#3Hm�3��3��3!׋2`�[3�53k�(3�i3�w�2�!@3��73X?�3�YL3�b+3wjR3��3o�W3*w3�3�sJ3��3|�C3NM�3˗%3
m3��3�S3�fV3��P3�CN3���3��2���3:'3yH63ӵB3���35  3d�2���25�4�{|3��J3��b375�2PQ3��3ZS3�0�2h�&3���3�y3��3���2%
�3j�K3*��2���3� �2Ԅi3z�3!e3�	&3X�3�k�2|B�3�6�2r�2��3��3mo�2��(3�>K3g �2��3��e3%y�3�n(3�3'�W3�43Q��2U��3C��2�x3R� 3Y̿3�i�27d�3��3�ͽ3��X3�{3�3��3
R3/��3{ȗ3w�Q3�[k3�s4�ϝ3���3VV3���3�63b�2�X�2�~Z3�^�3��3���3��3v��3r13	�4�h�3Y��3#`13K3�;3{LU3Mˌ31@i3gm�3"�3�j3�o3�3ֵ3ƘU3�` 3P�3u�[3��138#3���31�f36�3[�	36� 4бS3/3�GR3S��3�3�+h3o��3�� 3G�L3�c�3��3��3�<3��"3���3�>37�h3@h?3��3 Y3��3]��3�*T3�PI3i@4��w3m5s3J�3\<43h�!3�,_3�3�93E�3�Y�3Ϥ�3|�s3�ɷ2d^�3�a3��3B@F3��M3���3j�3�C�3|_3HcE3��k3�#�3I�:3[ѓ3@�3��E3�0\3�3�o3��@3�yM3���3��c3W�3�@3n�3���3�n3�|3*�3
h3��\3���3؛�3�dT3�N3$��3닇3;0�3��03��3;F*3V��3C]�3!@�2kjc3Ƒ�3��3��3.�2�3t^3&�3�3�mD3n��3�Ʉ3y2l3�W3��53s�#3\
4��Q3��83˼F35��3Kx3C4���3��3��C3���3���3��b3�'�3~�R3�7F3��3,�3�u3�173৅3��3h�L3��3�>/3-~;45�N3&��3-#3*;3ı�3BY3�G3�l�3NCo3��3��3�'Q3^�2YL�3~��3��2�53ǃ3�VM3I[|3���3�>3��J3Ԋ3��4t�b3+�b30[3a4�'63�3��3�,�2��3��3Y��3l�^3��)37�D3
Į3��w3��3e�3F��33�3y��3AW3T[�2��3X�"4�*3{��3�3�3&�3L�2�|u3�ur3u1�2:6�3� �3r`�3���3~�3�]03˨�3K#3�	K3/�24��3�3�h�3���3��33�3��4���3��3f��3)'4ȯ3���3�8�3@�K3�3��"4�3�f�3�3�32�34�i3�?3w]�3�TL3�w3�$F3�3]��3䯆3�R�3�4��13;x�3�V3�3��T3���3��3��p3�7�3�Ҕ38]4�.�3�,3e��3�L�3d� 3	z�3G�3ź�3�b�3\��3W]�3�d�3�63��f4��v3��3_��3|²3�>13N�3�3:�A3�ώ3�e4^��3�p3�(3 ��3&��3� 3��W33aC3�U4�(31�3�*3�42g3�>4Hr�3S��3ɝ�3$N{3���3� �3ݦ�3��F3���3�4x��3u��3V�?3���3'o13��3%2�3*-3�/�3D��3��3Z9�3��u3�
�3�z64v~3�K3*�3u��3�{3���3�ç3�X%3c��3724�6�3�qi3�H.3���3ʥ�3
bJ3>��3�r3��j3�.w3�k�3p�3��3�2&3�\4sRl3�M3�wy3�q�3BC�3���3Ď3-%v3�8�3�#4N��3��3�@3Υ�3'��3`�3*v3�ƛ3Z4�G�3���3�Qf3}r�3/3j64��3�ι3\̍3WBe3 �3�=�3�ל3��}3T��3�Q4%�4��|373��3+��3�I�3�ƪ3aG3��3�~�3j��3kA3���3N�3��4�x3RR�3'��3j��3��&3J�3j��3��3��[3�K)4[��3Ͻ�3r2h3�U�3ӱ�3P>)3�e�3�p�3LA3��@3�X4.p�3}�3���3hNQ4+X�3�$�3��h3��3^.s3�l3���3p�E3y1�3T�3���31�a3��3�&-35�3a�l3~tw3�03��3��3u�3�ҵ3���2N�3��4�r�3d�3��3ԊK3t,�3��D3GO�3��3��3�3P�j4~�j3�3S��3���3�0�3��3ɀC3:�X3�'t3`��3Z�e31�&3} �2���3Ng3��
3��%3u�3��2�Ov3��3�{�2Q@3!�s3�?P3N��3��3�\�3R�3ܰ�2��c3)wZ3�]c3��2�?\3�2=3�O3^''3�&�3I$'3�}#3�'P3�5"3юX3�n�3J�23[�D3�a`3���3x�L3��R3D��2V`3@�O3��2�h03�wP3�B�3X|53k�3�zO3	~,3]��2�	�3�(&3'�A3��+3�*3�=3uS�3�`�3���2z�93 �3�Aw3��F3P��2��d3���3%?23 g73��+3f�]3��;3Zc3��x3j`D3��3ل�3%P!3�I'3UIo3<%3(Ny3=�I3江3�3tn�3�ڻ34�k3��w3c�2fK3=3�H
3��-3��3��3!
3 Hg3�w3��53Ƈ3g�3s�21U�23x�2`533ҧ73��P3�d03�2Uq3#��3��3�S3��2Y�^3b�3`@3-	�3	 3%h3��03���3�V%3O�e3jN3e׭3��=3�Î3�'3���3ƨ<3RdL3(Yh3= 3#�=3�v�3'$�3@�3��&3E�y3&�3��3T�q3�306�30|3gd#3��T3p�03�2��47�)3�Ah3a�2�sA3�3�733��*3��3߲43��3U�13���2L��2�.H3��3��3G�:3F��2"�i3��%3��3�<3�'V3Z�'3
�3"�83��2'`Z3�mj3'3X�351�3�j�2�3�3�_Y3�P�3�8W3�36m�3ra�2#(�2ٽ|3V:�2��i3^3BV�3��J3��e3��3��3 
3KU431�P3ވ03�.3�43��s3,�3V3sҫ3�ʞ3��[3�l837�X3��3��3��}3v�2X�3�'�2�}�3��3AF
3G�3T*�3F�2�/q3&rv3ٙj3G�3K<43��B3* 3�1H3f�3MB�3	�q3Mb�2�jO3eT3G��28J�3��=3S�M3�3���3�A3]Be3#�A3���3��e3�3C&M36/t3��13��63g�3��3��53Y3$v�3�]3��33�kJ3��3��2���2�3�T3��3���3RU3"+W3��13��3�U�2�cX3�]p3��3kJ3|Q�3�jL3չ3��3?JZ3.�3ks�3�B�2Y�y3�3�3U�.34�[3Pk�2~r:3��2�aK3�P�2�n3���2%��3�s3��e3uP3X.3�l�2�
'3j�&3���2�[�3ȇ�3��W3�D�2}�2΁l3�<t3V�53��3��3��3��2�tu3c`�3��,3���2"��3��3�53��Z3pP^3{Q3�φ3�	[3�337Q3���3j~�3��z3'K3M�s3��C3>�3�at3�N3_ǎ3-83>�3�T"3�+3to�26y�3)�3x�03ŨD3:�k3��2��j3�%/3�3U�3���3a�J3�=3FEN3�,�3��@3�L�2	-3K�&3�3�3��93�N�3P%3Ҋ3"`3N"�3��>3��y3�!�3�3��30j3�!3�3R�<3�x3���3��M3X\�2>	�3lD3UII3�Ng3�A3�'�3a/3S΢3؈#3�43�3� �3��3�{S3^il3x�k3J�c3%u3¿�3A?3�q3��3���3��63i��2�	�3�]U3�2�j3�#3X�3x�|3�۵3tb3��d3�*T3���3m�K3S3<j03h�z3*�g3�Y$3>�3-�U3�ȍ3�)�3x؝39�3h��2�u3C�33��2?�T3.p3��73{k3���3I�3�@�2T63?.�3�v3�)3�<3f�!3�%=3[��2x,V3[�3f!�3��3,�37Z�3�Q�2"Xp3�H3z��2��\3{�73��3%831n3�#3zl3U$&3�[
43�3�� 3�x�3 3S<'3�@T3�q3��2�3���3�x�3���3D�2k`;3��23�3n33��2�=}3���2 O�3ڃ3��|3��3���3YFX3JB3�3�2\J3�� 3�3��363@��3��3]�]3{�H3@3�t�3۝Y3"~3��)3�t�2a�N3/83�6b3]W�3�'03��3i��3y3��W3�'}3Xa�3o+3|�3��T35�b3�<�3���30�3G+-3��&3�'�3xl�3��3�F�3 �T3A�-3��.3��4s�=3��3�$43�D�3�x3��53gV_3��S3��3��3Y>�33�>�3���3�3�O�3_�3:�F3�\W3X��2�߂3�׽2��t35`�3���3��s3�!�2�6:3�й3��<3���3�3�&3%�3��V3���3�Φ2�A�3�'�3X{�3�CF32�2�H63�R3l�.3Z%�3��E3&Ɠ3w\j3�4M3/u�3�N#3���2��3:ס31W(3Zvk3i�\3�N3��\3�|3Y8?3��-3W��3���3���3��.3!Y3�|�3�^f3
�a3��3E4� �3N�3o�3F˚3��3��3�,e3��I3��3Z/35�3�^3Iv'3)�2FZ3���3�F�3l�c3��'33�3h?x3�� 3&I3��c38KO3��@3�|x3�]63rn`3�m3;�3k�3o�3��3R��2�U�3���3�Y3b5\3�@3b��3��4�`>3P�39��3�a�3@ʐ3��3��2W<353��3T�332'Z3�tZ3���3#�}3s;83]3�>b3)`3(=�3x�3�b	3�[3Æ24݉3Q�3g� 3��3�K�3v�3x��3��p3i�3}�3�Z�3��3�Ր3Ֆ3\�4]!C3w��3�{3!
�3�#3,��3�33E�,3��3��3�ۈ3h��3U�'3�t3�]H3��3[�]3��\3��3�r3_��3EA�3W�B3\��2��M4���2S�|3��03��*3�A3W�3���3�¤2f�o3�o�3��3
�r3-�$3�=�3�̰3��W3�7�3C{�2�^�3'�>3���3fz�3	��3@Y3�\�3S
3P9N3U�T3�3��E33�H3_�x3a0Z3�.P3��3��j3�kN3�� 3]2\3�h3:.31��2��"3#[?3���2v��3e��3�,T3
3��36� 3zV3 �Y37Bn3���2Ag3L�34�36��3�3彟3K~38$3�h�3�c�3uL3�&3P< 3�n3���2���3�a3I�$3e=(3F�3L�:3�@3$%3�39�3���3}g�3\?�2��=3���3��3?/3V��2���3A433Y��2��}3�3��3�l 3yk�3�AO3���3{�Q38�4��_3�q�3��&3��2�d23sT,3+�3�IP3R�b3���3NV�3@3p��2i��3�"O3�J�2ADz3c��2��Q3��93�ph3 �e3��w3�l�2k �3o!30�m3�1N3��-3�$3�g3�\_3?�Z3$�\3��%4��r3=_3�'�2�8�3�w�3C�>3Ǒ,3�@3	NM3�3Bs3;S3}i13M�r3*�3�>?3+/"3��3��w3ob�3c�Q3���3 3�3�d�3�j�3��?3~i>3� 3�H38�?3xΒ3Q�<3/�I3�x_3l�@3.OG3�Gn3
s'3�7�3f�3p\�3�!3�r3�H+36�3��t3ه 3�aW3�53;
�3�'�3�c�2�P93�qD3TeJ3��3���2�}]3���2�z�3MD3��#3��G3�S4��3GT3�|`3=�@3��3'�|3��3�2>3dΠ3+9�3}:�3�v3�u�2a|J30]?3���2��y37vs2�YR3��A3c[�3�q3���2ѩ-3�U�3o2�2��X3g�t3>,3m5J3�-�3��3,$	3t��3�f�3ZɃ3h��3t�3���2��3EB3^��3՝23�� 4oj3��3��[3�`n3��2��3y�$3n-3@IA3� $3���2�/3��3���2=�3Mږ3�#�3�`<3��3�`a3g�f35�03��53��2�Ց3��3�E�3�}�37�3m�W3�v�3��R3�YI3"��3��k3��/3���3YW:3x�:3�3MY�3�\�3��L35#3���3��3�J3�P�3�EP3��K3/��2;ͬ3���3%�2�53���3��^3a?�3(�d3�ci3Yl-3
�3�,m3�~b3�ni3�!�3:)�3���3O��22~Z3M�u3�q3���3m�_3[�G3|!3��w36��3+�3aq�2�/�3u��3��3&PR3�N3�R36�d3��3�@3n�3�B�3Ȑ3�{3�k�2�Y�3���3o��2��3Vr�3B'�3P<(31��3�HZ3��73y�3�f�3�3Be3#�H3���3nE3�*?3�Py3��	3L�E3�u�3�rh3s~�3*��2�)u3��^3�
3t)3F73h�&3Lu3/��3��?3�4F3E��2���3`��3ܻy3&��3F3Uu3��3n�3�W)3�8734��3.9�3��3��21��3�{.3#35F{3�S3��3[�3T�X3G@3�E'3��3<~�3D_3��[3lG3�d33I213�jR3�=�3� 	3E�:3q��3��3;p3�\�2�� 3q	k3��3�B3վ3��3ze3*�P36y3��"3�X3t'-4׭83ɀ�3tO�3��3K|(3��?3VL3�!3�wp3&��3Ξ3��3n��2�Ce3|Q]3ZCs3��{3���2)m3��,3�E�3��h3�a3�*3kD�3!m3uހ3l�z3�N-3�l3)�3��3P63G93���3��3�t�3��3(q�3� �3��3#�3�3���3�3`_r3*U�3"&>3�p3Y�4uq23���3�{#3�(3��Z3L�v3�3k��2��h3F��3�C�33���2��]3*�r3��q3�L3�4E3�Ǖ3�+3�Ӎ3��J3n��2e�2���3G}3=��3�}3m�3�3#�$3n<3���2_�[3��835V�3���3=�3�`�3!�93��(3Pv3��3.�3V)*3�1�3��34_�3���3��4�<�3��4o��3�41�4Χ4���3j��3-r�34�u4!�3U�3ٮ{3:�3	��3�ɟ3��4m��3v|3�v�3H�4��4m[�3�.G4;�B4�>�3���3�ܧ3_	4�	�3K4��/4џ3kW�3?��3qH%4f'4 �3�="4j4ƛ�3 J4�� 4$��3�@4��&4H�4��41��3��J4N�g3H�3"�3�{4��3�[�3��4#V�3~��3��B4��3�9�3�y�3t�3�L�3�jf3q�3�ݼ3	��3��3�n14�7�3ct3v�p3�VV4�!�3Y�3E�3�"4#@3+�-4F��3�_3�x�3!{g4���3^��3��}3y�.4��3��"3VW4w+�3&��3=�3ɸj4��3�ҿ3�s�3�@4{t�3�u�3�f�364�3w	4@�3��3�b4Ѷ�3��\4_��3#ϑ3༗3SL[4`�	4Oh�3�.4���3<r�3
��3~�'4��3��	4��b3妍4oj�3�64���3b��3d��3�zv3{_4h4�3�� 4�P�4�b	4��4�ܢ3�:"4-`�3}]3�b�3��3pD&4��V3)�*4�Y�3E�Q3GUF3|��4�4��3���3�=4���3�3-��3��a3��3 R4`�64��l3Ý3/�3�G�3<�b3�q�37%�3P��3QYu3V�3d?�3"4��r3�4 �q3T�3*s�3E��32�3�H�3 �3>�b3)`�3?D4�`�36#w3W�3!�	4+��31�3:=4�Bl3�R�3m�3&4��30��3���3�r�4�C�3Y��3�4d�3��3<4{��3V�3ߔ4�4@�34���3=	3���3��3�g�3��3́33X4���3��R4!B�3/�f3�uW3�/�4��3�]�3��3hq3��3�I[3���3v˻3�14b�-4aW'4���3��3�4�}3Yn�3��3B�v3��3ݏ3�c4��4m]4�$�3]�4s��3��3�l4�y4���3�I49��3��[3�j�3g�4
4� �3��46v4R�64�1�3�S4���3�z+41��3�4���3��4%+*4�A�4{��3{Y�3_��3��/4�!4�QR4:i4��4�(4�24�n4;�4K�4�
�4x�3��P4j�34�)4y��4��3���4��4ìS4�K�3A�*4�4!��4Y�4�,4vX4��3?�U4.��3$�!4I(�47>_4��4�h�3�CH4��3���3�X4|��3�u4�R�3��{4YS�3�2"4F+3Z܆4�P4���3!�3��I4�:�3�%4-A4�<�3w�4�e�4�+4˓4���3%~4��'4�-�3��84��3�Ў4���3��@4.�3�Q4g��3	�4�O4��3�C4<n�3�k�3��4.,S4�ƶ3���3�M`4��R4�O�3�U 4(��4�r+4��f3��4G��3�Y4˲4��4GH�3R�3*�4�Nb4j�M4�df46^ 4�P4h� 499�3��E4/>�3/�l4b`�4���4WD4�3��N4��p4Lڝ3'�V4�!4�M94�̌3���4�d74k��3���3SQ�4���3��4(�4�>B4�p 4��3,7 4�~4�[4�<"42�S4m74D�|3��4���3���3�m$4pߒ3�s�3���3���4�\4��.4��3��=4�\�3j�4(u�3A�&4���3|y�3��!4��p3���3\sm4k��3Q�'4<��3@�K4~��3H�3Z�04c0G3�T4$4�3)e4
�3V�32;4�^�4��	4�%"4z�(4��3
�3t�&4..4��3`�4p��4^xj4��I4$��30�S4�"4/
4|14'U�3��4ټ�3*�4�3��s3�R�3`�4��30�3���3���3^�3��4.�4"��3^�,4\ ]4�:4/K4�KA3ÿN4��3���3�j&4%��3��44���3�d�4w 4�@S3�2i�3�?'3(�o373]n30�2�L3��3W�j3�\*3���3GĄ3|�[3c�3��3��3��2�0 3_�Q3cݙ3�N3%�o3��3�<m3		�3�j�3��
3�@3�(3��?3�~�25_u3�Ë3�3BN33d4�>�3��3ݹ2
MU3�\�2/L�2i��3�-�22�I3�3�Xl3��)3�Qw3k�2�4�32;3�+h3�13�?�3�2�BA3�p�3�3��z3�P�3~U�3V��3 Y�2D|3��\3�e 3ڷy3�o'3��3��3�>`3S�H3��3�De3��4�.-3�K3���2��J3ϓ3�C3��{3�v�2�l3"��3p5j36b3>�2�3�y�29C3��Z3��3��|3�!�3A�X3��3�e3t��2�a�3�d3�^83�93x�
3��R3��3�bk3f_>3�O3H��3Ȩ3
>c3-�H3L�3�V3�#3̲�3
��2H��3�G3 �n3�J3�W3�3�h�3CD�3�>W3��F3�G3�-=3�mQ3���3���2E�T3�y3���3�Oc3��3�z�3bF�3>�<3�DF3F�[3u�q3GM3��3�*3J��3�,	3�4Zv3��3S�p3�+3��
3��)3�A�3��33��=354Atd3�/:3B�2�Y�3'�3��33ԇ�23��21�3�"3�-f3,B	3��P3(�p3�s 4X3��c3��33=�K3;�3�چ3z3r�2RN$3#�3~�3�d3���2�%�3I��3�03��X3�*-3�f3��>3~��3�Î3W�2M�R3�-4E�93�\A3I53�2�U3��3|M93���262F3)g3�j�3�j35�2$3`�Z3�|�3�Po3M��2���3��#3�qo3��m3<�83>*34�4WT3�m3q�]3�o3��2��93z�p3�53�4[3%��3�ρ3��3]O3��3�p53Rִ3��x3�<3=�U3ؼ3�m�3Q�3�.3�]3vb�3��3�pA3�"�2�Ԩ3S�S3K�3��3�l3-V�2��k3o�3y:f3$��24Y3��!3#X�2�b]3��3��j3��2.��3CR?3��2_��3�ɕ3�$q3~:j3�{C3�33Qi 3�*%3[v3A)3eE^3���31uq3Ă3a�_3#S�3�43�{$3��3�0@3�KD3b 3J�3_3���3 j3ߒ3�ɇ3Uč3�nw3pq�3�G3�X3^��3�>T3�P�3d�3t�r3M�)3w�(3(�3��3�f]3�r{3���2�ٚ3�
3 Ng3�3�ٯ3�E(3_�3W�+3�c3��U3b�3��3�(�3�W�3z:�2�J3��4�O3ɋ3g�*3 +�3@�>3�(3�e�3T�29y3�!3j736^3�2A3%&3!�:4���2� .33r�3�13�Lh3<�:3�h�2�Xm3�=3#҃3��3
��2g�:3Fu{3�,3�_3<+�2�uq3Y��2LkR3�"3��3?�3��4��43�3J��2G:3�q3�F34��3�13Ӆ43k<�3�&�3�63N^ 3A��3y�3$�3��Q3>@)3�~3�J3(m�3Z�P3{�3��2�]�3��3�VM3��G3sl]3z3�63d�3� �2�v3O�3�a�3��A3X�2��p3d�
3�p3R(3���2xÁ3���2�{�3/�y3�1B3L�:3��3�ds3Яy3��23p�w3�m�2N�O3�#C3?;�2!�%3���3 ��3�ht3��$3:S3�VT3��2��/3TG�2���39�3i�I3�ta3��:37�J3�1�3įG3�A3j3JJ3��3�l�3uf@3٩83��w3��3�]3�xp3:f3�ʆ3 ϋ3\S-3�~34�3l]3}��2�0�3Ar3��3��3(�3.X�3��,3	�3J�X3z>;3��w3���3�G73D�X3��31��3`�<3�G3�
K3��x3^fU3�[�3���2�
:3J�3ڤ3��3ޣ�3̓�3!
�3�3j�l3�F�3�ޥ36�13�W�3|��3d�I3�j$3���3��3�#�3��F3^Z93�^h3�r;3��:3m�R3��3_�m3@�3�|�3.�3Rm31��3�*R3��3̾3�w3^�E3L��3� j3\E3,f�30�D4���3F|�3��C3Ñ3�
�3y�3�h_3ؓx3�T�3SL�3�^�3nL�3��3�@3è�3�i�3��3�0F3���3��W3�$J3'<�3�BV3ۊ�3O�4�4�3�]�34�=3�;�3}��3\|X3�Е35��3���3��@3��3wĒ3,k3��3@$F4��h3T5B3��32�13�[32�3З�3�)=3�qL3��3�k3��3~�23E]�3��3�U�3u8�3��p3��3�$:3Y�3��$3:3283
�4���3&s�3��~3t93.�3���3��3�&3-��3ԋ�3�a�3:��3�2��3��3+�3R��3�-3�ϝ3�͞3pa�3�;B3S�3�z3���3�:c3�]�3D&o3n3��3ݒ�3���3��3�3�3-�3܏3?�'32�w3��3��=3_�3SM�3@�3��G3���3b"G3}�3�$3F�O4p�P3�w3$�3Ń^3�М3��3	'�3��!3�~�3!�4Uͦ3��_3"�q3��3�P3��-3�V�3p�,3;3��3�_�3� Y3�~3�q3`��3�E35�c3�}�3	�3Ly>3Ϧ�3ej�3c3H30pW3x�54^�3b�3̺�2��3���3��3���3�7�2�@�3�1+3���3�e>3��3N�23�,*4�S!35�30�3�m3b��3�IT3z�I3�<m3%��3��3)�4��3�iC3��43#ͬ3K337Ci32�*3��3�j3r/�3�X�3c;�2�t3Ω04{J�3�*�3)�3dM3���3b�3a�O3��:3" �3��4���3���3sU3�c73���3c�3��A3��"3�
4a3�`�3ƕ3O�*4�Č3�4Q��3�f�3� W3�Qn3�-3b��3��o3',3k�+3���3� �3�Ē3�4*3�{3�8�3+�3\�W3��^3���33�D�3�3)<�3eaR3��3IB�3Ӑ3� ;3�y3%A(3�7�3��3�4	3�@L3喘3@��3�3��2?M�3~��3t�3ph3,3�7�3@I3�$�3��e3w[>3_�P3�4=�P3���3�G_3*\�3���3�˙3��g34U3/T23:b�3��p3��4�E3��3��3��#3C��3p<M3�m�3���3�u�3u�V3���3QN3Ħ=4�yM3g�v3Q��3� �3�G�3Fֺ3�4G=3���3
a 4엤3�ڟ3{�%3<
x3���3��2�3�p3�8�3 Nq3 !�3��3���2��
3�!4���3�z�3?�3��3��s3�}�3$S�3��F3�G�3�[4Ȅ�3�7�3i3NF�3�4�3��.3���3A�>3�Π38�3C��3^�3 î30�U3ԇ�36:/3��3��+3_҄3=A3ߗI3>��3�|3N�l3�g�3�؎3��{39��3��33��3�{3~'�3F�3�+�3��;36��3���3�I!3d�3��3�j3o2n3��3r�3ԩ�3���3?��35�.31��3
�4,��3ӏm3��!3~�3�S3�3>9�3\�T3�3�3�~3*@�37g]3�<03^h34�	#3Sw�3�j3OE3�~�3۾j39�3%�3�I�3��3��4E�s3�AA3Py�3���3�03��3nI3K~�3�o�3Zi�3<�3��,3�v�3��B4E�:3f��3\��3��3{�3צ3���3q
3�3��44��f3ſ3���3j��3�3_J�3
�_38A�3�p/3
4Xs3��3=��2�j473C93�l�3��Z3�Y 3���3p�`3^�2*��3M�3^�3J�3}��2�<38��3:˄3~(3�a�2tS�3��3�̢3&��3<V3��l3�3�N3�*3-�3�ڊ3��U3P�o3�[3��K3}L�3���3�?�3�J3��2�ٰ3��m3���2O�3��A3J<34x3�ױ3��;3q�)3���3�A�3�3\ 3�VB3�{)3G= 3e��3K�b3G.53�YY3.i�3�ސ3p3a^(3��P3 I(3|�3�JB3��#3��Y3��23A4�3�w�3r�.3��T3N߆3@�93�VA3V/3��,3��2aN3JK\3�=3��!3!�3ӡ�3m�03�o$3�%�3��R3�&�2��c3��`3	�%3<�3:��3�K�3��L3�O3��	4O�3DJ3.13�L3��2Y37�Z3�(3��3�\�3:��3��S3���2�y3ڞk3��i3J@3�O�2G�3�K3]W�3*S 3��3 �2���3 3�)3-a3j�3�Q34�38W3I43	�s3ہ�3�Ɵ3?�E3�^ 3+�q3�3 3I3�g3���2�Fk3q�3Y�3�I3k:;3R.3��3�3��T3�D�3X��3�)$3H|3�Ҋ3�#�2�V~3g9C3���3��3�@53�m3gw�3�3ݬl3��2�`g3j�63h�:3��>3��R3�3gN4��2(��3p��2~�73~��2��33�1r3�93e�3l��3��C3�Vi3Â3d�f3D93?��2�?p3���2l��3]�:3m�/3z�3�� 3�3�2WH4D�"3�53��2�(3�3"A3��[3�X�2�H3���3�Md34�2���2>03^zs3b��2EIG3r��2*��3��3�g�3Y��2�Ҍ3��<3�^ 4O�3�B3�[23��l3��37
3�hc3P�28�,3�R�3{֥3�V3�I03�q3��3��q3�=3��&3��r3Q�2!!�3�;3uL_3H3���3Ր3A�a3L-�38C+3|@23]6^3��3���2peT3X	�3�o3�U3�I;3w_]37��2��3�C3���2[�j3tT3 �3��3pϞ3� �2�|�3>�c3ga3��39463�R03��3P(�3���3GW3���3*8�3�W�3���3Z��3ޒ�3��33�F:3�e3�Vx3�~n3I��3�X�3��3D�I36��3�.�3��3�W�3p��3.�3�3�q�3��3���3lċ3�'�3aFq3�G3���3lF�3	��3&�q3䘔35�$4s�3��4��3�YG3��t3#l�3~GK3C�c3X��2�0�3��3Զ3;l�3�a�3F��3¥54�å3�nR3I,T3Xw�3���3��3��3�d=3��=3��30�#4S�e33uI 3#�243��3AX�3�!�3��4��/3�3M�3S-*3N9�3 /43�3�a�3Ю�3ϡ�3�o�3!��3�Q�3�g�3�$�3&13��3L�c3
�N3M�3 h4�̊3��n3qu�3��3=�3ݺ�3T��3h�s3��{3���3���3k"�3�`V3��3���3T�3�@�3���3yj�3�M�3���3Ŷ73{��3�N\34�Ҭ3�04XJ�3b�3૶3��3�@�3D�U3��3[��3�e+4֊�3�TU3��3���3P�D3�'�3s�c3
A�3	��2��3�{�3�n3"x3��E4�[3��53�t3xH�3���3<j�3ѝ3"��3�`�3
�4�M�3�{Y3�E03Ƽ�3xtQ3"�H3͙�3"?#3?��3!�H3��3E.3/a�3 ��3�4�F3z��3G]�3�f3=O�3g՟3�Z�3�X3,��3��4S�3��3��{3);�39�u3}xI3�S�3:3g3���3�t3v�3�Y3-TD3��3}��4�L�3��l3.F�3{�_3��3�.�3構3��2��3F�>4��3J6�3|��2���3p��3��e3&�3,m3���3�2D3�4�7�3�N#3h�y3e�o4�+q3+�3��{3I�Q3]Q�3K�3>C�3��3=��3�n4��3cf�3�3)��3jxJ3p3�7�3��:3'��3��(3�*4�bx3%�@3	�2��x3T�3h�3A93L=?3G)�2��3��3���2��2-B3�P3U�d3��3/�~3�3i}�2T�S3.�R3|5�2��&3�[3xo$3�g�2}��3�=�3��2�s*3J�,3�%P3JGF3�O3�RM3}��2��
3�P�3y�!3�63ƥ.3K8�3R3j?3j�'38#`22J�3 C3��l3:.3�r�3��2M�53��3���2M�3��93���2"`3$G3��2&��3��3��
3q3�D3G3+3k�3���2��b3�3��3Le]3uT�3d�3�A03p/H3��3�P3�zR3W�-3�� 36 3��.36�d3��2��3�]d3�K3��3+Ѷ2�	3���3�N�2�q�2Z�2T�3P�'3��B3��3�3�'3{��3_�3d�3��2�T3��2+�3�%3�3jC3��3T�U3��2��3��h3kZ;3���2*�53`C3V+%3z3o(�3��3��R3~5�26�j3�=3�\)32s�3�>3�'3��2PU�3	Ȍ2�H3`��3��n3O�3/�2�_m3~/3{3,
D3�*3X�w3(b�2��3�r3�_N3�I	3��3��3k�%3��3��*3(�3���2/E3�,�2p��3C4�3�3 ,3�3��f3�\3�� 3{�*3"R�2�r73UE�2ջ�3V3��2Y�2���3�ˀ3��D3��-3|�3ݘw3�!3H�3���2��83e@3��3�`Q3{D�2��3D1p3�2�3w��2��I3C�K3~{3Ai�2�M�2�r
3�P�3�;3%Ns3��3�M13�3��3Y@3d[3yEM3��3��4�Q83I�2g�[3�V3ބ3)2.3w�
3�K�3���2�EM3��3*��2M�3�_�3 s36'3�3�aL3oU�2l�33T3	�2�v93j&�3疄3߉�2�c�2��H3�A'3H�2Z0@3�P3�731T	3-M�3z�3N��3!�2A�3�C]3��/3<��3��3L-X38�3B��3�:h3/k3��3���3���3$�\3J]�3��,3��3�	�3F?�3W��3��E3�l�3�؜3i��3պ�3�,!4��3�x�3XEQ3���3<�E3��3�z�323뚊3|��3�aO3��3-�L3r��3�Wu3�nA3��Y3��p3	&�3��r31;�3�[!3�~43G�3}�48�^3,J<3M,b39��3F.,3S�]3�ř3�+3���3�-4���3m`3�� 3�{{3Nէ3��53��3^cb3�P+3�T�2}��3rO�3/ȇ3{��3�4�pI3���3_[3�A3��3�43Y�38i3CQ93ժ�3�o�3��3ރ�2<��3��Y3�i3�C3�U3_��3�;3���3�H�3,93ƴ�2p4�G=3��]3�3o3t8z3.\3�b�3%Lr3�-3��3,�4tHr3��3�'3���3�/g3Z�2��3��$3�j3�M)35�4	�F3BL�3)>�3���3�IR3��f3��3��3�ڌ3���3i��3�j3�H�3A�43�3J�3'n%3KW36r(3��s3�3j~3K��3&؉3S|�3�13m�{3�1N3بk4�0Y3[�3�_3��3��(3kJ3�p;3E�3�Ė3��?4�Ο3��#3�-3Hfp3K��3t�3��4�|:3�f�3�Ek3;��3��+3��"3m)3��4|�.3\zs3�l3��3��3��3<�3a3V
o3���3f&�3O��3�X3��3�`�3XH3O��3Ȋ3�Ҏ3��f3\�3�63�Q3�)3"�=4k�o3j�3�x�3��K3��F3��3�p�3w�3�`{3���39��3ۦ3�"3�,3�}3�Cf3|q�3n��2R�3�]53��3��38��2Ο3 [b4�IG3�W`39:�3j&3��M3��3�;�3��23i&�3·�3r\�3�LM3J�2cI�3�x3��R3��|3��3��k3�H3��3nY(36�32�3���3�o3J 3���3I��3�3�/3FO"3ښ83%Y3?o�3,Q�3�8�3#83�`3�T3P~3D^3�Sd3���2��s3�`�3���3O]%3n@t3�v3v3�=l3�3��j3��Z3�{�3l�3;̘3�?F3Cq3��3/!�3�w3n+�32p3�T�3�x�3!0C3:3r��3�}3C]�3��l38�q3~�3}O73J �3wC3��63��3�̓3�S�3qd!3'>3��4�^�39�D3/��3�H�3���3���2s37�y3n��3��b3�҇3�13d�T3�#3׋3+.�2�ǌ3�1(3�"3�x%3.�\3Sb3:}�2�]3*u�3���3W3T -3��3k��3Ub�2C�3��3���3>83�T�3b]�3��A3p+3���3��63�1X3)�93�O3�Ye3J?�3��M3�"3�3���3�X3P�3�]33&}�37�Y3r�3"j�3�I@3'�3�3q�}3���2vQ3�0j3�@54�DC3TWq3�B43�&�3�rq3z�u3i�C3��$3�u3O�4xPZ3��^3�yF3ժ3�z3N��2ޱ�3(�3���3�]�2�J�3.-T3b@3͞�2�m4�&3�f3���25�A3u8m3�23��o3��2v&3���3qc�3>�X3a��2�-3J)&3�e3X&m33ů2�Հ3J�3�}3�zX3Z�3�rj3(B�3�^{3��u3x�,3���393T;3e�s3��@3s�>3y��3G��3�\3��3g�3kj�3W�13o{�3��2�<~35O63��34`3�a%3+�@3�-4�x3��o3#ɠ3�,3��3<A	3��X3v:3`�e3a��3�ګ3D�k3X�2�Zu3rג3��]3B�k3	�26Ǭ3��f3	�3Oϊ3W'"3��324��P3d�^3}Ǽ3ץR3v�3�K3�v3�,3��396�3���3j�u3z 3�3���2�33�A�3��2Fb�3�93��3�T3�+�2?>�2R3�C3K�=3���2,�2�2�,-3���2y��2�:�2��I3.S33D�73���2��3�v�2-��2��2��
3`c�2�Ѩ2p�3Ą3�k%3yg"3��H3k#3931x3�K.3��[3|�!3�y�2��2D
3�Ą31�3Eu�2��2��;3�@3`��2� Z3[�30�03c�3ӑ3]��2��2R�	38u3�j�2�(33H3=�2p�2�53^k%3���25o!3�_�3�C3� 33�2,��2Z3>Ź2�3	�3��2�s�2z�G3>3��F3?��2��3��2���2��53R�>3ܞ2܊B3�)3�3[63�6~3�Ou3��2(��2 �
3�
3�)�2#��2?c
3��3!�2>�%3V(�2I3��3�֐3���2��2� �2�t3�!3E�3|NP3��2��&3Mʈ3�=I3j3�Ȝ24$#3��3G�2�3(��2N,J3�p&3�C3�I3�g�2�2/�3y�2�ȸ2�A3gG3�R�223�W53�1O23��l3��@3(�3�1�2ӗ�2��63�d2�13:2�2�33̩�2�s3�p3у3ɪG3���3
�2��313Cz�2��
3��2�"3&�3a!3��g3Q�3e�2M;�2;�h3Ί�2�T3�.3 ϴ2o3�	T3��R3t��2�3~_�2n��3Ε2W�=3�L3���2�3�i3�3��2�23��3[1i3G#3Yx3g�s3��3H��2[Ez3a��2b�3�2�2���3���2��2���2�}3���2��13{:f3�3��2P�3��3Ϳ�2��:3�r3Ńj3�%%3���2	�03��2���2�K 3T�2���2�š2�Z3F*&3��2/y�2���3��N3�F3��L3S�"3'�2��2	�>3`�2µ�2��23	�y3%��2#��2�j	3]�I3���2�c!3"�2��^3�1�2d�[3i3倯3���3(G(4�&x3��3ɏ�3��3��-3�5�3~��3[��3��3V4S�3w�4A��3��4�/�3o�>3�3H��35L�3���3��3�}3�_3�k�3��64�fq36x3.ŵ3���3�3_�}3�C�3�,3�p�3m]�3��3	��3)4M3z�3$�3�&'3�nf3�k@3�Ғ3h��3
4G}4��3Bi�3BE�3٧�3�ݺ3�t�3�?�3y�3�۬3Z
�3�F03#��3��4b4Ś�3�3���3���3m:�3�%�3�Q�3sR�3o�r3�T4HN3���3�	{3Ÿ�3�HV3�X�3Ս�3/.�3Ȅ3���3���3�R13��3��:4g�3�>3~�(3Er�3��31M�3;��3�hC3 ~3�ݖ3�u	4ɇ�3A$�3�֟3��3mT�3%��3Kc�3O��3{�3�S�3A}�3Y�K3�,�3D��3��4B(�3�03h54)G�3�c3�3�.�3wi�3�G�3��3e�u3ou�3�[�3��	4
�3Ff�3��3��3�m>3�|�3�ٗ3|�s3D��3���39�4�w[3�{3���3�S�3�r3` �3�}t3N��3���3�0�3�l�3H�31��3$342�3|��3�˓3	�@3�`s3�C�3/�3>�+3��3�м3{I�3��X3���3]l�3;��3Ô3�؎3�mt3j�3
�3��C4���3y�m3_�3��46M[3ֲ�3�8\3�{x3	Ð3 y3o\�3��|3�J�3_4�:�3v?�3��v3�7�3k/$3u�3帲33�+3���3y�l3<��3wh�3|��3�m3_u34��b3j��3��3��U3�.<3YlE3��48�3�ُ3/�!4|��3�ب3���3>��3ڕ�3n{3 �B33632��3�W3q�3�O�3�/3Q3043�=38�39��3[]�3Ϸ�3#Zx3�Ҕ3 ]c3,��3:�3���3�h~3c�o3R�3kT�3���3a��3���2;ބ3�k&3��n3��3��v3��3�׼3�^3�
,3��M3�h{3��V3��y3��t3�<�3��3���3���37P�3�&3�x3[E�3�ߋ3'�g3ŷ�3F�3�K.3զ{3>��3굌3�ܙ3�3�$�3
��3�#�3�O4}Z+3���33t�3�;n3�3|3�y�3e��3'��3ȓ;3o�3�ȩ3�C3�C3QO�3Լ3=zM3��3]��3U^n3�s3z�30NG34au3�=3��A3eIN3ŀD3G��3L�:3%�I3:�3�i3��e3�N�2��@3�)r3��$3pF�3�hT3��g3GEQ3QІ3�u3 ��3n�2~��376=3�Q3ޤD3r*D3���2͞w3�n3��2��]3�	4ɀ�3���2B��2���3�z3�`�2%F�3-Q&3�{�3U3�0�3�|"3�ZO3-l�2���3��h31Y3�;3�.g3$u]3�-E3.�K3�/3mi�3��\3�F�30)3�:�2�;�3ô�3��N3�3i^3�5�3�+31^/3O;�3�H3���2U��3Ãz3ޥ33�73LN�3�J3z�3���3;��2���3���3�x�3�+)3��2�#3X�J3��2��h3Ë3e��3l�v3�$�3�`I3q�&3$��2D ,4b�<3$/3R��2�Sr3�)�2ׄ�3��T3-t 3o]3���3�;�3�\3��2�~�3"�30�35J�3�y�2�`�31rj3<��3���3UI)3��/3���3i��2�A�3#k3a@M3ܬ3��G3x��3�W3��:3��3��3���3��#3M�a3 �3�$3G3�()3K��3�%R3o��3T+N3\3*3��-4$э3|?3
J�3�j3�[X3���3��/3m3�q�3W��3��3�4�p�3��x3��3�N(3eV�3�Ԅ3�/4�R�2��f3��3�l3N�2 Z�3�	3�iz3�$83��3�3��30Y�3 �H3]�3�%�3"��3Եg39#3�9�3\��2���2v�3P!3�3+3�o 3ϊ�3��3�e53�	3��M3��3�X3�0:3>63��2��63��E3���2@"03�On3Z�
3y} 3��2c�)3�G31&�2��2|3��3�2{_3:�3��*3c�M3�ؘ3wF,3�p�203v��2��2���3���3Ieh3F	3�a�3�}3w֏3ns�2o�3�oW3�m43~>3o:3�C43�H�25o3��)3%3+I�2��3ݛ3�'43�]a3�13�C�2+|3i"3z�2x�a3�t{3�މ3L�2{^�2�p3�"e3�#3��3<4�2�3��C3��3��U3�h"3�(3{�33v��2�3��3�_-3�jU3��3�A�2��M3�K�3��?3P� 3.�2(�F3��T3��2f�3-�2r�3�3�K3ڼ2��3n3;��3�Z3WQ3�I3��3�t�2 �Y3��93;��2��c3Շ3��u3T 3�Jx2K�g3� D3�n�2�.3�%3�_3���2��3��3��2�O3�3N�V3�?3]�`3ߚ53"P3p�E3�3��2�@3���3�2�3��23� 3�W�3�JX3~13�t3��2lAu3�H3��w3��3�3���2'Ⱦ3�3�x�2�S�2�37
j3S�*3`�\3>��2Z�3q.�3��3�3�H�2�m3�~3��3�$e3�� 3V�^3Q�\3�e3�� 3ّ>31>�2CT�3�2M3��3VQ3�T
3P�*3`&3!�y3 43=\�3�1�3�sj3w�3^9�2A93��<3g��2c�[3���2X�I3��3PG3�S�2,3b�2Z(�363��,3U�P3�+3^�3Λ83� �3F�2C{.3*$q3C�@3�¶3�903��H3�ƈ3��2ߒ13l��2�U�3�,�2�w3�736��2�`!3��3��2pY3��h3C�2��2�bG3�o03_��2 ��35Ϡ3�B�3v�i3��2���2�� 3�&�2�3�s3���35w�2�b�3�
3��%3�@�3�<�3ӅT3�C3�3���3k 3zx3��#3�8�2n��2Lr�3o^�3�j�3��3zr�3��)3�c�2�537�3�3T�2���3D�L3��#39�23�b�3��+3�Tc3,h&3�-S3��3��3e�3��2�3�,�3[`3�qb3��2�ZV3(�,3v��2P�'3�<3G#�2}�3rm�3η3��e3v�3C��3�s
3eF(3՛:3Y�3���2� 3�w3��	3��W3B�36k�3�X3E�2�&d3��)3]D3	�+3��;3�Ɍ3`�J3eZ�3�W"3d�3�03צ�3��2�13��3��`3 �@3cu3��
3L�3�D�3��3r�n3ƹ3��2��3��3�3sD3Gu�2�^J3�'3���3�3��2�c3�n�3�3�H�2?�3�� 3
�'3�v93#>3�H�2�943��[3�\�3:�33V23Q143V3yn�2��2�?j3+�3n|^3�+3Y�3� �3h4!�/3��30�A3�g�2��?3K�A3^�93���2�^83�n�3ê�3��F3�n3�P3�K:3rq:3��3��l2�ݼ3�c3n+3��A3��3IG�2nR�3�#3�t?3�"Y32'�2��)3�@23�kd3���2��e3�MU3��03�� 3��"3��63<�3��2e>�3���2�%3�� 3>�3��3�	3�3L��3
iF3��3,�"3�
3��3e3��3=3d!3�0�3�ݸ3��432��2��3-L	3Z9b3�t3��3C�3��3b~Q3j�!3ϝ�2鈱2Q}3t�]3+K3�2x3x{3�˪2c/3��3,3	.3d�[3Z�k3�R3���2�#3g1>3��3��$3��`3��3���2�3�3E�Y3�o�2�*3�y�3`s.3�'3�|3QO(3�f3�,3��3!3W)3) 3�K�3'b3�C�2�Ɏ3 %B3/>3�D3��D3*
3�/3O�B3	[3�|�3�E3���3�>:3?�3]-43y�`3�~3=��3;ބ3�3��3��3��3���3#3�|�3��u300(3IV^3Bj�3(+�3�Թ2���3\�O3v3��3k��3���3:ܛ3_i3�T3��3�+f33$3���3w[*4b�=3	@c3aq�2��3%3{%�3Ѓ3zS3˂3{3���3�F3+\3��T3B4C*?3�&3�i�3���3!��2�	b3�P�3��3�_3���3�T3A~3k%/3�f3�ٚ3���2v�3S�m3�693�H3��3�l30�f3�K#3�-�3�@�2��w3S<k3��k3��G3c�R3yP3�Q;3��A3��3[S{3-3�}�2�3^�o3�$63$�3��%3��3oRu3��3p�,3�#3���3��3P =3�ɛ3YJ3]�73:�\3��o3[4�3�x�3a;�3S�3�%x3��r3��3CU�3��3��g3L3�3�<3d�k3�Ii3�ř3�3#'�3�3tH3�}3�\�3�S3��3�M�3�_�2,E3B��3���3A�a3�*3f��3Q��3�vu3�ߝ3�723�y�3x��3�(�3� �3ۊ63b+�2�-4�543�~�3RL3 Z$3�.3���3
Ԕ3�N3��d3Ny�3�4�Ud3��3���3Ka3��!3�>{3[S�3F�K3�B(3�Z�3��s3��3�$i3"L�3�!�2��3�Mf3�{3�]w3ˀ�3��3~�C3�lo3�ѥ3��3Ź3�X3�:3�>\3XR-3�:3��p37��3��}3ؑ3��W3l�3�3:3��4'�H3}��3=�Z3��3��Y3=83?��30,
3���3���3��3�<�3���2�9�2.�3v�3�ȅ3.�V3z��33R�2&%�3���3ˎ�2�� 3���3��M3�3�_3'Y3k�X3�3��m3�)3Ց3A��3ة�3�^3�N�20sn3��h3˸53�3%f43�w�3>�3h�3�w�3Bww3йa3���3��3��3�S3,G�3}E3�j�3:� 3^��3��b3K�&4���3 ��3�	:3M`�3�3�f3P`�3���3iLw3Q�#3���3�*�3�3�)�3��4��/3� �3�s�3�9�3i@`3n�3��3��V3N��34zZ�3�)�3j�H3�N�3��e3 �%3�Λ3g3g3;�3��3��3*3o�3MB3w�4�\[3�ѣ3��3���3&�2�%�3���3*��2O<�3q4�>�3D��3�33o�3��3��%3�3��W3��l3��J3��3aV�3��u3��3>?�3ٶ�3�K�3��	3�p3wC3/�f3��3nI53sr�3�*!4�3L�3��g3L�3�}�3&Q�3[n�3�|�3��4C�u3$��3�|�3��e3A1C3��3��3�[�3��39�3�U�3N-�3�2�3M)3��3�X 4Ϣ�3�#�3 r:3��}3�C�3x��3p�4b�$3�~�3��a3��4�7m3���3i3�k4�_v3~2k3��3J�3�+3ڱ�3T:k3qK!3`s�3B�4�x4u�3Y�I3( 3���3E�z3t�3y�V3��4�+�3�!�3jRV3���3�u3�/4t�3"33*�3�%{3M�t3�H�3��3HM83�ٓ3��F4���3�vD3���3��3��3�A3��3�;f3�u�3�]�3D��33��3�UH3��03|�y4��Q3���3"
�3G$3A܏3��4\��3{�P3K�3_�4|�3,ۛ3H�)3���3���3��63^8�3u�3�I�3�Y�3�!�3�i�31�3t�3o�54g��3$)�3��3}�3!�|3k��3,��3�3j՗3NB4^L�3�u�3�	$3||�3q��3>�3�#�3��a3�a4)�Z3�3��3�	N3S6	3��34��3p�w3���3c*�3�GX3��3��3�-d3L�n3`�3(�34p�39�3���3�U_3Y �35yy3�3���3�k3!t�3���33�N3MY�2"�3�L3��;3��_3��'3r)3�93&6-3N�2�573�l3?�_3�c3z�2�Y�3q�d34�3��;3�D3�93�Q�2��S3��63�\s3�(�3��3y�23�k3T�2aV3.!I37�3�>+3��g3�*3�3��F3\�3U��2b3�3pO�2�]�2Bqz3�R�2u��3S�53�B3��3O�"3�f�2��J3j)3Q�3(r3ၒ3�#3�Pw3b��2��3w�x3���3	3o��2���2��32�3�3�D�3���2�z&3�3ͽ3̨&3��.3*613e;N3;��2I�27�D3-B�373�;3n=u3!�2��[30��3�#3])3L��2�be3qZv3)��2��m3I(�2MW3#3��^3��)3_�3�C�29�3 >3���2P�i3��
3h"J3��3�}3���2ѱ�2�l�3�
�3:��2>�2 �A3��)3w�2��3G�,3ㅕ29�;3c�3��3�g3z��2�̗3`)3='y3�^13�� 3�3��2��3�`3�3��3�Jv3c��2C1�2��g3�gq3^�j3��<3�3�[3T�%3�83&�03#3|-�2�V�3L��2�4P3�P=3z�y3��L3�JZ3_�X3�<3�33�@3�!U3m��2<i3�3�>�2$F�3��2?�F3��n3-M3�E3`4q3��3"��3�j�2�^3�2�%3�5�2q�73߇�3��2��2��d3��3�4|3�M�2D�3��2�3}t33��2�I3X��2�!{3hK3so2�B�2_��3�K3S��2�P3��2>j}2:�|3m��2p��2x�-3�C�3��3�f3`w3��@39�33e>3y�3ϭ�2㷬3���2w:3�l>3	͖2��2��
4�h�2��2��2��2V��2|�2f_�2��3�}3w��3�Vx3�|3�u�2&Pk3o�>3�x�2vq3�K 38�3qq3v�N3��,3b��2ƹ�2V;T3?|�2���2,\�2M�3��2��A3i��2�M	3���2i3}��2o.�2b��2#�3k�2�/3���2�[3���2�A�2�E3D]�2�2E�3�gE3�,�2��3`��2��3.�2�U3�X#3��2[D3��Q3Q�33Bq3[��2 V03�� 3�$�2_ �2�I�2���2@q�22�/3���2�Ă2�J�2�K3���2�W�2�D�2���2z��2ȳ�2�73��
3�b�2��~3��2���2bw2�G3��2u2QO�2�6�2��2��2N3�$�2��2�}!3;/3��j2���2�V�2T��2|��2F��2wH3U��2W3 3�733ƝB3#�73W��2�3�F(3�@�2�2Om12
�3��2��2X��2�]�2h��2_�	3���2��22�2m�2 �2�?�27�	3��2��2t�27��2�\3=��2��2)�636��2W�3`�3!�3�� 36J�2���2ֱ�2��13��3�L3`�3ɠ�2ծ3 �2�%�2y�3��B2]A�2,3^�3�'3���2�:�2o��2���2C˾2�K�2m��2���26�3�8�2���2�m�2wu3���2�l2j��2� �2p�2Ù�2��22;v2���2�Ja3�I3�^�2p-�2��3�@�2(1�2-T3PT�2���2�]�2�	M3x �24B�2X$�2���3w3�)v2��3���2�d�2Dk3�3Rq�2H��2�l38�<3�m�2o6=2�*3��2x��2�h&3=_�2��3b�Z2/�3�&�2���2�>'3�ܦ3G�2��2���2�U2r�2�2g��2r��2���2l .3�x39E�2��^2_3�B3�_H3�7(3�
P2j�3�<�2(�_3꒡2sd�2�=�2 q/3�=�2馹2�n'3��2�Y�2��3���2���2y�%3�T:3�l�2m�"3�:+22V2_�2��g2��3�Tj2pZ3�m2;3���2G^M3(J�2�f�3@!g3��03�&3�)3���2�n%3��<3eA"3q
93T�r3Ƭ<3|�W3�3�NM3��3F�!3_�3<3>��2���2`^3f/}3��3��D3��3��3,�B3~3Ֆn3��'3���3�5u3�q<3>؄3L��3'yc3��a3c��2|=�3�<"3�$3�r3$�2Ϫ�3���256�3G�3)��3��2���3�I3�n+3�L3��2�D�2��13Q�l3)93%v3�]�3Y3y��2/ �2{�3�t:3xu�2YSd3TxD3]�d38+=3 �M3(I�2�v�3:�#3�f[3*103a3o�}34303j<&3�Λ3-g�2n�k3���3�`P3Y��2[�<3��w3b�3���2��"3*63�i3���2Qw3-*?3r(M3��2N�3=4�39�,3��2���2ӝ�2	3�%?3K3*3O��3U�o3J3�N�2a�P3�3�3�(&3SN�2��73S��2{�3�&3�B3D,3ޙ3�C�2�^�2�"?3JwO3��
3%W>3�w:3���2��-32՘36�.3R�2�E�2
�3��&3"�3`3�d3h=3j��2 ��3�93!_
3��2}��3��Q3ǰO3��g3�(L3Bv3ѳ73a73�LZ3�(3݌k3vOF3�\ 3���2�N3s~3�Ac3��3�h3b<3�3E��3ܝ3�[�2��T3�Y�3:� 3�1H3^�X3��3jD3S�E3��3���2`Kp3���3��:3��U3B� 3�I3�Gb3�3u�H3&�2乎3��3�m3�?3���2�q3��3`O3|�3g�|3��3_3� J3+�_3r/3
\�3;�Z3�s>3#�83�l)33 3��f3e�2���2K� 3�3qhv3x�C3k�	3q3�g�2��3�*3o��2�h/3�j�2��2���2yH"3{��2�$30�3�l�3-?3w33��]3�6D3P�3��S3l��2S�3@�3�Px3�3�B3;3za3��3ܱ3�y3"G3''C3V�53S�&3_�3��3��2܃3��3�O3h�U3C�O3F��2?�3� 3j3�K3XG3K0u3@=�3EqE3��3^�3G6Q3�)3b�m3U23+�o3�n3S�3m�-3F"d3��03�o33��33jn�3�d�2�!3�]b3�?3>�D3�3%B3���2T�k3sd3B�38�!3dD3�Ц2��s3��'3Ъ<3��c3j��2�
b3�T3��'3f)F3���2qm83Qֈ3���2x_"3�kd3}�?3׭3Z�3EL33�(�3O��2z��3[��2�S3ًJ3یR3[��2+3��n3�c3�73A��3���3�iH3���2��&3 3��23dq73'tL39&�3��3�u3	`j3��3)@3?�
4^�<3��S3<�G3.Y�3m�C3��W3Dn3�޳2ʨ
3�OD3|N3��S3�L�2L433,53��2�~�3j��2��3��
3ԶR3�W�2�D3Ї�2X��3޼63��83E�3h=3�3��P3E�
3�a3c3���3$��3ۮ!3ő�2zs�3��/3�	3��,3�3�F�33R,3��_3$3�lK3Q�b3���3��S3E<~3��3Y�7333�`k3��3J�2 �F3���3
!P32>�2^>3Zw<3wO�2��3��'3��2�G�2��E3�]�3�&3?�W3���2�m3-%3��2��3.vR3��3i-Q3��3e�J3�403�B 4�U>3"�j3� 3ꕀ3��3f|3|�Z3jV3��t3��2
�3@�K3R�3���2v4��H3��3b��2�A3�3�/31�Q3yo$3��@3�U�3���3~B3��2 �*3��x3`A3'�23���2r��3P��2���3`�83_r&3�k�2��3��2iG3�4�3J�\3-��2��2jhK3��3	�3�F�3)�E3�t=3w�2��A3�EC3�Ч2��3+��2	A�2�F�2�K_3`�x3-�u3�W3�)�3�2G3>�r3�[ 3?��3�L3ڗ{3j��3��`3l��3�{�3N�3��q3D.,3\��3�"3��3ZV�3�ֆ3,Z�3��3���3�e3(Ϟ3��b3�I44$D�31+�3Q��3G��3�AL3�8�3�r�3;�3㾿3���3<�3)��3�� 3�	;3��3�V3 �3Z��3��3&�T3h��3��3���3�w$3�]�3�'@3O�3k13+��3��2��83��3p@'3Q�3�4S_�3}�^3�a3kݺ3�Q�3��J3�_�3M;3M��3G=3�L�3yx3��3�f3���3bÑ3R�3�mQ3�3���2��o3@��3�E�2��3*�3���3���3�_3�[3��4��3:=�3�3��3d3���3R1�3��I3�e3��3��3�;I3Bw�3�	�3�h3n��3�Ҕ3�>?3�P�3��3�=�3'�3���3D'u3��Q3�c�3Uj�3j�.3�T�38�G3��3#3�#b3h&�3hKU4"�3���3�My3���3�L�3֗3Pa�3�X3pQ�3?L�3]4�x3JT3��4M��3&p63L�3��P3)j�3�3�;�3L`v3f�3�53�ԝ3%/�3�=�3�*R3�P�3���3���3rz3��>3�0�3�w�3���3��3�M.3�	L3r3��\3Z�30�3�`�3+o3��3��3(L\3�
03�G$4�@�2m�3[��3�M43��B3��]3ya3A�o3�5�3N}�3�m�3�3P�3��3>�>3{�43���3T%�3�v�3�q3ݒ�3"��3S d3�ʻ3%� 4s�3
�m3Y�3|߲3�93#�_3i��3��P3�$�3�>4֧�34ȍ3n�3Rh�3kN�3L�e3���3.73o�33;C3 �l3)F3?z�3�Ø3�$;4�m3y��3SE3��43�)�3��I3��3y_/3���34�n�3�O�3O��2�Ps3tcs3�V�3��3�t3U��3c3vq�3���3���3���2���3P�3��3:\S3�*�3GB3q�3��m3��L3�k'3}8�3��q3A˝3�=.3���3RZ�2R|�2I�D3��Z3�G3p�3�te37W3PP63�+3�q�3�% 3�Za3��13d�3���2_}�3j=�3�A�3)z�3g.�3W�S3}�032 �2+'�3��N3�/K3�B3���3��o3�0<3�3��<3gX�3�a3���3�23��)3y�=3a�a3���21o53lm�3�3��35�3~U3bf$3�)3��t3e�3K�3��3�=!3���3�.�2�:�3#8"3jՀ3���2nV�3
�W3�v3��Z3�%3��(3�u|3>[R37)3�3=�3v�3e�2/��2��e3Q��3�43�_3Q$3�J&3]��2�)�3�� 3 "3��3��3�3*03LN3�F3�(13lo3C?3��3\oi3?��3�=3&ٓ3ǰ 3� a3*cw3�p@3�=k3���2�%3(:3�Ր3v.r3j��2�#)3�ٕ3��B3�O~3r3��U3�3�)�3S�3���2A3��3W�s3�_�3���2Q�)3�,�3ǈ�2�L3�,33K_�3R�h3<-3���2�nC3��2l��3�xY3p�53�I*3�c3?9R3Ź63��3KM3)c3���3
�3p�I3���2>��3y�3j�2��3H<�2-�}3t3:�3�-3�93�K3?tX36E3��3�C&3�#33[M3m��3@��2Z��2�}R3���3�u�3x�3�+�2�?s3��&3��.3�U�3���2�Kg3>0-3�	�38T�2��03U�63�w�3�3�wJ319|3=�-3��/3)�43i�I3H�[3bc:33,�3�8]3MA73b��2�Ec3Ik(37�3)�K3!3�&23�?3�[�3�3�3�j93�48k�2�n3��3aq�2R�3�lB3ĐT3�"3u��3В3��3Fv>3�<�2'A3fo3T""3�vB3U|�2�\3ވ�2�{3.;J3��t3�1(3��3t��2�23"h3�.3<I�2(�,3��3T�43�� 3���3k�V3�o3F�C3l�v3պ@3{�2N3��O3��83��2���3��.3�;�3��2v�3�]P3�eU3��3�\,3�3Y{V3�T�3�U3#�c3���3�ӣ3V3	g�2�hm3��U3^�U3�U3���2&O�3 z3�y3~�53�L
3f�2��3j�2YkM3a�3�^3�̹2|}%3�@3��2:_E3ċ�33X3�&3(�25�3��k3���2�o83[7�2a!<3���2�32�3��Q3g�3���3�o�2�P3B�A3��z3��2R*3�2g3���2��<3�A�3,�3��;3n�2�83�13��2�= 3co�2ٟV3�)3()l3˟/3�YL3ĺ�2[:�3��3n3��3>��2w�!3�j
3��39�_2:O3�}f3a_3�73˶3�x�2�
t3ֺj2�)3ǔ�2�c3E��2���3�+32�32�B3�J�3�_�2� A3�k 3n�3��3��3�>s3�g�2�3��3S��3?�3tV3�Z3?3v�3�QV3��24AX3Q23^Am3� 3��!3���2���3�3qM+3�N3Y>�21/�2��3-�#3��28�U3�9�3OL3?�3m�2F`.3k�n3��3�m�2�73��83��2bP�3K%3_37k�29ޣ3n}*3��$3#�V3�H3�B(3�33�(%36�23��J3$�38�3�2�2��32j�2�Y�2��j3g�3ùN3F 3=�P3��'30� 3v3+�3`�3��&3!#3 �r3T��2b(3f(13�߉2k$f3F�3��I3m,3��3�� 3��W3�F3�V�2D3��3��2�ʛ36�2��2ǣ�2�.�3l��2��-3��3�0�2�:33��3~�f3 "�2JdU3���3,3Ғ<3��2��03)2;3��33��*3�T�2�]z3&��2�k�3j�-3�ޟ3��>3���3��F3>�
3��U3S�3k`�2X�3m-3)�-3̐/3T��3j3��3Gl.3!��3�S3g"�2EHR3�Ve3J5o30�2��3�&3�	>3��t3>��3�?�3�qx3�ɐ33W93�D3��u3Pp3s=�3*c;3'[�3!�3�l3�A3k3^3�M3\`�3�;7335D3�xY3��~3���3y�U3�yU3p��3�t3�mg3J�33g��3I�3��.3s$�3K��2m�C3,(4�;{3x�q3��2B��3+�3��Y3G��3�J73��n3�3X@�30�3���3��3�3��?3�X$3�[3�
j3!�)3�{w3rR�3�=3�H3���3	��3Pqy3<y3h��3�H3��3�,�3{M32��38�$3<�m3@GV3,ć3|�Y3���3�h13~�=3��V3��G3�4b3*��3��O3iB3��W3�=�3�_k3N�e3�I�2�w3�yH3s/*3S�3H

3՟3~�3��h3WX3�J�3j��3:��3��v3h�H3L�n3EMt3�?3��l3��3'�/3T8^3�3IW�3�{3w;`3j;3H�g3�3�y3�=L3/r�3>�=38�S3�O@3�)O3��3��4�c[3��C3��3��53���2�=3�u�3��3fVr3���3�~�3��3�0!3%�3W�E3��P3�Ob3.��2�Ƈ3�k)3�J�3g�)3 �t3�N�3ݝ�3L�2y#a3Y�3XX�3��23�(�3ç�3���2�.3E�3~�N3@73+�"3nŒ3��3�a3�3[��2Xѕ3�WN3-�3O�*3��*3�V3\o�3�(N3�w�3�tw3=�3�,3y�!3���3=#3o3#t�3��3�jb3�13�Y�3���3Q3~�k3��&3${B3H>3���3�rT3�8+3��P3Ǐ�3E8U3�l3�u3en3r|_3���3em3�=3՛R3�?�3�đ3F��3()
3!��3�3#03���3�*W3�)�3�!3�t 4�u/3��r3�T3FW3Hw3o��3�<3�}63r�3�Y�3ܺ�3ބ�3�Vw3��3�Gz3��3)3�>�3ҧ�3?vS3�[3F��3I@k3#�3�λ3.�y3�p�3�P3��
4	jk32O`3PV^3�J3.Kn3��a3PR�3/�3`�3��3~AF3�D�34^3IR�3$h�3Z��3�s+3�^�3'�Y3��63f�{3$��3��N3�iI3���3y��2�nB3c��3���3F�3Jm38�3e�3f`93һ�3�~3���2�O�2��3��J3b�3�XT3�G&3l�B3�3��3��j36�m3w�`3)߷3��$3�CC3%I3+��3�rI3��K3��~3�Y3(�f3ed�3b3S	13�C�2k3�gT3��O3��-3�c[3.�3��c3sK�3��l3��3�jY3���3ż�33B/3�h�3õ�3\ �3��3p̛3��3yt�3똠3���3���3<�#3�Ӫ3z~�3,;3�Ck3�Ɠ3���3W�3h�3��s3�'234AQ3�X�3�A}3��E3���3�6S3��&3n$�3v\�3�3<��3z��3��3&�s3_��2�P�3LG�3�3O>v3��2�JN3��3��k3��R3`4337P3�#�3���2�#�2nK3ˁj3mh$3�j�3%5�3�	3ఁ38��3���3-��3K�*3|��3;�83��!3��m3�5Z3�\3f�`3��4�`3:�x3h�_3%�4WI3Ww3�43�3>�3� �3Ȯ3� -3�3��3�i3�L3|�3bl�3��l3x-3.˘3�h3��3s$3�1�3X�32�38��3�2 4ۍf3�_�3pP|3D43t�3UV3v2P3�p�2��3F4�ݡ3~�t3���3���3�ˌ3��p3�#3��O3O73|&3�@4�3K�93���2?�3�W3Ds=3=��3�̧3�_�2�.+3{Z3X�3)r�3���3��3g\�3�Y�2^��3u�3#63 I3݇3��-3��3��3��^3��[3�T�2��c3�!83sYx3'�3Ȁ�3�3�a%3��:3v��2,'3&��3��3��M3��%3�s3��u3�j39ǳ2T�r3-es3}�2�ޖ32!@3GB3֯3��3�a3��\3�LN34�]3�3e�%3@�J3�T3�-3�� 3ǁj3Ƿi3�L3��3��3�3N�93B�3��43Q<,3�t3�3Fah3%��2__�3^xt3���3�e#3j��3��3��u3��63�lK3�(�2ħ�3]��3��f3=�2I=3�;3Z�*3�I3z 3��Q3M�2�ő3��3:B13"�=3j��3G�53�ye3E�m3�q63tm3��~3p#3���2��@3!�3G�^3]QJ3�3��J3m�[3+J�23��2�A�3�03��3?l;3+%3g03E[�3���2wB3���2�F53�O38Ѝ3��a3Z��2��2$�3�8�3͘o3��2*�03�aI3�K3U�{3}h�2��3� :3I(F3]�2�3tv83���3��T3��2�*�2ޠZ3jJK3��.3R�O3!�2�3�ܚ3wdn3�-J3+TE3��I3��13T-3�Ύ3+	3��33ï-3)|T3��M3���2(:�2W��3��2m3�2�2�|3��-3q873�k3�E<37`3;�3+*_3<|�2�2�2�X3 i3�>�2|53QK�27�3/�3	d�3��63lj3ǥ 3�Ñ3���28� 3	�$33#3���2�3�o)3���2�E3BD 4�i�2��d3b��2,a�3&3���2}sp3�D�2��U3�^�2R�3�E3�m 3�q�24p�3��3ך+3�i�3�c'3���2��3(�`3\��2C'3�{3��r3���3;��2S�3F[3�2x`3��35X�3^33�b3$��2R,3H��2j�3H�(3Q�.3w�3F�=38��2���2	�3��29{3�X3@�3�E-3��3׹�3 L3�Q38�*3&L3��3a3�3I��2�\_3��2�݄35@3�3I'3,�3���2@{3w3r%3�@3�63*a3M�3��2�3��3�3O3�DW3�3C-3P�*3j�e3>'3�$3�Z3r�*3� 3�_�2��J3*�2�у37�3� 3��J3F�p3sJ3�� 3}ǉ2As53N��2俴2�Z�3� 38CG3��3�N3)3�3+�3���3�3��3+�2hx:3�K�2��23�r3*3��[3 �X3�&`3�1$3���2�Im3��3��3��3)��2�gQ3���2�@3`��2wu3k��2� 4�,3�'F3x�23<�2H��2��G31�3{��2:}_3gY�3�k�2���2j߰2���2�d3q�24@3de%3ui�2��2&
23y�!3���20^k2�F�3��2F�'3�=_3�3��2��2TD3���2AQ3_U3�x�3��K3FN�2�O3۷A3諘2|1B35��2�_�2mA3!��3g��2���2lN3�Ÿ3�G3Nk3�3��31ݹ2+i3�^�2��2��93�a3�l�3▇3��73�3�9
3 P3��43���2�ֆ3#��2j�3�3]��2��3(�4Z(3F'3��?3Ѳ03�ˎ2��2w3��3�� 3�r3;OI3q�3�2D�3�?3pS)3QE�28A�2��3!��2�D)3�2l�3���2��3n��2���2bA�2(��2@�2��Q3l�@3U�3P:3�b�3��>3t�3R�2�kB3���2���2��33�z3�3���2RI.3V��2�2X�2�H�3߹,3>7]3��43rL3E�2��3��3�R�2f<3|{b3x�P3�43-��2c�A3�_!3s�3{'3��3x�3So3h��3�� 3B� 3^�2���3�>�2�13�+�2�J2�j�2���2�Eo3A��2�7(3SP3�^3(�3Ό�2�n3�R3���29�3���2��>3��2�]3�z3�{�3*��2Y��3��2�pY3��3u(?3׽�2�d3��#3��2��3���3��h3�BF3h�	3�\3PG�2Ȝ�2˛$3SJ3�F3X3c$�3I�~3��3t13v��3˝�2o�l3��>3�K63ʢ2��83/�F3q�#3Vf�2$�3Ѣ;3\WD3�i�2��3P>3G� 3R�3�s'37E3Ty3��3V�33q'3�It3���3�\>3�38q3dgu3!Y3Qo33��U3v�2�j3X�3��K3:d.3on3��\3v��2�%3�i3̒3�@3�;3:��3��V3��u3�V3�ʓ3�3b�3t�23K�`3�3�_3��	3<�2p�3[��3��g3�[U3z# 3�I36�u3J��2���3kt3_�i3�� 3��3-%73_y,3�l3~η3hK3363�ѭ2;�H3U�@3φD3J�H3�U�2��Q3��n3�_3Jm33��2�l�3C53L��2�L3 �3�z3M$J3���3]#l3h�3޴3-��3�3UA3\[k3*<3B�13#F3t��3W�3��3��T3��3��@3^�23f�e3��m3�3lO�2M�O3�D�3�B3�P3ddF3Bo3H�D3��3H��2��'3xK�2�)33|3���3��Q3@(�3A~�3��4�M�3'�_3�3�F�3FY3/6@3
�E3�)�3i��3M7k3��38\3�Pt3C��3�64G�93^ڄ3y�63�`3+�C3�=3��~3��2�DZ3y�3���3� J3�3��A3�F3_�2{#�3�23��m3v�:3,p�3�t
3c�2��X3���3�j"3c�;3*�3�$3��13�"3�@3�G�2u�"3c��3w�3�}l3�
3��3���3���2dE53�93_�[3��*3��3N3��3�F~3�`�3H�=3!�M3��3y<G3�V�2%�;3��*3�H3���3"��3W�C3OA�2��2Ĉb3�_3�*�3��35t�2�H3�3�x3Ĥ�3u�3�N�3/�?4�b�3�ž3�z}3�]�3ۖ03�PH3#�3��D3q�l3��37��3+�j3��{3n��3��3�>H3�4w3o5�3���3PP3�E�3̴s3�kB3ngC3�f�3��3���3?��3���3Dx3-x93b]o3�Ԡ3�>O3��3�G�3umV3]"W3��3/�3��n3�q3P�x3{�^3�n:3���3Ž3�}y3�Z�3�4�T=3=8�3�S�3H.�3d��3�ͤ3��3	R35K3f�3\�3���3OyD3� �3�+�3x�A3Es�3BN3���3� �3���3�?{3A��3��C3ֈ�3��K32�l3���3�!�3| 3U!+3�>�3t�3h�3D��3��3���3qM3%�3Mjh3UU�3~1�3��^3��3\Kd3��3ȏ�3�2{3�43�4��g3U{3���3i�3�k�36cP3�]3x�L3�[L3d�3���3�30aF3�	�3���3��33n>�3!3e�3_hA3��3�@3�G�3�+h3�_*4�̆37"�3��A3Iw3�*E3n��3��3�#3�GU3�8�3�4^�3��=3a�W33��3��_3$ǥ3(\X3��3��|3$C�3ΪC3��q3@�3��Y4c��3�aX3�@�3�,*3�T�32g\3H��3m��2���3W��3
6�3�S3*$\3�V�3Z��3`h�3{�.3�cV3� �3��K3Z�3⹇3n3߳3��4Ą3)��3���3�H`3��r3^��3�oF3�W�3Ӆ�3to�3���3W�3;�H3W~d3d193	�Y3�xh3/o�2KL3��L3dX�3�Ľ3G�3�wm3�f�4��3�t�3���3��3OMY3z�s3��3�13A�3B��3>��3�R3��3?�3�˶3�`f3ƅN3ϚI3���3Z�k3̓�3��l3��"3�p�3[�4"��3D��3˾[3��@3*��3��3$�3��2���3�y�3�'�3��3N�3 �r3�w3ӯ3(8�3�@3�*�3���3��3���3"!�3�J?31��3�3H��3í$3�Z3���2E�b3�X3� 
3��;3�ǵ3��3�G�3��73,�3f�'3_{A3�;3�0h3�ޘ3j��2�\�3TO3��3�=3ӓ3�13�G3��_3t܊3,W3<3���3 �D32m3���3�Ϥ3���3�_3��k3�+�3�83��H3���3��3]�3�}�3��3�3���2�d�3|�.3�f\3 ��2s>i3
63$�i3�n�3HqY3�"d3�Q36��3(%Z3zа2��3t�C3�q3T@3��3���3�3��Z33N�2a�D3�r^3SJ4"3/',3�k,3g��3n��2x�Q3U�3��2�bH3�T�3��G3W�$3U 3G?3��y3�z3@��3#d3�R�3}�d3]�s3�j3ވ�2%��2���3�/3��3�33���2cS�3��3-�3�_63)�.3C��3�\3���397�2jX�37:�35}3م�3��3��o30�H3��Y3
_�3�/3�aI30_�3�,3L��3�X3�43��C3�p3?$�3��3��o3���3(K�3ב�2�n�2ᣕ3]�W31�?3LR�3o�13q�3�g�2�$[3(^e3�/d3P/3�O24J3�2�vN3�3 �O3uD3a�3��3κ3�`U3�r�3��3J�Z3�
3�ʮ3�3��2�9�3E�$3�;�3��3�w�3\�43��3�a3�N	4C<A3�u?3�H3��23�03՚_31�3���2	o3K��3h�r3a�l3�X�2�1�32ӕ3��)3�c�3�/3�Nq3�	�2��3��;3}O3�fA3���3�B\3;{�3}B�3���3pB_3
33�3^x3K�3�V�3s"�3�L3��3�L3.��3��S3�χ3?�73��3:3���3v\63N�
3X��2�4>4O4I33�x3�c3�=�3�3�Y&3�^=3Q�3�[3��3��3��3
��2v�3a|3�`E3�F�3�!3��}3NN>3��3{4=39�3��43\ٺ3��~37�3� J3�g3.�J30�3h�H3J�J3��I3�a�3ؐw3��3K3�4��$3���2$�P3y�r3�|f3�d(3�u4ϓ�3��3��X3>3
4G�g3��33.+3�g~3cb�3�?�3"4�3�3�rZ3x�
4N��3#��3�2j3ϼ�3lX�3�R3�6�31[3��3�X3B��3=�3I��3��3�34A�\3wߚ3:ؕ37�3s�Y3�S3]MX3/]`3�=N3&4��3���3���2(�3O�c3���3�D3��^3i��3��3fu�3|C3��4҆>3
�<4!�f3*�3x��31�3��	3��X3�<�3��V3~ϔ3�-4y�3H7�3��p3���3x�3��W3ҍ�3�(3(B�3�!{3���3"�!3B�L3��3 ��3`�c3+�i3HVu3��3	d3�Ȏ3$s�3� 3��3#��3���3S"�3)�e3ᓳ3���3�6|3�<K3�nE3h�H35l3�]�3vJ�3[=�3!�f3�&�3�c3O�3��x3%=3��3S��3�$�3=,33E��3���3g�4�G�3$�3ߧ�3�ޓ3�s3���3�\63�6�3� w3F
�3-Qc3�� 3��I3��4��3��3��"3���3~�f3d�K3,Z�3�Yk3di�3���3�g3K�x3��3@�3�Dr3�z3|ܺ3�&!3�#�3<&3��h3Ԇ,3��l3XK�3�g�3��g3�7K3�=38�T3W�O3��3zb�3z�3�I3�5�3�b�3�U3�H@3$�3�2�3�03�T�3��3�13�3ܶ�3tjo3��3^LE3�C�3xm�3O�j3T�3'�3'x�3�*3�\�3��_3��}3h�3{��3���3�3B��3���3D$3^m3H(3��V3�i3�f�3�{T3��^3pN3��4%�2�G�31;3�RE3��3��]3L��3%3��3���3�o�3"�3��3�/�3��3�3�2A"�3�93T��3wa3���3.�K3���3��D3"�3�{03�[�3�3Hk53'�2�-3A�3�F3�|3���3֔3��>3jXK3Y�P3A<O3�f3�C3Um#3��3թ�2���3�q3+$�32��3��3�vS3$<3��3;Qr3��"3VH3��Y3���2��A31��3p��3�Ќ3��2>e�3�KM3��2{b�2y.3�	�3
u3�S�3���33�^3y�2�>�3e<B3��n3�B3�҉33j_3|3(3�$�3T�3�63�C�3+L�3�a3:�2�.�3��N3$� 3�X3*,30w3���2N֖3�O/3Ln�3�L�3nt4��"3�S:3:��3q�E3oX3�3��3~��2�*�3dm�3�n�3T�z3Y#3��q3�)~3�M3??�3�^�2���3w��3�Ε3~3��3eL;3Ϋ�3  r3�M3�F�3>�`3��r3�Z�3@͒3�	30ݏ3W��3�`�3m!3��2��3��J3l�C3S��3�7�25��3��03�bs3/&A3�v3��3Ga�3M\3D�3δ3W��2��3 �3xz�3�w�23"3&��3uv�3�T83T]3�Cg3��z3��3s�~3�3�m�3�M3�T�3��@3�e3!��3l��3�,(3WƜ39^3P�/3��.3��h3<u3��2�B[3���3J~3�3�-	3'�3}�F3�53��P3�Z3I�3���2��3^\3�w3ժ3��3P�Z3�T31�k3E�	3�&U3*�<3�^D3��
3���3��3h�@3�^13�~!3�[�3EC?3UM3X�3}�$3!�3��&3{��3͜3��U3"�_3�~�3���3�D�3���3 B�3���2%:/3�2�3l��2�FH3��3�8�3R��3%�3Hc3V��3�K3�b3�g3K��3�K53��3�Y3¾p3td3��4͖934ٔ3�{3�	3�:36�53�)�3��*3U_[3��3Ev~3P�3��V3J�z3Y%3�8I35��32��2ᯗ3�k3Mϐ3<B=3n|3mu�2z��31^3|�2�n3!�?3�n�2`3��3VoI3Ly3�,�3)yc3� $39�2r�3�=37r3{B3��3�03�53�A83El3wG�35�X3��3>�	3#�3Z:3��3�BH3��g3]3��2:3P?3xD3\�M3�83N�.3~~X36B3�E\3��;3e�
3i3�2483�'3�3U3�d 3�S�3C�3�^G3�%3i�3S23e/3|��3Fb�2M�T3���3`�X325�2�2f3��3|b�2�63��2�;3|D3��K3�93,a&3�3�+�3� 63s3�=43�T�2�� 3���23��3�?3�jx3��3 k+3�u43P?�2CP?3�e3�Z�2q#3RN�2"�3&ɤ2S:t3��3�3�3���3�=3"�3I63^�2+n�2�3W33s|�2?�w3t��33R3�3�u3�3:3��3�n�2ρ-3(�2��23�3+��3�n3�8�26(%3�˦3δ3/q3��03CJ�3��31�S3%�,3���2��3�_i3�{3��3�o�2��>3f!t3iT3�W3���2+�3#m�2��3 r3�3#9�2��3p��2�<�2�3ZU63�j�23�3'!�2ǂ3z[R3.:30�!3+�3���2޾3O��2�3���2�1e3c�3j�3��'3�,3�3���3��2��3�h3��(3��34�3�#3M��2Zg3��I3d�Z3��b3U��2��l36U)3���2g�%3'��2��j3%��2�dj3�aE3�+�2�P�25D�3F�2��"3� 3�m�23��2KU3 H-3>��2�m�3i�3�J�3��@3 ��2�D	3�N3� 3%V[3e@�2p�73�~3�;3\�@3a��2��2���3�c�2_��3ֶ2��?3���2�034h3���2sQ%3x�3/�]3�?3N.�2�W3.�3���2/�p3v��2��I3�3�#;31�)3���3{+3f��3��J3֓,3Ye3by�3G�3�^�3`�3��#3N6<3 �3�rg3�>|3{8P3`j?3�#�3V23��3Dy�3�2^3�/3v��3�E3
��3��b3/�3���30�3!�j3e>3f�73
�>3g�3S�/3^S3�ۭ3�}�3*��3%�Y3�J3gk�3[�s3Մ3��3vH�3|�r3���3��}3��<3�Y]3 ~�3�2(3�?3�=3١�3��F3g�Z3�U�3�3��`3%��3�u�3p�r3}��2\N3݄�3�>�2�с3�'3�a37;3 �3�I/3�r�3�St3�u4֓3�J3]w/3��13gi/3�_�3���3��K3�I3�*�3�з3�q�3�3�3��3���3k&X3���3��g3Θ4K.�3ͤ�3���3��3D�3g�3�bC3�C3�YT3��3�53䝥3�\32�3�r�3
a�3���36q3)�
3�83y.3� 3#�}3'�73�O�3;� 3�$�3J�3;7�3\��3Ȓ4͖3��3_�z3��3�>3Bl3n�3$_C3�5q3�7�3�q3�l�3Q�43"��3j�|3�!3�;�3�Q&3�lv3�a#3�*�3�O3J�u3��3j҉32Q@3��r3��2�;3��h3|�03ؑ�3h�%3�8d3� �3�3_<H34�33�B�3��A3Y0L3֕^3�.3��;3�wn3d>�3z3*ST3��3#e�3��<3I��3f3-3�o3Vř3}7�3��N3��^3:�3��N3�
p3<�2͔3�q3��O38'�3���2��3��]3UO�3�W`3kE33�3�4?wU3u�3��o3��3^�3�Y13h�K3F�3��3��P3]j�3_^3��3�0�3ae3��3��-3pt3��31b)3�-�3ӏO30p�2~�23D<�3�L3��,3�K�3�`j3�3��F3��3�l3�qE35�w3;a�3rN_3�(38�53��3�?73w��3^3lvI3�,3 w�3��f3��H2l=�2i��2I�327��2p��2��3���2��2��2Ԛ�2��]2��2E��2�S�2|�2�F�2]��2+Q62��2�Æ2ǥ21�2�2���2~e�2��2��3�ۿ2sA�2�c�2��2$'�2��2���2._�2�5�2V��2@��2g��2��F2��2Z�2%��2��2�	�2gf�2b�2�w�2D;�2��o2u�2�31G�2ֱ�2�d�2v֧2��^2�i�2�>�2�Vv2�6�2Wl+3t��2s;2��o2Q��2�J�2O12@��2E�2q�2��S2���2���2���2���2M��3$�2_U�2�q�2&��2Lv�2̦�2ʧ�2|rQ2�_�2�73]W20�2�52��2��2��2�[o2��2���2�C�29t�2�	�2bA2�J2*iw3)�2�3�2��2*��2�.�2v�2^C�2� L2�2�43�ї2!Ϣ2j�62�U�2l8�2�2���2�o2��2��@2c23�q�2뱎2@gG2(�3n�2���2	��2)�p2��I2���2��2F�&2�
�2���2�a�2���2G52��m2^��2�J2�z2pZb2
� 3
�F2|�n2,��2�w2�Z2A�2���2H�2�ܖ2�l�2��2��3���2!!�2��2g��2U�2e��2�'d2پ�21�2aQ�2}��2�K2*x$3�ʛ2��2���2z82���2HxO3�Q^2�$�2�-�2G�n2ڝ42���2v��2��2+�2��3��2��2c�2ke�2不2#��2���2�)�1�2�k2���2���2r��2�j�2'It3X�2�\�2F�3��2��2,v�2���2{�G2��3A}�2Ps�2]a�2O,�2D�2��{2�J�2}P�2��2�p3Y�B2���21��2��D2�;2�?3f!E2��g2�-�2�|2��Q2QB�2F��2�32��23��2T&n2Y��1�"�2�f2�x2�v�2�S�1�2DI&2^��2���2�K�35��3<2�3eTR3U��3hD3
��3�3z-N3p�l3닎3�=�32�35h�3��K3��Z3Fh�3G�3�3)�S3v�!3{�Z3ڿ�3��4�rc3'q23�H3���3�jV3j,i3,�q3+�R3�F3�T�3I#�3�)3��3r�3��3��3X��2	��3Q�a3�$�2R�,3pq+3k�s3
�V3J҆3Pѝ3B�3�8d39]�3l9�3��3n�3��3��R3��>3"h�3���27�^3���3(�3D3�z.3��3��V3M{�3i��3P�2O^�3S՝3�]x3o�13��{3f�13�4.�O3�y3�c�3u�3{n3�҂3S�x3�I3�53r�4nk�3E73�*�2��13]f�3B�k3� �3�H�2~�W3�WF3�ϙ3=�3�wZ3^�3�Q�3Tف3�i*3��3m�}3h4H3�Ha3+��3rQA3��23�$�3 [b3<�d3��35�3�ӡ3�b3�C3!:3���3S)3���3�A,3��135��3E��3��.3�H3�H3(�?3�ʈ3���3��3bDv3MP�3��3�Oi3�4�3H��2Ԋ3|��3�	H3Ip�3��03�A�3�A3 �/3v�3��'3=_�2K4��3�f3��3{^o3�#�3��3��3�i3��Q3�Y�3��H3<b�3�13T�v3�3h�~3�ؘ3�$#3�"s3�rk3�/�3
YB3��93��|3��3�y3���3k�2���3�@3|E|3i��3��3dE3��3�C�3���3^_3�`3[:�2�f3gX�3xy3��2��	3.U4e3V�+3 �M3���3��;3\0�3�U3�"3F�3�Օ3Q��3#�@3���3o�3�"�3�z30��2�M�3H<A3��;3p�3l�'3v��3�13�u�3�c3��3l]�2V��3�_3���3���3��S3I�S3�n3�x�3�t3���3��3�
4��3�u<3�)O3`H�3�}93���3�,3[.�3��#3I��3���3�I30\t2n�3{�3l�B3��2�� 3��3IoI3P'3��+3J��2���3�v�3˻M33�2�kb3AK3T��2G��3f�2S�3T�2�m�3�63=�[3c�2FO�3^3�%3�5)3�03�U#3�-L3qqG3'� 3&!3�^34�3.i3m3��.3� 3k
�2��:3�la3�3��2��>3ӓS3=A3`��2��;3b@3��^33��a3'��2|��2r�M3�Sd2]�#3�R�3�13�s�2cɞ2j[�3b�/3�O�2 �Z31��219,3�3Ɵ=3>R03��/3p��2���3���2�>3:	3%�3(�2�B3�|R3��,3]��2��3H�}3��2�O�2���2E�(3W��25��2B��2�.3	��2]3�J�2a*3�7�2�
�3AZ�2`or3Bm3�F3�;
3.)3�3�+�2�3r�3�B�3��3�~�2g3�3c�2xR3!�3��u3v	�2�(�3 +3�>3�3��s3h�F3�O3,30�3�23
r 3�j3��3�3/Z�3��3���2��2�s3�MH3?��2z�S3i	�2D�3�K�2�03�l�2�?&3}��2�׬3�+�2�W3���2�3z��2�3�3��2��
3��?3�O34�=3(��2��83�q3���2�
3IE�22�
3=�V3A�N3�3Wf3]�33��3T�3n�"3��I3�h3b*3�>3L3�2��%3�ۀ3�D3t�D3�e�2p3��3э�2�03�=�2~kE3!c3��3�K83�#�2=�3�t�3U�3�T3�d3���2Mص2��21C3���25�73G�M3t�L3�.!3��2��43���3��2B�M3�2��23���2�>F3��2�h�2F��28�3J�2�W:3���2��3���2�3�3���2Y33�3�L/3|<3p��2�&U3� 3��3G�p3�Q�2v(3��2أ|3zr3��3�=#3���3��?3O\3�_W3���3�mP3�B3ǈ#3��3|(3G��3��3�3���2�s[3x��3�=3"NQ3MY/3 F3QK33�c�3��L30o�3o�_3�h�3��'3Z�k3��3'��3uÛ3GF�3���3�hV3��/3ŕ�3P�33��3O� 3oȝ3ؚz3NLd3�/363q�^3�|C3\�3ngY3��=3|�3���3Ī$3T>3^�H3T7�3ׇ3jp3IDG3�m*3\HI3�)�3f1V34u]3���2`�O3o��3�3-�3�B%3#/3`8Y3i�3I�3�TV3r�3���3W�93�+;3�y3�E$3F��2�(�3�cq3=�3Վi3T��3(�N3�Y3Ō3u�P3r�=3���2J|.3�)3��3#R
3D��3�3�23��2���3�lg3>3�3:Dr3���3lY?3I�3��x3SBX3�43��3P<�3Z"3�2�hD3��535�3��k3��@3��\3_�3�Q�3��3���2K�3_r4@ad3�H3XK3��w3�Q�2_�3W3�v93`�+3,4]߫39R-3�)�2e�3�3I!3�<3�3�N�3$R73� d3R�3�I3
\�2T�3��)3��o3��3m)=3YT3�Mg3v(/3Sq3��<3(h�3�8R3�	3�I3��^3rnB3`
3"�x3�b43�j63f�3I-�3�G32u:3F�2ow4`13��3ycP3UZ{3��3?$3l�3Z03��37��3�d�3���3��2�1�2�`3[�3{fg3�@A3�x3^��2�]�3�}'3+F7313G��3%�T3�,�2�cP3���2�39ub3dC3��'3I2~3Q�63Ѫ�3�	:3b{�26�33�@;3w�2<e3�5�2z+(3�9:3{d�3fR3��2�3�(�3��2�y36<(3�x@3A�/3��73��]3�H�2��}3=�q3�Jw3�!O3}�-3�x�3���2�q�2p�j3�2��3�&3e<�3)3:/�3��+3(x�3�o�2Р3���2�PC3$�2��3H�33g(�2k;<3�^3��3�*3���2��p3�J3d�u2���2�~+3���2��2��3�)�2��3!�2�h3���2�G�2�3��%3��23�K3�SP3��28m2���3$$�2�W63V�2ǡc3��G3��2�;$3�|3�q�2�3kz3dA�2p<3�:�22�O3�g�2G��2`ߡ2�a3�
3��	3�'3�-�2yf3Ov�2�ل3�1�2��2��3��3��g2͵3�)�2�%d3���2DRD3���2c�Q3FA3�	�3;�3y!�2A��2�u�2]��2Λ�2C�3?=�2�93�i�3��2`x�2�X�2�03�t3�?	3��2��	3Cs�2�N�2Ȉ-3D2�20��2y��2���3=��2�S�2��3-��2�D�2�r�2�<�2��2�
*3~�u3��p3��2/^3 ��3�3p��2�%3-�2&d�2�[�2�[3*�2�w�2�q(3�P3�2�0�2�413��2��x2U��3P�K3�A�2L-#3"&+3��83�3E#�2�X3�&3Cͭ2rE�2�D�2<��2/��28B3��3���2h�2ĵ3/�63>��2a�3w��2&M�2Kg3:�"3.J�2�;.3��34	33&6�2���2�g3��2=h�2�0	3!c�27�_3��2Cg3��2��H37�3��~3��(3��2��2�2I��2��"30Z/3���2��	3��3��<3uZ3uY�2a31=3���21`3W֠2��!3F�2a�J3�+�2H@�2<�2���3��3T�'3p�431�-3
3nYB3�b�2m��2o��2� ^3�Q3���2^��2��3C0r3��2���2�cN2Ĉ13�m�2�#J3�	3j�2���2�є3�1�2e�*3@�3��p3�M2�v�2.U)3?y�2�3wcN3��3��2+�2�%3õ2í�2�+3ӎ�2p,63	��2�A3�3�� 4>a@3la�3���3S�M3�'/3D7B3w``3DsZ3ؘi3Z�3 +G3��4B'�3��3a#3��3�b�3a�j3�ը3}��3�3�+3mE�3i3��3�X3gq4�m3�ƃ3�43�d83}�S3�U3Q~3��3-�3s�4Nv4�o�3��Q3cߖ3�m3RQ*3��A3.B3�F�3��&3��3�pv3;�3�p�3Ĕ4n�3Ue*3
�~3�3s�93�03�3�3B:�38�3欍3ގ�3�y�3�t_3�%�3��3�T�2�	�3s�3c�;3�9`3�J3=�b3NÊ3ex3Y;�3�63
V3@�3�^l3qD�3
�838hN3�\-3	ވ3\�4�[3�O3ob.3|-3�3yog3귤3���2xد3%��2S��3�c3�3Q�3V��3��M3C"B3v9�3��3��|3� �3~3��t3��3���3���3_��3��3�+3!��3;)53A��3A<;3��3�3hN35�3O�732�-3|��3�4~3.�3��3\�z3Қ/3rT3g>3��3�ت3e�3/P�3̟�3�.p3b�3�ѧ3��2�4L3#�>3���3$^�2!��3�Kb3��83݇k3�]R42��3�"W3~�93�Y3�GL3!o�3�$�3�_3 A�3�
�3�*�3=�S3�D83��3s�3Mw&3���3��F3�5�3͝A3���3� �3���2�~3�4f�R33[/3243)bR3�"3���3��3��c3�~�3�2�3N�3�3K3�_G3�Y�3�S�2q��39�>3�H3���3�;�3w�3u�`3@�3F7�3�<�3���2KΈ3��3��w3�~3��D3e�S3$i�3�4,�3P8&3?�3�}3���3�O�3�3��3HlZ3��	3���3�E3�e:3�&a3G�14�93�93�ܒ3��3m�]3fC�3�O�3ǁC3���3���3m��3���3���2��-3�d3
!3���3�A63�	4�7R3x3�31#F3�ڮ3�A�3d�!4��h34(\3� >3c�3�Y/3���3�;�3�zN3�*�3�̿3s
�3w8�3XV3zn�3.$X33�13Q�3�fC3�6�3�XR34T�3A��3贺3.s3dV�3n.3�N3Sߩ3'q32m�3�3���3Ա%3�2F3*��3�Ȃ3���3�k3�:�3�1~3��2�4�3p�3P��3��J3��3�53)P�3�W3
i�3�i?3R�3M��3���3(�A3� �3V�3��!3���394���3��3v�3рL3P�P3'JK3hO�3�g3FE4�g&3��3�Bz3��3�aF3��4� ^3��m3-�z3��U3��3�$T3tV�3{763nIe3w��3��3t§3�`38�3�l�3�3U_�3۩3��y3e� 3S_3�13d�3cl�2��3�$3y:,3�3�m3JL)3�O�39�3���2Lo�3�1 4�/�39��37��2��3���3��>3{y�33US3b�A3�-B3�x�3
G132�+3�ؚ3z@�3m��3��a3}ٖ3�Ȱ3��3�ri3�[�3��J3�.j3�E�3���3m'3��2%�o3ז3u;�3�S3w�3�'�3���3�;�3� M3/t�3��3��3k83���3+��3ތ3�7�31@�3��3@#3�B�3en!40�3��3�N3�4]`}3��k3���3@8|3 �3_fT3H�3
�3���3�@+3��4�e�3��38]�3��3�443�R�3൴3�>3�'�3-Ѱ3��3���3$3\l�3-�p3�j03���3�� 3��3�3ȠV3N53ݗ3x��2[%?4��s3��Q3怚3$v�3�f3�3e��3�(3��3M��30@�3�ю3o�/3�w�3	W3��2��E3��3��3!^h3;҆3�ߛ3�3�v�2�� 4y�>3��m3���3hK�3�
3��)3_��3�.3!��3�A�3��3�\3��3hz3tJ�3c͌3�t3�u3g�3[�.3��3ӇW3`�h3r�3���3�`d3���3�V%3�Ƶ3��2�I�3��?3*K934k[3,��3�V3��P3q�3�Y�3_<73!�&3'5T3E
3yF�3�t3?��3�Ň3��Y3��e3I�4�$^3(�2%��3F��3�
�3�3F�3�A3m a3��3S"�3��l3V.\3�D38u83�S*3�Œ3�d.3��n3"�3�j�3�+3�4=3,�32��3�)3BbF3�H3{Hq3ҙ73�l3Jd�3~,�2ޓ93�w�3-�3�V39��2:G3�Ϗ3l��2�t�3�1X3\��3"5x3 '�3qwa3U��3�ʕ38�3�3��3
f@3���3�Z.3J�3��j3_03	��3%#�3�O�3��N3y'3q��3�q�3�s3aCz3Z�93� �3lF3K�3!�43�mT3%�3�U�3�nI3�)�3nS�3ؑ�3��43��|3x�3Mfs3?|�3��	4���3ŀ^3��3�|h3(�m3�[(3ʦ�3f�'3�`�3�M|3v�3��w3�LW3��a3Z�(4Un3��L3[=3��3bK3�V3�3�3�ҡ3��3��4��P3�1�2E�3��3c,3�,�3�Q�3Hy�3⺚3�*�3}(3s3�}\39*4[�q3@�H3V,w3�zf36e3�/R3�B�3�n3P��3���3��3�)3��3���3.�c3 �K3�q�3׾3gZ�3�23�B�3l�X3!?63��~3��4�]3��{3a�)3�D�3�a"3o�U3�,�3��3=A�35��3L��3���3B��2'A&3雂3�%3�E�3�+�2�BO3�;,3%�3'ӊ3+�V3�Zc3>4�K�3�a�3B�3P	3R�3��C34�3�3J��3@��3�45w�3���2ޡV3�a�3ݧD39��3� �3W��3��3�zy3�3��3I�63;�3��%3�C�3�τ3�S_3+�93�a�3L�3	�"3���3h�3-t�3�f�3,��2��[3�'�3� �3�n�3g3b�/3���2'��3�=P3~׉3[��3,��3uv39��3h��3��4} c3N�3f�i3�H�3��3e4�Q�3ﮚ3?ޕ3�A�3��z3��3���3�Ş3i�3g�h3�o�3v�3��3@��3]�4��3�>�3f��3��39��3[h�3j\�3�J4���3F6�3��-4p��3,h,3��3�0�3E3�v�3`�3	4��3]S�3��3��3'E3�v4�*N32C�3�d3�{�3j��3�-H3�	4s~3z,�3��44��3��3=8S3l|�3�z�3-�h3u��3�23e �3XM3P��3�a�3u�39x3s�4�3<��3���3�+j3f�O3*��3�+�3ɯ�3X��3h�4���3��!4��f3�/�3�C�3��M3eg�3{�g3�U�3��x3Me46�s39*�3�,3��+4Q�3s�|3�3���3�O�3V4/t4�~�3�k�3��
4C��3��3�E�30z�3wL�3 S3���3͆�3���3��3���3���3T��3��3}A4��3s��3�y�37��3gp�3¦3���3�3�'�3�4z�4	��3�V3��3@ �3�G3f�3֟.3���3��<3;��3���3 �3�#Q3�yF4�t3�`3��3'�t3�jS3���3:5�3�D3"�3Ǜ4)f�3>�e3��R3d�s3y�3\-3�3� &3{�3��39�3J�l3Z3�3�ta3��40��3+��35��3��3>F�3I>�3��3��v3��3|�4���3���3I.3sd�3�U�3VQ�39 �3�z3�l�3CDZ3�w�3(�p3ʓ~31�`3R04�u3`�*3�V�3?RD3�'P3���3���3�DG3ʣ3�<�3��3ܧ�3'.{3?��3L<�3)��3^�35S3�^�3��>3�7�3�'�3�M�3L�3�:4���3i�d3pg�3Uz�3��m3;�R3P�3BKF3?k�3=��3簥3��3w�s3�5�3��F3ׅ�3�v�3���2b��32�(3��3
��3o�^3ڍ3a��3��2]�P3:F3)��3q)3�V3��3)�,3�y93:đ3�3Wy3���2Z]a3
�3;T3D�3e�}3<@D3��3���3��f3�6�3r	�2���3���2�K3H��2�L�3�
3�73��\3�73��3�/�3�3(Ǻ2���2�Ƃ3R�2��3��43�M�243�13F��3�3�.$3��3��3s� 3զ�2��3�3`�3��3I�3�'3p�f3G��3xm[3@.3:_�2�$3��53�[3�Y3@/3�҂324�2xS|3\'3Ȓ3��2�8q3�S30�D3��~3\�>3O�@3�U3zU3�3��x3 :�36�K3��93ܧ�2�[3�?L3G��2�� 3��2ށ|3�w�2|N3+l3(-�2�2��33�3Jd�3��G3�\s3:w�2�yB3���2vČ3X�a39A\3�53��3��e3'_�3��2/L.3,/�2@9`3;36�D3���2�f3�$3J�3��A3��3���2��F3�#3L3ؖ[3�D�2쎃3��3��3��.3�H�2��V3 3���2�c3�3"��3�
-3��z3���2�lM3]�3 I�3 ).3EN3¼�2�3�e37�/3'O3+�o3qC�3�4\�}3��"3W��20�`3��3!3�iS3�Z3g6�3$�_3�!I3$m3���2���2���3��!3�3�� 3v�$3{3$�3��f3�w�2��Q3`�3�ȕ3�/3��63��a3�Q3���2�/�30�P3�3��3-0�3T;�2�]834�3�g�37zH3kM�3ⳗ3�~P3���2�E3�D&3P�3��3jN3�ن3+�3z�3FC3�!3ڏ&3�<3N�*3�R3gs3��3"3��23tu�2nZ�3���2͓23"J�2d�;3���2J@43ۚ�3^A�2�pC3p~�3�z3�`V3y��2�+3�
3� 3��13+�3�T3,��2;`83wr13A�3��2��3��3��^3�WL3@ӗ3�Sa35_/3�23�B3�#&31cR3���3�*B3̋�2�z|3]3
-3��93_!�3��3��B3 ��3�l3lΏ3*�3ץ�3BbN3s��3�So3R�53w��3�n3/d3��3o+{3%	�3��3$t�3��%3
�s3nW�3H�2��%3�4}3�?>3.J;3�U�39�3=�l3��3��3��m3�s3)=&3�Gv3V-�2��3��~3\�3)�3F(�3:y�3��S3�[!3Z�h3=0�3E�!3Hni3�.3~'M3��2�3�3q�2oa�3�d�2���3/��3��=3��?3v93\I37�Q3\��3� 3��3}��3�I�3G�3�W3@�3�J3�X)3��O3��K3�d�3R 3���3xH�3Q�+3�X;3���3Ӗo3s$_3~�|3g4a3�q�3���3żH3�N3?�c3��3G�3�8b3&3�53��3;R53.�3�|23g�3r37�3��3>qB3�E3���3�a:3�,e3�f~3�Od3c�3ha3S�-3���2~�3|xK3*J�3lp3f�3�{�3女3�k:3|�73�;^3	E�34��3{�i3�D[3�H`3�Y3'�3��3�"�3&l�3��3Cfi3O{�3TCi3�=3�ja3NR�3b�z3o�3iv3�!�3��3�]A3�|�2m�3*��3��3��{3�=3+�E3�#:3o�3P~3F�a3��P3V>;3C�53B3|38�p3m�&3v�3Xn3��3|u�3��3�2&3�3� 33�Q3���2G[3�*F3P�3f�3�j{3�b23L*�3Y�E3�ڒ3ґ�3��j3e0u3V+3��3u�3�F�3i�3��3V<�3��D3��y3b��33r�c3��(3]�V3?��2h��3���3�2�E�2'��3�3��3k�3R�;3�3G�H3�-s3%U�2Z�^3���3E5�3�QB3-.�2]�3H�23�H3�GU3u"�2#v{3�1+3�^W3��$3�^3ĸ�2�a32�3��3�*3�qE3`'�2`G#3��3��2*��2P�53�
3��%3��2�,3�3>T�2��2S�%3am�2��2�l�3es83	�2��3=(c3�O�2�2�3쿭2DK3���2��3ح�2�e�2�nP3�3���3�ts23~��2r2�2E�3K�3�3r�Q3P�3k03�#3�V3��-3
s�2Iw+3�~3�E3�G�2�O3K�3���2��'3k�<3S�*3oZ3�y�2��03�wA3ܑ�2��3���2��2Ң�2O�25�3_&3e3�� 4aP�2��2�-�2l%�2)��2�~�22#3��2���2�3��G3c�2�z2�1�2V�!3�2�c^2Y�2�Z�2[q�24E3nN�2%�2���2���3�2^%3�G�2�8�2.�!3+k3�>3�_�2Db�2��3�3�-3�.�2�i83�b�2'B�2(�83���2F��2;��2���2�G)37h3���2�d�3�3D�2?�(3�f	3���2t[3��30-�2��2�n3 �A3j��2〨2ew�2B/3b��2�23Qd2�3:�2qY3Ǭ�2D*�2��2:�3��2s��2��2/J3^��2���2��&3�؟2k��2I3i3�.�2�p�2�Q�2���2��2a�2U�w2�V3���2<�N38N�2��3�3��3�$�2��2m*[3e/3�13nL3$3c��2,�3��3��S3�'3���2~B3D��2�}�2��3���2g813w� 3W�3���2,��2F��2e-�3�e�2�3PO3��3G�2x-:3/�2�T�2�ގ3S�3�$3��3�C�2ٞ.3�;3 %3���2ň�2�P 3�>�2��3S�3�G�2zl�2Ϋ3!ѓ2��k2M��2�3{��2�p�2^�u3Q�2��2���3#��2��2��2��:3C+�2-�2�cL3�e�2$�2�B�29�J33Z�2�P�3�s�3l�3m�G3x�3�c3��3�A�2�<3� �3�TZ3�KL3o��3�S^3f��3��3���3��N3yz�2:Y&3�4,3�'53�7�2���3%�43�c�3�}3��3{�3��3q��3���3�A�3��f3֮3���3z�W3��3�9�3�c�3��3B	�3$ވ3��83�%�3�3�U�3d��3g?�3�Θ3䍍3YU3�\�3�͂3��3bf>3](�3�Ώ3��!3�3�wf3yXz3���3E��3/�i3��T3�w3�,�3�3P�P3BW�3\K�3�;�3V��3O-3��3I�3��3�)�2�&3w*�3�43�?3B��3��z3M3_cw3��3��k3��3��30��3�~�3�zQ3�Ys3�@?3X�3��#3@��3�'.3�3�"3��3.k�3��X3�{�3�EB3_�3�-�3�h3�3��3��3�1Z36�l3�3Iƪ3.��3�)3��T3d�3��3�pk3���3�@�3�PR3�P3!��3�33���3]˚3�;3��3MY=3^��3���26�Y3��3�3y&�3H83$�}3�@A3�"34D�3�j3�p�3�� 3�p�3%�Z3�=3�:3.	4��3 �3���3��3�83l՘3� �3R��3�u�3�W 47�3��3\�3��3�GT3��83�3O�F3�׀3O�}3�3�4�3��S3��W3�	47�3li)31�Q3��3��13�b�3�ϔ3�)g34��3uSs3<��31	K3lE3\��3U3)eX3�0q3Q�`3>�3��k3�-�3!�3x�3-63��3K3E3�U3�j�3˿E3=(3^X�3H֛3��B3�,�3���3>e�3��3���2"�B3j��3�&3��3�3@�4.ъ3���3U(y3��R3k3i�3Ac:3�s3"�{3j|�3`Ӟ35�Z3+��3޶	3��
4Ċ�3A�3��o3�j�2�d�3�M�3q�53�#�3$(�3�j3� �2���3��V3�	�3���3eR4��H3�p�3���2��3�)T3T3r$q3�Wj3�_3�X�3��3mm�3��&3
ڝ3�`�3��43S�W3W�U3|P�3h93F�3�63�}�3�3���3#3-�3R��2֞23���2�V3%�f3�]3�5�3�E�3Xf3�w	3��3]�3e�63FQ_3& .3�Q3�.�3me	3�u�3H�3Jx3-�3�^�3��3P<�3e�/3��3��G32p3{\%3�-�3�r3�
�3<��3�G33� �3@l�36�V3�c3Z<w3��`3��3��3��"3ߠ�3���2׿�3��|3�P3+N�3�b�3�3��73J�M3W��2"P3 ��36^39�d3�,�2��\3�n03P�3�R83�y�2NȜ30�3�Ϲ3ab3��[3F 	3�+�3�nq3�;�3f�+3��U3��83^��3òq3�� 3�ex3��3V�3CF�3�43��3��43���2j͡3P�M3'q3N)k3�"�3T
@3V:3P$3	��3�<�2�*g3��3.�Y3y�>3��83\*O3�$3�23@�4���3�-3C=�2�Lv3��3?j�2U�3�r3�#�3��3�U3�;13�VU3��03o|3c%3~R 3T�^30�K3A$K3�{m3��3f23�_�3�#�3�	q3�3W�3��3C��3�fn3�
�3N�3�a3�gC3�`}3�?3k3�Q30��3QI�3��3_3ɉ�2g3*A23���353���3E��3_��3G63���2.,3Ϫp3�A3}�K3�Ok3���3߆,3j��3j5�3��`3	a'3$��3�?3�13J�3zY�368L3��3���2�=3F�V3�3�3�$�3�(S3�d3 z3=��3��3�w3�@+3���3"��2ɵ�3��{3v@3�2��4��3a 3*L�34A3n@!3�^�2�=Z3�1G3E��3@��3�o3/g3���2]3�_3!I�2T�O3�*3Y(3:�2�s�3�'3��48��3��4<��3'�3��l3�pt3rh3k�3FD�3ꫀ3���3{M�3oQ�3�O�3�Q�3qA�3G��3��3��3���3�q�3+�3��3;�V3RW�3�]3=�94�}�3���3�{3���3~DE3D��3h��3m��3Xou3)J4ϵ�3�<�3�^3��3��3N��3)l�3O7�3���33ʔ3s54�F�3Q=�3�973NV4Y�x3��3�]v3Ә�3��3�8�3�2�3�]3�~3"��3pB�3_�E3)t(3�w�3�J�3�-�3���3��53�3~��3gг3m�>3��3J�31F4��z3R8�3<3>x4�3���33!�3��L3?'�3�`4���3�<3�
(3���3���3�`\3��36��3_��3�53��3µ3kf}3S�3��3I��3& 3k̬3ys�3b�~3���3�)�3�g�3<e�3��4�W�3�3��3���3?4�4l3�]�3
Ƨ3���3Il�3��3���3-��3#`U3��3��3#��3޲3���3J�73�j�3�<�3�x]3v��3��4LW�3ɮ�3IAz3�p.4_��3ǔ�3�o�3?��3���3_�3^�3|R�3L��3<Q3���3���3⓬3"�3�̪3���3�<4)��32�3 ��3T�@4xM�3���3�R�3X��3�3���3֑�3�\�3�q�3��n3�4�}3�ǜ3�<�3=44�I3w;�3��3|�3�cy3M�3�]�3_�3��3�Q$4��3-��3�D3���3�%�3	�B3z�3L�z3T�3�%�3�9=4��Q3�x3�k 3A24���3J|4��3�Z3�~�3�=�3�4_�M32��3�&-4K��3ꣻ3��j3?;�3�:4Vߑ3��3�x3�Y�3��3�3��3#"I3T�o3m�W4b��3�n�3�7�35�3�[z3FC�3D��3�*�3Ͻ3](4�]�3�8�3�93���37W�3�P3f��3���3���3A�3Ah 4��3���3r�3Ү�3σ�3�B!3��3��3��2�>w3i�S3�}3�-3X$q3$o;3G��3�YV3z1�3�M~3�/s3��T3�،3�3h3���2:ߦ3�W�3.B3	�|3|�3�03�2�3HMh3��/3��3T�q3�W3/��2.sH3(n�3��T3�R�3���2�H3��D3��Z3A�'3�f3t)43�Q<3�vP3>u3oD�3��&3���35�3�3Ɏ�3�%y3�gG3d�3�̦3�fs3#UF3���3��3$�X3'G�2�e�3.�S3&�3�3�^.3��3���2���3��3�*3�w23��4��3 %3Ċn3_��3*�U3�.o3�k3[<3�n�3Sғ3��3��33��2>��3���3�0b3��*3{3��S3#r03ة�3"l73c�"3U�2�ܧ3}��3)a�2 ��2䥀3��3�$k3��v3Ҟ03g�A3K~�3(�3��3X�K3�Ò31Q3;3��A3� 836�3ΩA3��3Qdo3�p3|3%3�,�3�743�3a3w 3�	D3�tF3�]n3=�e3��2��3��3�z�3U\3�ee3}Z�3��z3M93���3@�y3�n3�#�2W7q3!23�338�*3D�4��P3�$~3��+3��3Q�~3ɃQ3�.T3��j3��q3���3QF�3(kX3�%3��L3;�3���2�k3t3r�w3��t3�L�3���3��S3u�?3���3�Y3�~M35Zf3)߃3Uʷ3�Xg3mU3�E\3b]q3H��3`�3O�\3�3�T_3��\3�$3�߇3A�A35�;30h3��t3	Vl3�nj3��3���3\�33Į�3�̈3��d3��X3��R3��b3۠{3��	3��3��3�3�� 3�H�3�s3��3���3��[3n�3׭3� �3��/3���2��:3��44.�L3/�V3�I�3���3R�}3���3TI�3:�?3PS�3���3�T�3�F�3p�!3p�*3�Q�333_� 3���2(�3 Ё3;��3[�3�3�T�2Hn�38e�2+13�_�2 V3�1�2T/3�3։�2��3+3~��2� 3(L�2�*3O"3�3F3��J3[�13m:�2�CX3R�3s��3�X�3�V�3X_3��;3� �2��@3���2�^3��{3CKs22�03܋R3��	3��3��3��3%��2r��2I��2Q��2�|3��3k�3���2�3cS�28@s3�y�2ɴ3��2G/37`�2z�(3 @3n̸2̧3i�)3���3���2;��2~I*3H�13��2��3A��2j�)3���2�/A3U=3�y3@�3>��3�!�2x23�>�23O�3`F3
�/3��3~:63X�3Gi3&3�U�2��N3	YP3�5�2��U3�:3�f3L�y2ʸn3��2)Uf3�$�2��r3SY3���2��'3n}�2��2��33�Ё3���2��(3/n�3�GC3���2� 3-*f3�Q�2f�2R�3��2�n73P�2q�O3L�,3V��2i��2�3�� 3yg3B�-3���2ϫ�2eS�2^��2��2_R�2�]3a
3f)32H�2/�3 -3��!3�5!3[� 3WE3��3C3kb�2O�!3r�C3/T�3�%3R��2%=�2ෑ3���2�93 �<3�U�2�30�3B�z3���2"�z2��n3"9�2���2<�3p��2b�3+�33�632�3v�2lD/3��N3���2k+3��w3h�.3Չ3���2�V3ڋ�253�dL3Y�3N|3%~�2U*�2�l43}��2l� 3���2�l3��G3j�l3��3�B�2Y!}31�3Y�$3NC3��H3���2�73�3�Q3��3�gV3�[�3��3f�23D03��3n�37��2�_3X�2V��3QY�2'_3-[�2���2t-E2���3�2�;�2#�3֏�2�>�2��2�� 3	A�2�3���2o�M3n�3�#�25�#3<�I3�J�2��21�2��3�ϱ2E�83�J3+��3K2^3�4'�Z3��}3�T+3%�4���3~�3�eQ3��F3�0�3>"4�Ũ3"�[3��03�z�3��|3"X3*"�3n�&3i�3u�3�:�3��~3(��3F�3��.4B�L3���3�i�3�4�3�
�3���3R#�3�ca3�A�3�Z 4�+�3m��3�a�3E/�3P�k3��`3���3��@3��3c��3�4\��3�3U�3!�(4�E�3À�3�I�3�!'3��c3:!�3a7�3W3�,�3gT4[`�3��?3���3Ӑ�3�h�3�\h3G��3��3��Z3&�37��3��3W:�3�Jz3r�4���3f0M3|�3?ҙ3*�p3Z�3���3ǆF3�F�3�X4z$4 n�3Ec834�v3_E�3x��3�3 ܆3�Zm3�-g3�d�3�<G3��?39U=3��3�v3pK�3<)�3�23�9�3$^�3�~4�jn3s��38�3��4��j3��3�l�3��3Z�e3��3�3IǦ3��v3�
4�~�33�3bˍ3�N.4<YX3s�>3�%�3 f-3� }3�L34e�3��&3h��3D�4v4>i�3��:3LF
41��3��3��3T�3o2�3dT=3b
4�G3i)z3�3�3+�I44�3l��3c��3yM�3*�x3��3sV3�Df3?0f3�4	4脏3��T3a�O3�na3�3��c33�3�.3hٷ3�W/3�:�3�b�3�x�3q��3��P4	=�3�FU3q 	4�=�3�`�36
43ꄌ3�3�4�3�=�3�>�3�&�3V4#3�"�3
�3k3S&�3��3dT�3�t�3#�|3\�i3P��3*��3�׋4�S�3P��3�y�3n63�֝3r��3�]4�t�3do�3`4��4�d�3�C3�+�3o[�3gz�3�n3P�[3�4.$&3���3.��3�E�3I�2�;d4⛢3�N{3�ʥ3FY�3��83.h�3��3c83�(|3`B4�K�3Ψ4?ߒ3Yy�3]�}3���3�m�3�я31��3��3,��3�B�3h��3�3 X�3&+	3̲Y3#�3]Ő3J"�2� j3x&3�>3��
3	!�3��/34~83�G�2��=3�5�2�|�2?KG3��.3�@3��2_=�3M3�9)34��2���3�^#3+_N3ɐt3��n3��3�`3��93M�2s�2��3�3�3�:�2��d3Z�T3s�2l�63���2�
"3�)3`�I3Ngx3a	*3D�*3�Z�3E"�2d��2I3!r�2�3��2sf�3��2��@3��3\x3H<3��2Y�X3��@3{'�2�>3�J�2�3?� 3�-U33��2VIr33U.4/�3�-3=�J3�,3�}q3Ê'3ܪ�3��2�F?3�E�3>�z3��;3�3�2��-33"�3�L�20�3��G3��~3�r�2xHx3��3Vz�2q�2��3	�T3�F83���2���2>�A3D3�43��3%�R3�Ҟ3�i3�`}3���2>s23z�3��2A�3R�+3ǲ23� 34�@3�43�Q3�S�2䓖37 �2�2B�3,�?3µ�2{�I3N�{39��2cJ�3�n�3'ܨ3q?-3��C3K83�_k3�c�2.�T3+�3&
13RҐ2�Ѡ3w��3�C3q��2�2�3�3��3X�33�{�2>�"3=%[32�<3�#3yB(3g��3�M@3�3�g�2��3ձ3/ɿ2q
u3��2�3�3��:3A^�3���2^O�2P�2J�3<H3i8�3�.3�c3�O#3OA�2ںW3�3bPP3��|3��3i�43��2��]3��3`�S3�j3�J3�7m3T�2s%d3�X3��h3��f3��3�,3�=33R�G3�3���2�k3�z�2V�3���3��3(-g3���2(3T`R3��3��E3�E3��@3V�3��w3�b;3O��2@��2K��3��T3?,�2�DN3сA33�T3�
3ֽ�2�3+L>3{�3�13��2i�.3WI�2E�3���3TF�22�a3}_�2�]3e�A3��v3x��2��4�C3�C3�2(3�;[3�H)3�(�3Z3m�3:�i3.��3+y3O΄3�jN3#�^3��{3[�3��2�a3K�W3~`3���3�v@3;�3��3�3f��3(�G3�^3 �635�3�u�3�X�3�$3Ќ3��3=��3��_3���2$(3�La3_3�WD3��W3��z35
=3���3v�3�R�3�b�2]�3㏐3>23b�@3$23���2��J3�8�3˼+3��r33N�3v�3�W3|{3*��3��;3�3�b�3ߴ;3�m3�3�<�3��b3�p3��-3��3��3��3zSD3�9a3�y 3�O=3A��3Ud3���3 ��3��j3a�u3�[N3�!G3-�l3WFJ31�/3"�93��3ՆJ3^E�3��e3S��2�:%3��35*3�!3��m3q*3�RU3��3�|3@5P3)ϛ3\��3���3Lt33Ճ3*��3a�b3RI3���32S3�v3���20i	4�DU3�;3�:)3���3/�3/�3msj3lE 3�S43�lA3f�3O3UA3���3�3�h93�3�2\s�3_�3X�3ݔ3�c3�q�3��"3#�3�s!3�>3^NN3��4ȴA3��3:�23�3�#W3QO3z�3��@3Ãk3��3��3��=3�� 3���3�GT3��3�0F3�+D3�P/3�23I�3�ZL3��R3��X3P��3L�3
>�3>�93v3�V3md�3!;�3�3�ɭ31�3�ѫ39!�3�|3�9�3/ױ33A3oq�3�j�2W�3��_3��3�a3��=3}"h3�\�3�b3��k3U��3��3�R3��x3�vj3!B�3�Ǣ3y��3���3B�f3�e,3�O3ϙ3͵�3�!n3��2�F�3�E3��{3h�U3��q3t�83^�3"�V3xv�3�C3��p3��3� D3o�s3��3��3���3���3� T3�P�2�v�3��t3$��3��l3V�2�0�3��'3u49��3�3y�D3X��3o5#3��x3(3�(�3M�&3|�3�<�3�.3+J3xs�3Q�z3�3;3��D3���3s^3!��2�n3ծ53�[3-��2��3�D�3J��3��93E�3g�=3<P3���3-�3�?F3m�`3�m3Xpw3�2_3\��3թ�3MU�3��3�J�3� �3��h3��Z3ՂG3n�s3ە	3��323�Ⱦ3@�F3zd�3)a23E�3 ҈3㶊3F(3��53�3�(3 {L3=�3�(�3�o3��:3k�`3��63�
3�+T3P3��3S�E3��3A;3���3W)3���3��f3�U 3���3�{x3��,3^ń3�`�3�3]�3�3?�3C�[3�S3�c�3� 3 �3��]3��93[R�3 BM3�^�3�*3/Wp3"�i3���3y�3yn�3�Ŏ3!�e3�4Z3�Su3�X!3�J3�(�3�D�3@D�3��73�93�˰3�o�3��p3g�3�Lq3�U�3��p3b�Q3Ig�3��3Z��2Z'�3�<�2���3�3A&:3�P)3e�=3�J}3�93�(�3)-�3-��3��b3i�>3���3��F3�� 3�om3)�M3��:3p_+3���3r13�E3 b3@�3]#3�.3y�d3C�H3��[3ʺ3�=O3�	3�z_3�1�3[��3�J533j�23_�@3C��2��3��3��c3a�73�/�3�@374r3��B3�4�33Z�l3�͟3���3o�3ѩ3��K3H��2[ې3xɖ3�E�3�|�3���2QE,3-J3�!3ե�3��3
 v3͐3���3y�33�793�#+3�,/4��03��'3W0�3$�-3(Ν2c$3�3-z�2�2�3��3�3#s3���2Sm	3�?@3Tj3�]O3�h32�k3$b3��3sn\3 �3��'3�4�k3�;3�MA3l�%3ӂ3>�W3�R\3�/3��L3%�c3�Z�34��3o7�2
6�3k�>3��N3R>�3�/�2��c3|	3���3��3��4qf3/d4�H�3E��3� �3dQ�3o,�3	��3è3v(�3���3��24~]�3�3%ݗ3�R�3�	�3�i3lY3�?"4��3̃s3�N/4+2�3���3d]�3�4���3���3obJ3�@�3�W}3��3?�3E��3 ų3T�4��3iT�34��3�_4��4L�u3��3�{�3�L�3o��3�\F4�F�3 �4-�3|&e4Ǹ�3~��3j�3U��3�U�3�У3�4GL3�3���3]��3s�3R�3�9�34?Np3 �3�C~3zu4��3��3�^l3�K�3Gk�3��4���3_i�3�e�3�+�3n�3���3�^4��3�I�37949�4�	3�j�3���3�|�3�y3N�3�DN3�3d�3:),4�%�3�y�3J��3D4�3>��3�r�3~�3=�3F��3���3���3�ڲ3�4kF�3N{3��N3�M4mw�3�x3���3���3tǌ3�N�3SI4�#�3��4G�3�~4��3�X�3���3N2�3���3�g4?��3�^36	4I�:4r
4j�#4C��3�ޚ32��3�C�3�[%4,݉3��3��3rL4�k�3�63/4v3+�z4�n�3�Z�3j�3�3���3��3 ni36�3��3��&4���30p3�`�3�A3���3A�3g�4[RI3-^�3��n3�4�D�3e�3�x 4��K4B��3'�3/`4Wt3l��3�k�3���3�T�3�;�3!4O�4�{�3|��3�	4�(�3�[�3��44�3��4���3�4i�4Vޅ3�'3��4�3��3}Ҟ3�3�!�3���3m�34�i3�x�3I��3�r4�K4�ʑ3ʈ4��3?�O32}�3���3��54���3L4�B�3ܭ3��23�~4�6�3��3���3B'�3�X�3-�37��3���3P4
�4��4��3y?~3-4���3�¸3���3�y_3ܵ�3xt^3��14?J�3|b�3�83#�,4M�3��3-�]3�u�3�_�3P4^�3�S�31#�3}�3�U�3�4h�V3���36�3�F$3l��3���3}V�3^4m3���3���3G��31&�3I�30;�3��3K�33r�3{��3-��3��4��4��3��4�Q�3‏3h��31l�3$"�3)��2�N�3VZ�3Ƙ�3�ə3e��3���3�}�35�73,,)4!T33Ը�3�M�3��B3���3}�X3ন3\un3�m�3��3�3�3�3|ɕ3M��3DY]3&��3�ׄ3�B�3Ǫ_3V9�3�<�3�)[3$]�3��4�~3�5�3:�3
�32!b3��3K��3�(B3$��3�d*4	"4T�A3� �2�I�3�V4�r{3L�3�sM39٘3��3��3w+.3���3�I4�I04��3;��3-{�3:&�3�3�v�3��3v�^3��3r��3g�3C�o3kJ�3GF�3H'�3�t83#�T3�؇3M��3�,m3z$4+ }3��4��[3U��3�N�3p�3a��3?c�3�<3���3^�^3l~@3�
�3D�4��3|l�3��U3���3��3��3
��3�].3bu3��3��3���3U=m3	�S39v74;�n3xť3�q73�zz35ϛ3���3���3��B3�=�3�F�3Q��3�l3�3��3G��3�^t3���3a�~3ow�3��u3���3K��3�-�3;��3/4�Pl3�>�31�H3U��3h��2��3���3��03��3�!D4�E4x}�3��H3ӷ�3��3Ld3	G�3X3>#�3@}3Xc4pl�3�d3B�3!64�z�3��3�iq3]�`3�]}3j��3A4��D3��3�#4��
4\!�3>�3[&�37rl3�*�3��3g�3�(�3zaP3�,�3ͭ�3n�v3��_3�fI4,�43ŗ3mE�3�C�3i�P3%�3�b�3563Zl4r�d3��3��3R�Z3��3q	�39H3��3��3Il3��3	�3�͖3l�3I��3�zA4�'�3og�3�³3,�3�}3o|4���3��@3�y�3w�3_+�3"�3�^35_4q�3wX�3�4�3�(l3���3�cm3x��3��3c�3��3WX4<��3�a�3K�]3ܻ3�м3�P�3��4��T3��3���3�?4�]4#�?3R44�?�3�ߡ3�[�3�G�3���3E
�3g4���3��3�133+4
��3�q4FD�3��4��3˗3s3�3���3���3QuR4�P�3��3g�(3��3��4ݪ3	$4��3g�4;N3���3�ï3�3�~L3(X?4�(V3XΩ3�K�3KA}3Cj3�6�3�654
�3)��3�4N�3�h�3�K3�4 k�3(	I3�H3��3e��3�Jy3*�3_��3\��3���3�4���3%T�3�s�3ڕ�3W�3�84�V�37��3��3l�b4�j�3*׫3!9�3]��3��3�̃3Ӿ'4a�o3އ�3q=M3�w4[�32P�3}3��$4U�j3P��30��3	X�3n��3�h3�3��23��3�K49B�3s��3>3	��3���3��3�`3~.�3us�3e3?�4���3Jf;3B�3��94�y�3 ��3C��3*��3QO�3��3C�3]L�3��3��3�X�3l9�3&j3~N�3�?r3���3���3��3�G�3�b�3#��3Y��3j��3s�3ő84)j83<L�3h��3��3/3{3E�3q�3�$3{Su3�_�3��3�ؼ3�F3s.�3���3�u3��3 �53�t3��3�/�3��73�3�3bL�3HM4���3���3	�3�S4���3b��3��24�W3NW�3B�)4�׬3m�3uw73�C3`��3VG3�5�3p3��4to�3�1�3�	�3 �O3)�03�4]9�3��3��N3�y,3��375�3Ph�3d
�3/y4,)�3$��3p�3.3[0�3�l+3ăn3��3�՚3i�3�{�3���3�;�3�3ǌ�2�v�3��+3���2.��2��2�2�13)�3��2� 3g�J31�83$[3T`�2��=3F$�2���2�n�2Rh3��w3 ��2_�U3�_�2��^3��3��3d$3��2Ej3�3�2p�2�j3�U3�$�2t�w3qR�3573�3|T2��135�3�ר28V3�4�2;03A��2��h3/L�2�N3u��2��e3���2'3�,03��33S�3�@8343T�2w�2�V33�3�X�2��3��2`�z2��_3_��2ֆ3���2��2�^3��3{3a�3B 3�	3��23?��2<�2��2�J}3)'3瓶3vՠ3ӭ.3�"3��2k13Bq�2N%�2�R3�j3��s3�!3G�&3!�3�M
3�e 3���3�2~�E3i=�2$z�2y�3_�2E�2I��2���2a��3�_53<�2`��2`�3�a3��20�n3VI�2���2��2SU�3���2Q39+G3���3�53~��22�2�p�2p43�>-393]`3���2\e3�sX3Ѳ/3���2�*3�{63TO�2p�2���2 |3���2�G3�T�2�2^�234P�3��3��3�3A�3��2�R3z*3�3�2Y3�[36v"3s�2"|�2g�53��3L�%33q��2)63Ac�2�SP3|]3��?3�t�2\��3��2ү83N��2G��2�p�2i��2-�.3�=33��3Bx3ɽ43(�3��2�*3��t3ѹ 3'�3=r"3�N3�2���33ע2C��2�>�2��3���2�K�2@�	3�;3t#3�T�25�]3�)393ʂ�3��t3�b3Jݱ2D�+3��21/3ӄ3�]D3|�3��2��@3'�
3���2-�2�43t��223��3`�&3�T�2E�<37�.3�n�2�@3���3�#3mB:3�ۤ2m�Z3G��2�,3X�3�v�2�=3==�2�NL3�:�2��3�C�3��3�Rs3��3�3�N]3魴2�S3r��3�3�F13፡3d�;3c�T3�d3I��3i��3$%3��2�13� 3��2��3Y�35v3<�3��3��2�3M�934��3|��2���3��G3�]�2R�O3#�3m43��3��2�>3nD3#�R3�:3��2��3�3Л�3Xq�3��^3ƴ,3J��3Ӽ�2�63��935Q3�f3�yq37j3�_�2��^3i��3�Ԙ39'32�3��23�(3ڴ2 �3�#3�/3��3��3��"3 4�3IA3.�3[�39'Y3'w3���3�N3�-l3�>�3>�?3@6�3O�3��|3$3���2��3�3�j�2��3�?3��f3.!3��f3��3}�3�3O��3�53�	G3 r�3g!73J�$3ת"3n�63���2<�3�3� �301z3A	3��3GW3Z�3m� 3�u43��G3�qa3��3�!@3E3��2O�3g.P3#f3.F$3��3�n�2��3�c3�H3�ex3&�3��\3O 3}�2:��3ro�3ACS3��,3M��2�U#3	C�2��3a�G3��n3}z,3'4_�U3�!3T�3[��2��)3��C3�Zi3e~/3�@3���3���3�}�2��3��3T�=3��P3]�3���2��/3�,+3�9�3�3��"3K�203�3��3g�3{�V3���2Ю!3NW3�'v3Sh)3;K+3��3�В3�8(3�x2/߉3�K�3;�3o�w3.�2��3%�3f��3�^3q�33�QU3���3�D3���3��3U�2"�~3>;3��b3X3���3Gy^3�GN3��q3��R3�t3�I3�.P3O� 3�Z3��^3˺3]�3�d-3�H3x��2���3C]63f>-3�\3)�e3Pc�2��&3�ܝ3.U�2��L3J�4w�u3>ӯ3��38G3�_3u3��l3���2ن�3�3��3\,h3��
3a;k2�D:3���2��3+��2��3��3`�;3��3��3�W�2��U3t�[3)�2�ߦ2X73�$3�D�2B��2��)3�/�2
��2s�[3W�N3Ғ3Ct3�aw3¬)3�|)3��K3�� 3��2�<3@:)3-$3�) 3VL~3�(g3��L3Ml�2NNy3?j�2�H�2@<3�3h53:�3uJ3u��2KN�2e��2���3֤ 3"183ۣ#3��83/^3���2�GX3\I�2O�3�%b3�O&3P��2}�Q2��`3N��2���2�T3;�3�@{3f��2��D3�39�Y3�ro2Rt3!a13�X+36�3��2@X32�\3�<3�(3�Ag3Vh�3G��2km3k�3��43ED$3��2�~3�� 3� �3F��2)tf3�H43���2�z2�.�3�?�2U�2��Y3e~ 3��2�E3C<3:�2H43ab)3�3C��2{��2HB3yl3��2T�83��2z�!3U��2��3:�2Rm�2f~�2���3:$�2ۨ3��3�L�2��2���2� �2Ư�2�r3�Zo3z_3s	a3�k%3�;3^v�3��2&��2��3�3/�3��2D�3�33�w�2�\�3���2��2��2dV39J�2��63Q�B3!�2��03�
�3V@�3��3s�2�3
O�2���25��2I;�2�#I3G�2">23,�v2�J*3B"�2���3�/-3��H3�* 3~Z�25��2ΕX3�\h3���2��3H6v3���3��3u�2x�'3��?3�"�2��3o3٪3A��2!1N3}XQ3q>32��2z��3��3��3 $3�a�2Sx(3 �#3u�2'��2��3��3)g3t�2Z��2�3qQ32�2O�R3���2�%�2�(3t�:3���2�@�2��2�e3�u!3�zr3$�3��#3r�2��23F�R3q�2ۖ�2��3��3�?	3���2�!3n�2�3(�K3+��2�03�3��3 �3PKw��V �  � PK                       checkpoint/data/18FB ZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/19FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�U�f����0�#.{��6���"'��^���P�4@���3�1��1��6p�6��S6`_L4��4v�6�Rȶ^��6�,�6W�4��G�6�E(�9%�&y�Dc��ꇶ����6��7_1n6<ˏ5�Ɔ� �n2�
�6`�:�>9�6�P�5N�����䈶8I6&��N�U�7i��N.]6|-C�������q�6�@�6B��ɹN6Ժ��]��6�nŴ�Q��l�6��j�"de�Bʶ��6���5���hA�����[�P��3�Ek����6��9�@��5B�{6S����Y�Fț5布6 ��4t	�*��6\�*� U5Sa%6��s50[�hO�Q78�5�F�6q.�5@��3i�76�t���KE6�Kb�,��4j�Y��55O+I6�Q��v%7Σ�6�?�6@����ec26?j�*��6�,ȵu�5�����k�5R�6�2�����@"z68�e6�ʘ�Їn�4ߵ�16�(���N�~�6fnE7}��:	�@Ic� 煳� 6Q/6h���x8��R�6�#����5��_6�"f�-��Ή5.��5�)�6E�64�����6��i�y�����5I�7�!�5b�R�σ�6�c�6���5J3�4�G�6��6�� �ŵB(�P�)39��6lƵ"�5�����5|ȴ�|�6�4�5�+�69�HzO6jv�6����^ö�,
��;��h �4	6�4�,�5�����OI�2�Z6��Ƕw9�5��^5�87����ft�6\W6������5b�7�[�5X�6+���!�5;��B������+�?6�l�5TZ5�� ���7�A�<ن6�i�5x�75�'/4 �26�6 ��6��V5 3��_7+n��%ƅ�����;6�b86�� 6|��67L̶�m�6$�r��o�Fz;5��?5F������6���6��K6��q6�B7@�y�h�^�W�ܵ8�61�46��s�,��5B�6�|���_(�Λ76�CմH&�����6]�76��	7~����6xJy�  � ���B@*�|�'�6=5��v6Ί86�l �B/����9���d9�6��絒6=���m��7��5�ұ��K�~Q�6O�58/����˶�25���5��P�"y��U�6�����7�R�H�Ķ�� 7��5�|�4���6�<��	���7fM�6�1p6P�z4����Z��5ⴳ�zժ6�@���@���m6I'"5f��6m�+6�3��JT���R� �!�}�I��6#\���/�5ÅѶ�\�5��N����6^54��R/�$��8�P�ǳo����F�"M��:�5�i�С�5F�)7�v�6���6	�7ȏF�0�,����$37�p߽�������h�Ο�� k��w�6�"��.h6ȍ����4w����{�6�S쵖�6��y5J��,&�0��5�q�┧6!� 75�Q6�h/���6:�b��W�4I�� �i�4�7��5nq���J6�9���6|I޶p�,�N��6^�"7*kӵ ؛3�;7(�\4�:6�
�5Є�5i)Q6{^u5\�+��a��I�3��B5\%���(7(�B��ǡ��f���aG6
������TZ�zK϶h5�����6N�&6e甶~�%����8���:�Ƕ��1�z�56然�(�������������6�5�4ʐA61z������E����>��6p�.�0[�5���4���L~������׵T|�6e�m5x:�6��6���В�4hb��@y �B!7�NZ�d|�5H��6��6!.W6J�E6�@`6YEO�y%6���2t�	�6���0U��r�6b&�� @^0��6��F��
E6�2C���!�F�6�f���55
c�5�z5�a��t��5t���;e���µ�V�6t2���"��X�^5fʶk�Y�B��3��!�⶘	���M.�'#�66t�����(b4��6��t6<v%����6�&����y7�܇6��B7j,�~�)�&tP�\��@ݴPKH�EP�  �  PK                     1 checkpoint/data/2FB- ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ۍ3c�+3��93�Ý3�J�3��3E�P3v�*34BN3y73em�3�/3�ӂ3���3<t3[3;I%3/&g3�+�3ʍk3��z3�fa3o·3/�13�3���5�-5�^)5�ڇ54i�5895*%?5�Җ5m�/5x�V5�Hg5��/5ф�5�0q5�5Bz�4��85@�b5!�5UC5�I�5���4~�u5�m$5c��5,+1y<0��0�0/U�0���0=7�0z�0Rٜ0Z��0��0q �/�0��-0���0���0L�0W��0bV�0�~�0I�0���0tYO1,*Z0U��0��2��20e2,MO2 �2�&g2��!2�t�2gZ2��2)�e2�h2�82s��2��r2H}2z�C2d�2���2C�2A�3�#�2;��2v��2>��2��>3(m837�2GC3��3�13�3�؁39�2?d3��x3pb33�83�3:�U3�-3�a(3���2j̟3�Q3K�3]`�2��83Z3ط43���1�[P1��H1>��1���1EW�1�j�13�1��D1֭�1�Q&2�21@C31	�1��1��d1X-2|],1��2�fl1�wb1���1O��1��1`�1Y��1�x�1�=�1v�1���1��Y1�ڇ1��o1';�1	f^1��1'�1d�1 �1�; 2�e�1e�1�G�1/(�1⚲1�?�1�g�1�^2~��1��1�{2[^P2��190�2��p2��2��a2��2��.27�c2f�}2�$W2�2�992��2��*2Ƹk2���1�q/2v22���2�B2�T�2��k2�ڙ2ɟ-2�'�13�1�2@b�16��1�!s1�q2^̶1n:�1�1�1X�1��2�=�1��1�7t1 �1���1:� 2�̿1@2T�2;��1�2�/�1)�1�.n1 1�_1���1	1Xu�0���0�U;1c W1�u�0�51*�1��02�P1`v1��1V�1�p1�Z1��G1��B1s|k1��1�!H1�/�1�>1�1��1���1�1�l�1;��1��1��2�3+2�r�1�EC1���1/��1*h�1�ص1E��1�e1J�1�2u��1�i�1m42+ov1z1�0ڠ�/O�x0�G�0��j0X��/��0r�T0���/��/�΢0��0�D 0{;0�h0��~0~g0���0��F1�i�/�U�0��/ֹ�0?�00Yf�0$��0���0~ag0���0�v+1� �0��1K�0�O�0s|�0qL1+�0���0\��0:J�0�U�0bh�0��0w1�0�=S1���0Ε1=��01�0ܽ�0�1�/B�\/Q�D0e��0���0m��/s�#1��</Õ^0=]�/��@0\�0�y50�,�/UI0���0o@}/K��0MG%/P&�/�C00訃/��0[s�0���0��)1��.0�1���0��+1P�s0��0�v�0œ�0uU�0߉0(`�0|��0ֽ�0�d�0ʃ�0��0�n�0��0���0��0d�y1��1���0�Ã0c�1ë?00��0���0���0~�0��1��1ı0l��0Z�0�	�0 �1�_�0�%�0�"1�y�01�h�0j� 1y� 1���00��0 1�U51�A�10y�0OW1C�01�/�0A�518m1��1UH�0���0��0�8�1�e%1J�0�1��0W[r1#_a1�w01�?�1k�~1v'u1�J1�2Q12V�M2E��1��2Gca2��
2Qy2�2���1۹x2(vV2y�72�42c�1�%�1�82�{�102��s2I�1`g2�xS2lrj2�(C2�g2
�".l9�,�f�-�Z.�Ϊ-�5�.9�D.^1.�{�-��-��.��.�J\."fZ.��%.���-�Z�-|$-�,-���-�j�-�K.K�&./Z�.��-��0�F90�8S0X1�^�/ehi0T��0̌�02��/ǒ�0��30n� 0L�=0!	*01�0C�/���1-1c^�0���0/41Uo0GQ0j�0���0Z8�0��o0�r0i�"1u�w0�C0 �0DzI0Cj0�[�0�2�0g-1��1Lo0�$0� �0���0�1��0��0P�0v߭0j�0TԳ0�U�0�p�1��`1��e1쁮1__�1��W17o`1$n�1��1�N1�P|1�z�1�1��U1�:�1G�g1��B1��1�h1"�1/ c1'�(1�\�1�h�1i�1Ó1.�0K��0^��0n�+1�.81`�1 1a�C1��1%1p�51��F1��1��0���0h�1w]�0�06`0|��0���0_�p1��+1f�61s*0�Z/{3/��.u(/ � .�/m~�-8�8.7O%/�K/��-��/��W/��/��!/��/¤�/�V�.�.���/�3/ZL�/�-I�0��/(�
0���/��I0*�/N`l0J��/!�0Ք�/�OE0ءn0Vo	0��/��0iܩ0�md0�%0" �/��;0=��0u��0�>�/�~�0@�0��0C
�1K�T1& 1Р�1���1�m�1"~�1��1أ�1��1���1�u1[�O1%�q1[)1#x�1G��1A�F1Ҩ�1�d;1
q�1�=�1/j+28T,1_��1�۞2��22�32oVj2Ȉ2�
2'�g2.2�582Yzv2"�2;��2�r2w�w2�D�2-�;2؎U2L<G2�tA2��2��2 �[2?m�2���2%��2�s=1��X1r�0Kp�1ہ*1�X1�w�06�`1��0�B1�Hm1pY�1]951�(1d�)1��1W*(10�L1��`1I�E1��t1��1�761�n�0��1��.��.�K�.��.�}t.��4/��.��.;'.Z��.CR.v�F.v��.���.L�.��/k�/NW/'/r/�/�'O/P��.��k/�8/(nA/��e2�SF2�8�1m��1�m2�Y�1�{2j�:2Ou*25�Y2��m2�7s2D2�ie2�;2�M�152��1��2bv�1�12P�_2[�q2i�o2�f_2�)�1�|[1�3�0�]K1L�1,:41TgM1��|1\1P�1�i1UL1�4�1G0y1 Wp1�1�HJ1�ő1�1U8F1/�1��0�B1�V1���1#L�4�9\4�o4�<B4Ҩ�4Y�p4��H4��E4.a4��*4�rX4�`S4�'�46��3��
4)2*4]�y4k,4G�L4�(4�T4�4�Ζ4&�/4�2/4%63�5�2��2P�29��2" 3��3nF�293��2���2g�2w#3ԇ2W 3a�3/N�2���2;�%3#��2�ŝ2B�2vv3,3��"3���3 tA3.3�n�3�ip3�l3�Z�3�$|3j6z3��O3��-3Fl3���3�S�3y��32K3��b3<\D3��,3iJ�3�3�5�3F�3g�3���3���3�l�3�[
3�2�3{��3�3k�3�y�3� �3�#	4��3Yڶ3#��3���3��t3\�3��3o�3�4�N�3�Gz3���3CO�3/�3��3�5��56b�4�-5W�m4�1�5u�4��4���4B�5&e5<� 5���4Xc�4�֫4�51.�4$��4^r25���4[�44r�4
�B5ֳ�4w��4�T3�-3�9�27�3�e�2	,3��t3�5@3�(3�/X3ܯ3��3��2��2��23�Q13��2^=83��`3��/3~�3(�-3Q�X3�.V3z�3��e3� 3���21B33�Q3XJ>3���2�c3�3A3�;�2�%K3�3�-3E�26� 3��2�tM3<�3��34�3��Z3��3Y�I3{3�`>3 t`4D�3�O4/BQ4�	j4ɬ=4�QR4	z4P�4��R4��4�%;4b�4�Fn4��04�c4��@476%43�4�"4A.p4g�T4-�b4��Q4�&4\�;4hH4]{�3�sm4Jxc4��4��#4,b!4%\*4��4ή?44�r!4n�	4�~54]�4�.]4w�s4J�.4Ke424��3�"x4��4*�[4 ��/���/g��/���/�˜0�p�/�j0;A�/�� 0\y}/�u�00=0}�g0϶�/�	O0z��0�0 #0ƨ�/'a0D�a0+��/��0���/��0>Ġ2<A�2�y22_��2i��2�}�2OQ�2�T�2��2j�2262	�p20N�2�U2�ߋ2�V�2+3�22��2E��2^�2=��2v0�2��2�߷2h�~2���3x�4i`	4�*4t4�4I.4Dz�3:��3eX�3${�3�L�3��3�4빤3�)�3��3��3��04͉�3��4�5�3� 4�'�3��24C}M3#�V3	3(#3��3�FY3�.3ߥ%3(�	3��x3_)R3��[3k�2�R30	3MV�2��3�PZ3&�h3Ȁ3� #3ղ%3�[T3\6b3f3`�(4S-4X��3@ X4 �'4��4w�3��3۞44�O4��3 ɐ4��-4��4Ӥ4�<4��3�	4��4J�u4J`4�'?4~^4��4�E�4�7�4�24���4#��4��p4�y{49�R4��4 �4�|s4\�p49��4#E4:I4v��4a�4#� 4Ifp4��Y4��4j��4k�4S�4�!.4׎3��&3�
�2��m3�W3�3Mw�2�53���2���3U�'3�H�2�s3>XW3$�13��!3��3��d3q)$3*�3�2�3��33m3g��//Ak/�cE/e�/ �m0/d�/�Y�0p��//;�/=��0���/��/s&�/�$0�q}0DR9/�Y0�l�0Ӵ�/��.f�/9R0�Š/��/���/Knp4v$P4�vM4k�4j��4ï34ĪC4��w4���3��T4��j4�Wg4�(43�}4h�94c!h4��C4��'4���4.p74z_�4��s4Qp�4\�w4�4F4C��4	�+4&.4���4~N4���3ْ4FJ4&�3�94yEQ4y\4��4V�04��b4l�	4��f4g44�,@4Sz@4��4U�4Y��4�{4�e4��4o5�4�p5�Ӹ5�YA5T�4�u�4p��4��4�g�4y��48�5�e5���42н4�a�4�Z}5�s�4��i5Y��4_5��R5+�$5�Z�56�4es�3Ѐ 4�Z�3~^�3�\�3��4��3@��3�ޏ3��3'E�3@Ƌ3���3T �3�$�33��3�;3S݈3a��3 \�3�s�3��3;�4þ�3�C�3�1'3�ٚ2�h�2S�2wt�2M�2��3�F�2���2oo2P�2���2�2$�26{�2��v2	(�2n��2o3�D�2��2�8�2���25�2m��2�!�3�M�2���2Zi�3���2�173�3}""3"ɽ2{3q3�T3�>�2�#/3n�#3q�&3J3�O/3�r�2s�53t�-3\�+3S]?3�0f3)��2��J3Nb�.l�.��q/0R0ޥ�/���/�ZQ/�&�.�c�/�V�/6�/�w/%�X0)�v0S>�0qs\/i�G0��/;�0�@�/m��0ز&/ ��/��/]2�/�\k3��e3T��2}��3v�W3�Fs3�Ј3Z�|3*BC3iv�3	�C3|=�3�93`.�3��f3�R�3��3�A$3���3�8�3���3}�3�3��3Uԇ3dM1`�1#&p1l��1��1�c�1�^2�W�1/�1�I14&�1��"16��1�	�166�0�c1cf11y{1��1�B21�n�1��:1�`q1S�_1�?�1PK �JD  D  PK                     < checkpoint/data/20FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�@�3�S:3�\4N�4 ��3�;�3���3���3^�4i�3��3��4�,�3K�3��3��3Ծ:4*�3�ݥ3��3&�4���3[�3t�3��3p��39�A4W.4�~�3�)�3l�3޳�3��3��o3Z�3�Q4�
�3�3�h�3���3E�3�K4! �3��4�o[3��(4���3@	p3�4b�	4���3*��3u}3$C3U��3�K�3��364v[�3��3b3�3���3��3��m3���3�V�3���3(�3��3���3�?�3�K�3�K�3�4�e�3A�3wrZ3P��3���3��3�q4�3�3���3�Љ3?r�3�`�3�T4�=�30�3rd/48�3m#4�4^�f3b�4��q3N'�3�xm3^�3���3�P�3�'4�.�3�$4V�4Fm3/��3}�24s��3�3�O�3�4L�l3�o3��3/ƫ3��30�3MX�3�Ϲ3��3�޴3�8�3Hܛ3�4��D3�fU45��3�w'4a�3�v)4�J4���3@�3���2���3��3`��3��3crS3y9�3�3���3^23���3a74.�3�4���3@�44Ύ�3�A34ߊ�3�;�3�<~3��3��3��3p��3���3��3��'4��34�&�3IR�3��4<��3�d�3F�y3�Ϣ3�h�3Fe�3���3�f�3(��3��T3Ȝ�3|�3d�3�O�3X4��4�4��4F��3�G�3(�3WPF3h�3�� 4��3i�3��3o�3+	4�m4AV�3���3�J3;�4�8�3���3�)�3�S>4bb4{ȴ3f��3���3j^3�q�3�>�3�a�3Y��3W�3v^�3��4���3���3���3u�M3��3F�44�#4�24;8~3*L�3��3��4��3���3�3�3�˪3;Q�34��34�K�3X"�3_�
4)L�3_��3#{�3��39�3� �3窗3ذ�3;4�t4�L83B�	4�g�3�h�3���3���3G�}3@+�3�]�3��3Ϸ�3���3r�v3y-�3��3��3�U�3$�3)�38��3��3L!�3/�3�u4k]�3�3�d4-�=3�T_3
�3���3s�4q�3Tr�3.W4M�3�3��3�׹3=�3G־3���32��3=�I3e`4M�3T��3��23��3+V�3��3��3@�4N}�3��4?�W3�4�T4���2s�3EK=4b� 3tj�3$�3d,�3��#4j�G3�4$Ә3�?4��3��3�E�3��$4i��3�~�3�5�3��b3�^�33g��4 �4��14�\�3]54=�3��3��3�3�Je3��4��3�/�3�3g��3s��3W�3I�{3;F�3]�#4�)�3��e3m�#4��34��4���3�m4}{3M-�3�)�3�I�3���3�i�3l�4T��3�3`�44f��3��+4���3���3o��3�q�3�M4���3�J�3�~�3�W�3���3��h4���3��3z�3���3Ɨ
4�%4���3	��3��3^�4�Ơ3r��3��3p�3a'�3<h�34�3�h$4��3�Nj3SY�3�[�3�_�3e�3o�3���3���3<��2�3�F�3^��3�4)��3�L�3�G�3y~~3���3w��3�#�3+4���3eX4Fu�3N��3�4J�F3�W�3���3h��3��3���3��3���3�*�3�3��3�G�3,��3(��3��4��S3�c�3?�3���3��3d�4�v�36�3��3�v3���3�t�3��3b;3�@4B�3Pj3�J�2���3��n3�4R��3&m!3���3'��3���3�l03���3�{�3hP�3-�4C4�3�3Q��3���2B��3݈^3���3hӔ3�4mѫ3b��3�*+4�3��3���3,��3�?�3/�G4"�3KdE3�3T~j3ul4��4F4�,�3�94�u83ӓ�3Oh3PK��Q|�  �  PK                     0 checkpoint/data/21FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/22FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�+�N$5��$�
������$���ٵ0a]�D����H�f�iB4��J���p�\h� �D�������>q����ڵZ���X���z�4h�� 쨲�������5 mg07��� E�4��4 #�}ۿ��U74ޑ5���_��6����^�N>F�����x�³�?.3 ���"4񹳵?��4s$ִ5Mt$�J�촞c$5�
̵���e��z��ޏ8�0�H4�W����[��N@��`7�d���ݴPv�����	����8���.ݻ3��괏竴�=�3�ӳ�@Vz�~ȴ�m=� �Ҳ�!������T9���0�Ywc��̳����Q���������Zv4��N��s�N��$����N
�P�׵�#d��K6�"�SZa������x3�1�Wb-��gL���ɴ��÷!56���~��_s��>�\0�l�,��P�x?��+T	�������ԇ�"D�� L4��5�x�3�v��
-�5z[�eд�a�4�쿵�ݷ��i�4�D���9�@jv���K���4Hvڴpݟ3����w44���3�[���pʹr̎�a}.��;��gT��k3"�N`*5���"ސ3v�3�4"9'�g��:q����c��M��3�P��\O1��Q���ڵw|д�H����xq����BON5��R!	��B��J�� S����O�m�5�q'�8I�R[�a��3��O5��� �2�)մ8������ ǳ��4�W/���h4v螵	�B�޼��p�;3���<��4�C���O4-2��ԡ�t�3�o�4Q紘�3��F�G!���d@����r�=�vÀ5�
B�z�r���}� Lʲ�m �j�#4��ޥu�7װ��Ĵ�k��CG��V�Sd��������(�������@�{4�E�����kQ���.��H�����eP5$<�4�	���-C5fC���w��G��\�0�m>���?9�8n���$��=z3�Δ4W���	��@��&[d�,+��Z�4� ���ݴG�\��KJ�J|}��i~�кϵ��b�F�$5L��Y�ݳV�|���
��俵|eǴ&I���α�������R�UV��˴8�2��t�_��´�4$���-f�+֗��g`�z���H�1�^;4��4�xX�4�(F��Ųi ˴W�-���&5t��92�l�Z4�h�Iڴ�[״F��P���?��*.���o��{�7����3F�"���`I�1�k�������`�����"��>n��F�����+�&��,�������"5�*���д�X´�.K���v7]5 ]5��5�?D4'I�4�+��8nT�67	�-T��\�4��4+Տ�̾I��?�4�X������I��C��<��4�P�4^f�3�5BpG*���7��*0��.�:}�ݱ�����v3�8'��W���دM3X4�4��2�#��j�34��8�����G4x�᳥�ܵ�&5#	�30�3�J6�����Դ�0�x�^��BxW�h�̴Ȗ�3�C�4*��\k�p	k��˛2*~����k4LV��U���{��>���@�j�
�u���F�(5b�����y�^�5��/��?���~M�����4����-���w�4#7������Ȟ���������h�%��45"�&2����4c2�#���ܶ��Q4��Q��ח�<�<Q����2��g��5G�6�7��ܭ5!�/�P�&�����ೄ��V��:����39��;��)�-���}�E5���,Q�4ٮ�ޑ����3��l4]�I���M�z[��>�/�&"=�{/��)%��4���|۴t���Z ��p��A8��Q�s�x.��E���̴����Z3�����m��lC�������a�Q�4/���@
��䋱�
Ե4�����E�8��4��;4�K����4r
��I��Lk4ށ4�tǳ"o�~�촱��PKN���  �  PK                     0 checkpoint/data/23FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�ai/��*/*�/[I</6�U/BvB/�k�/R�5/�rM/
�P/]�&/��/K��.�$/�Y�/Fם.
d9/��C/X
/��.��S/�=/�Q/��^/.�F/C�.$�0E�/�B$/<`/%�:/:�4/ʓ�/pK /Ƙ?/��r/d�}/��/��.2Q=/��u/n�1/��/e/n�/��]//��.z��/��/���/%�u/�&/aA�/-.�.���.�l|/��/���/GK�/�^	/�~�.`�/'/3/3�K/yb/}Te/=�.�t/2E7/YL�.;�/{x�."?�/3�/b�=/��/�΍.��J/���/�/��$/�w�/�K/r�7/	C�/N=�/���.+Q/�'/��.[�/�~�/7�7/��.f��/2X/[�'/\�L/�:�.@O*/��/\�/T�/��=/TK6/��4/��/ol�/���/k:�.�<�.u�(/ԩ/��.j�/r��.��.ͪ/��/3U(/ hz/��	/}/f/�?K/7�/�G/�h0/S�A/�3�/�5f/�F�.��r/���/d�/v�/��/��!/J�/���/r/JKI/��/��J/ߪ*/�c/��B/x|�/Έ./o'	/��/�Vu/�͒/��@/��
/���.��V/��L//��/�F4/�3v/ᅃ/.l
/p�C/�o�.c� /M?�.R�.��`/�j/���.�/;/�/;�&/*=
/��.D;/iʱ/\"/(g�.�#B/�/��*/�R/�/=��/;��.���.Bg�.��/f�/%�P/麡/®)/���.�VM/r�/�<�/iw�.�:Z/P�$/Ɔ�/�$�/J�"/���/�`/��O/�f/��./�ޅ/#�9/z/��%/�4#/`/J/N/��S/��Z/�i�/�8�/� �.��/�F�/��/�k/��/��/3��.�<0/���.��/q�x/��M/�2/�o/��/< /
��.W[�.���.,�.��/ܽ/{*�.C�/�a-/#��.C��/S#2/��/���.���/�7?/�m�/rg�/�!/���.��x/�-k/��P/g�@/\��.�'/C�/��=/ ��/�ی/[�1/k̭.w6#/�Xy/k��/�ީ/��/�}J/#Դ/���/��/HJ/��,/AF�/�		/��{/c/j� 0rH�.	K/=qM/��/8/.VA/ӟ/wM�/���.rV/�&�/�l�/��V/�Z3/y��/YF}/E#�.L�/�|�.�9m/�̕/ꊆ/v�/�H/N'�/�g$/��/��.\�~/�Q1/�O/��/y�/E��/w(c/z~�.�:/9Ή/�Ed/ua#/�_/�?�/D� /U�/���.��/���/�//�5J/��}/�1�/y1/q�/<�.0O�/�k/���/Ix�.��)/�/��.h�/3�/K�n/�W /��	/��j/g*@/�A�/Q?/Z�C/���.(�d/�/?�a/���.U�;/�W�.��`/��.�R?/#e�/��/�O/m�/o��.Ɗ/=�/�s/8/�/��/�%�/Q�/L�/ذ�/�(0�ֽ.,��/܊�/G�o/��/���/1�)/_��/zXq/�[�.�f3/��/�/�&�/�2}/nY�.���.aCF/��4/��.g�/�K�/�>�/�u�.C��/�/��1/Xj�.���/��//�5�/�0/T�$/�/�
B/���/��/�c-/gj3/��/�!�.��j/��/]k/�E/�|/��/a�I/�X/΋d/�K�.�i7/Iv�/2�?/�/R�*/��/���/>AD/��a/���/Ɖ�.�	[/&oV/��/Z�(/k��.�/�.*�/�-/�D/h�*/�T�/�Ŝ/O,/�O/ڿ�/�>"//O/_��/�>U/�
	/A�\/:5�/�G/hs/F/@7?/���/�/���.�v!/���.�c�/73�.���/��(/�k/��/`;/�/�^/��T/���/�/��.��0Q#�/�"0/��K/
�0/��T/�/�w�/'�?/�J/"��.���.�Z�.PKNR���  �  PK                     0 checkpoint/data/24FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/25FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZT�8�q��cL��=��$�Ŵ� (��W6��C��DC�30߳�N���д~��4��5��e5���h"8���d5��赹X�5N�5B�E����5��V�<g��� ���߳R���;����5\�6��k5�}3�$���R���5��]��5�b�4�����.���𠵸�/5�z�3��oܴ�rS5�۴�����-�*�5�Չ5
n��H5����F�5 �4�3���5����p΃�����5$@D4=��?	S�I+���ו�����u�n� 6&MO��6Ĵc����F5B-��
}� ��4�5Ȏt�|�J���6 ~H�Bk�4�9e5��m3 �e���%���6��T���5��.4�R�3�$5�����W�4�K�Ve�4��E�d�(4C+25N,Q�9*6��^5j�5')��۝�Xn@��Q�5D��D�$4���6�4���5J�(�>��\O55�~5���/�y�/�B�5�ɬ���o���5�<6d�7���2����2 �Z�b#�4.&#5��&� K2k�5a�/�3�4dUW5.����.V���|2m_3+��5��5.Z��v��58`�����n��4�36 Q�2�$���52 \5`p�4�3�g�5���5�*��Y���h�y=s���5��9����4*��a�4�����5@�C4�٤5oB��:53��5	?�\>��0�2�Rڵd�4&�5����j(4.R��.�O��PV5��ӵ���4�۶2A6������r5�n�4(ﷵ'L5r�6:4��5�����4m4���nl��򿵦��4��B4�N=1��S�b� 6�)+�ӛ5P�4 �#3U0>4��T2�5�
�5�14�)´Cg6�Hµ����y���n�4?5Dku4��5����Hu5ȳG�M���IⳄA�3������545� T5�')5+�5̔��b�d��IoZ5��5j���|�4��5�"ɵ~�?��q	5�Q� �����5�9�4|6޵���4������&����'�����:	��v5��/5��=���j�����c�5?���xL��᳉16���4�sɵDPV��ʏ5-o^4�X���µ�����Ӝ3HT����.�X�6�w�E96+�����t|#6�U�4@�2���5��U��>εpO6ߩ�5#�5H���`�����2������5_� ���ǵX%<5���Ur�5\r�5�9��'I��=�� ����ʑ�B��4fز��'�4��ﵰz�4�}�Z��5�"M�]�Y��� �i��Z��jm4��&Y�BMP����4����fP3��26)
�5�4�5z�6d 9��u@�Z_U��T���;�����z���Di�j��5$�����.5�Z8��U3�ӵuO�5D\���5���2OV�ME�L��4����!�5f��5��&5�,��$�5f����?84.0����w��Ҵ��3�`�L5@��Zj5c���H3g�����P5�/+6��`�ʲ�s/6I>��ʕ4&�4Н4�.G5dJ�3¢��yR���i/����3��(��-6��n��_ֵ���45&�X(�\����6�^���l�5��
5,m���I���մ���;�3=�Q!5�ɵ����p!�U�鴖��5��3 4�3|���{��[��
�+��54,����a40�30R���)�)�V�\�5 �<4�Ʋ5�2�5,_!��$#�)*��J���\
6d_��	
5ZVU5B
�4�'�4�5��b5�Jl���5Vr��D �v�55��ܼ��M��5�D���'�t'�5�sa�3`5��J�9�|��4t7'��zs�����4`jb��̠4�&�%���鸵�x"54 (�����gz40�����۵��8�l��(��[A��5~��j���i�4X��5�VP5r?�� �5@I�T�.)6	}�58-H6~O�pj�
���/�Au��PKD���  �  PK                     0 checkpoint/data/26FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���1�K01��2�q	2�M�1$�1�� 2L�1�	2ur�11�2أ2ʪ�1�Џ1a��1D�1F. 2@�1���1�7�1�C2��1�Л1��1�:�1�Z�1�G72���1�`�1�v�1+��1�x�1�.�1Hi1ѯ�1K�2��1��1���1���1�`�1/�2�j�1!2�?c1�� 2K��1��1y�2y� 2H��1]�1P��1�?1�}�13�1Ң�1w�2s��1� �1�&�1�B�1;�1V��1���1�q�1���1_l�1R��1ǃ�1��1=[�1�1d� 2Ե�1H�1��G1gL�1��1r�1�1�1���1
a�1�̆1� 2���1�2���1O�1O�02C��1oE	2D2�R1V2��b1��1�h�1:�1�1���1�p2��	2c�2�2�s10�1�52�]�1���1c�1�Z�1u$`1O�Y1���10��1t��1Ze.1x�1���1��1��1}
�1#��102�N1�:2,��1�\2t��1�2k�2%��1���1� �0���1���1<�1K2�
o1,��1�$�1o$�1�11ӫ�1*�2�0�1-	2�B�1-�52 h�1�Z42��1���1De�1�8�1Ų�1%��1���1⍿1�i�1d�.2[�*2��1�r�1��1�ڔ1���1c�1���1��1T��1�q�17V�1��1 j1R��1(A�1�#1�A�1��2�;
2�2|d2���1A��1�'�1j�d1���1��19�1=�1c��1��1��2�� 2���1u֯1��T1�!�1���1}�1W�1�U)26�F2Oڠ1���1�̞1(t1f8�1?}�1���1��11��1@��1�2,S�1	��18��1��71t"�1�r2Ϫ
2*"2�k2>7~1oe�1p��1���12F'1U��1Δ1I[�1]e�1��1��2֖1hms11��1S[�1�>�1¿Y1gg�1ր�1(��1P��1\�1�2�
2��C1�� 2�1���1B�1:��1�c�1ᠴ1�V�1���1���1�m�1�Yy1W��1���1] 2E��1� �1��1�F�1�	�1���1 '�1$@
2Dn�1��1%�2��I1��t1"��1�]�1Fj�1�;�14�1�M"2���1��14��1�_�1��1(��1ٕ�1р�1�tD1�nO2���1�E�1��`1���1J��1���1)�1��1�ݨ1�u2�օ12��:2�1��1%(2��:1��1 ��1�-�1�S#2�o1��2ߐ1��02x��1D"�1:��1_e2��1���1���1�$H1N��1��1 �z2M�2��20~�14��1��2!��1Kݝ1��1sFo1R�%2�ŗ1⍖1�z�1L4�1%��1���1]g\1pM�1'�2t��1�!p1��2�;2�2s��1E2m��1��1p8�1;��1K��1�x�1��2:�1D��1��#2*��1�6$2 ��1��1��1R�1t�2��18�1���1�&�1W��1B�R2���1��	20��1��1��2�q&2:O�1���1��10�2�,�1�*s17��1�ǧ1�w�1���1���1�2z�1���1E'�1�2�1��1Μ�1��2���1���1�{1N�1r��1���1�2�Ե1f��1i��1�o}1�q�1fȤ1zG�12>]�1�S�1I��1��1��2��p1�'�1)�1R��1"��1�U�1�	2���1���1���1s�1+��1*��1=��1"ۏ2"�61o�1��2\��1��1Q�2.��1���1
w�1�E_1���1P�1}��19�41q�2�S�1���12�1���1�}_1�e2+�2kM1o>z1���1U820�D1X��1���1�]�1�R(2O��1٤�1���1�"1wu2��d1��2��1'_2��1��u1�&-2���1[��1��1�M�1��10w>2���1�K1ad�1Έ1��2�Z
2��2�l�1�&2W91��1�'w1PKe"ڼ�  �  PK                     0 checkpoint/data/27FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/28FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�T�{7�'8�N�8�緶6��7<	�t�7���6@X�6���6�+8�@5��9�5J�6��D`8��(>8�C>�_�5���6�36����6F48����\�?��!�dEc7:��7�|*8n�(��)�6�4;��{��>B8��;���8fܞ8 �_6h@�6։�7x3g����6��T6��A�l�d��"
���跤).7�N)8�&����6���t��7���6��77�+�4�f7�}ӷj3�sѷ�77X�6���7ŗ9�r�����8X:�[̷���8OH78I������V7V�÷����7���6D��"`7�s58�
C8���6���?(8C���ܶJe'��f7�.�6e{#8fo�8�ٟ�N9�u7�L�[����3q���Π8�R׷|D?��n�8���'�7R���08�W#8X>28.�78ID7�}7�hο�|~���=�(�޶Sh)8ā�7fg8H�7�x�Bz�Sh7�$8�����Ҷ�[�i7&8�n:��x����6N@C7�8r�3�Љ���g˷��6��58�;��-�|7��8#�68��#8�>��k#�7�-I�𶧶��7[�<� ��ط�6���v��lI����8),��$�RV��5����6��.W�7< 8�Ip7|�	�0�@��)8�(�\�D�t�%8��<�6/�7O�B8��f7,��f 68tw:�x�7�V�6�'�5�]7P[R7�28�%�8�S7|�;��FZ�(%�8\Ϸ7��v����ض�97�a(�h�ȕ��@�7�<D7b�Ϸ`M��x>=��|B7�@��6�F̷v>!8�Q����$�7�"8���N�C�a*�{_8�^)8��������x����7� ��8��7UA8P��6��>���@����6���7�=�ك&8X����ѷ�<8'<8ϑ/�'�B8�mm��c��8W�98p�7��7�H<������ȶs�986ݞ�Įs�*e�7�6�������6X���2
���7 4��ÿ480�)�h}�6�޶�48�K68�<�6��6��T�$@+�C?��8���6$#*8v�B8�A�ҷM�8C.��xն�<8|�B�8��6Hd�6��6��98��� ��6`�ɶL�����p��7��48��6�9`8��`�P<��N�`7J>8�
6�����7�b884�W7��8P6��d�>���7B78��c�\�7�&8��7�oӶ�%���60g%8�&�8 �����5M�!��?�H@�6�^k8^@8��=�2�7��ͷ�B8� �O*48��C���%���Z��7�R8��'���	�zB8h�7�֫7p���<8PR7�!7�\�����0s:8�8eL7����ٶ�ܠ�U���p��K��8��r�78��6��6Х�0�8,�����6 ն`f�η�7H��6T8pz�6f(������Ϸ',�8��<8�� �X=�7 1*���'���28+�)���6�H�f����6	 +�$X��778A��8=8�з|܊7t2�D�=� 3��緻�!�Fd88lB8����Ja�7�|>��88��#�4
[7q'8�����wV���,��dC�������6�e78��8�S5������GŶ�B7Ш�6�e�6�L7�׷j�2���74�B7@��8X��68��6�\� F	7��6`��50���	�>���7�388���� 8,8��V���6���7�Y18<���˙��_*���6^�7�C7��7�ԶW=��SƷ 4�5?���]7�k��CѶ�<8h[�6ik@8 $��՟8��8�X���^8�E;����.�'��$���<8��68̯^7����k6�O���.@������ڴ�����p7jiϷ��ڷ��>�����L�7��<����6��D���A8x�6P9��b8R}�7�h58�~!8��$�b��Hg7J�8�bB8��i��8(�R�2� �6F�89�8�a�*�9﬛8��/��<u�0���˷8ɂ8A!7S�9��9��Ö8$|Ҹ2��8���8K-���΄��}�7�a870�ָ� �c��E�9�~8��7���%�O旸��͸��ڸ �%���7�?Ƹ�9#M�>�9��۸�@� ��7Cw7@�6�k�8L�8�g�8!Ay�����0'�����8�$!9��8�������$�8�hz8A����7,/58@��6-+8Vs.��88\�ٷ��и�'�7 �7s[��lH���TQ8�&8ԕ�8��89�(Ÿ��շr[&�,Z8
X���H�8�Hȷ!5���+L5��Q�@�Ǹ�#�6}��8`,6��V8�r���g$8س���W/9�����w۸!'U��,+9��8H|�8<>
8@�޷;x4���D�6e49����K����1�%S8�*�p'�F:׷p��*=�8���7�J�7����4�_�挟����7ճ߸0G��Iad��P�5.��PRL8�5ϸu��T�9�ߔ�fm$9(��Tb���Pd8�и�n8�O"8w4*9@��5�,޶�ݡ�R�8����Va8�4=���7��]��_��F9���7�)���t�7V�8�QX6���@�����@8�{X�5�7V����\d��Z�70�ζ�(8����m8����t��7�]Y����7_��86\�ͺ�8���8���7d6��÷m�������8�*.�r��8�u�̋6)�I8�:q��	9p����.%93�`8D�K9�=�7�.�T��8!?�8P�7@��4���(�D�@�5&�8��ĸ��X8LK9M�S�*>���l���81�w�JL�2��7\*ظ�
�u������7U��8=@�0޶�a98�l�b�'�T	��#O80ŗ8�~�8�Ŧ�<zӸ��'����8�N7S���1�8JT�8�ַ�8r�9�ȸ��෬Q���{G8$���#θ���$E̸��<8�^����c5M�B�Ht7�@Ÿ}0�726
9����8
�`���3�Ӹ��Ō7X�7�6P7�?�����7���8�~<������=��$�и��7�L�a� �:5�����a�8,�X�6��8��'8@͝5�7��7���7@8��?ME��3�7P�7�̰7������8���na7c��d�9��8F�d��v���J6��+8��2�Კ8Z�[��X�8�sL�&��8uv88�ݸ��y�>��8��߸��8�m�8�W9/"�8��!-�
�w�@�6FO8Td�7�n8���6�
m6~H�8b\}�V�N8�S~8beE7̹"�H���s�8*Щ8��8F�'8��+85T��Vh8�/�8���7���f�8��̊:8,|�6���8���OZ�`��8�N�7L�x8I'"9N�8��ȸ�E�8Ԡ������ �s�ø��o8mz8��8<���U9ܪ8+'����7�%����8^���[Y7(pQ��ڸ)�9�6�8K##���޷L�
8���7�1;����V�J�aG�8\�������C������8�*@7j��8����8��Z7 �
6Q��8��ʸG$�8#2�8��7��8��������B�8x)7���h��?�tE��X��8H3ظ���7���8�9�$8H�8�9 o�n��59�08��9t�ͷ@����6ʸ�T���.�N�2���+�����8X4ٸ���7EH9�䂷!�8N~�8�dݷ�8 �4�t�	G8 T}8Xq�7��8z(-�@h�7F�o8��W�\�H�r ظ�c�6�1%�@�)7�2R8�͸�w�]�*�z 󸐮\8p?B7K�W�"U�%U޸�\���θ.�i8@��8��!9Ȧn7�[���,��G~�7�V9�
Ҹ�_�7��p8h-�7:�9� ��]d�$
����R�8X����@7
�8B�V��$:�0D	�Nr��Lm1���!��h7�	�5�9�����6lL�8���8�̙�mښ8����JT�7��7E1�����7�7�vY�|Bd�*l^��X7�8����z���o7�Z�e7�K��ǌf��b�i!����I��?�8��h�ppa7s o��I�8�蛸�1^��d7yB���g7S�8]����"�8�F�7/�8y\ⷬ���#��8�JQ�fk��~�7ӌe79�98)�`�<.�RX���8*5�7{��7Pd7}A�8�j7�O���ę�[S`7=:e7�P�J����J`��_��x�������g�N�8}�B7��d��h{��#a7ݕ�8"�����b7�A��(p��o�7P��8(0�8 �G�V�7���S�8��]�L�6���j�[7��N7g雸c7�9s�

d78�W�����φ8�$`��������8�E�8��8(���ƕ����W�7���u�A�J�/���b7a)s�W��7�x7>�]7O�_7�J7 ����O�89�q��?[��8k7d`T�a�y7#M��!��Sub7�N���@��ܳc7kY���f����8(rd�>�d�Z�d7\���`����L79Pf7L�6�
�8��8�Md7����J���Q7To?�c�8ۢ���o`��,����F8P%M��E���Ov���Z7��]7i�%�85#q���G��/j��7!�l����7Uoj�Q�g74�8�_����8D�08kE_75�7�n�@�C7)1e7��8��_7�ә8l�b7�_��7i�����	�d�bd7��7�Z8Z
 8Ȇc7!|�7;T]�ξb���8��]�'�[�\�]��ߚ8y\7IW]7V��ߨc�R����'\�`d7�G�8w�N7���8�ɘ8��X7/�_�d�_7����_��/c�W�`7�U7�$e7uT��*D[7��^7Fx�8��I���c71�\�`�_7������c�Fd7�[���`{�}/����8�K�8.�����S�#�8�b7��c�]L�+�]7�ؗ8���T\7ꉚ8��^�h�^7㕁8B7��i�f7 ��8�a�b�8O
���a7e4�8�H��,7����8�h7�����`7)[7�|=7R��������W�_7�a^7u�����87�U��Q\7���8�W��Ƹ[7��87��89�~�n�S��7�阸����K��8XH�8���8�W����8�"X7��\7��8Wd7��a7�Q7$��6��8���8�,b�^�-��.�8�ߑ8�vb�ļ(�(ʒ8�q`����8h웸�J`7Sl��[�g�o7�VS7�n7d���ͭO��U7.�8�� ��P7([7�_i7XK��nJ�8����/.��Y�m7��k��"��S�8���8R�`7 9U7�[7�|b�Y���F�`�l���}����c7�;X�x!�8����[�A7J�8�d��?d7��b�Ta�8���8#U�8WI]7ְ�8���.�e��e����T���e�Y7L d7E#^���]�X{�7�yZ�=ᙸ��_7Ɣ�8��}�7�ƛ�q`7<h���
a��P_�"�g7БW7O�Z7#�c7��7�ֆ7�'h7N��X-��H:6�#ՙ���e��`�qњ8��i�+�o���8�`�DH��rk�|�M81l��L�Y7�\�m�'��8�f7�U���	8sPe8qre7��T7 Q�8 *f����8��d�mi�ܴ��h_�\�J�8c^7�Xf�cy\�iΙ8Q`M��a�P�d��3f7ɚ���7�jf�SW��T�{\7Q4�7Toc�8�����c�=\_�$hX��ޘ8 �_�Y�d��[8EG�Қ��١Z�o1R�k7�8�����l��Jr��"`7×F�h=t7ރ����X7������`7���8�:`�􍄸�rp8{"���3f7��8��]7 {�'#�8�r71�`78��e��7c�J�d7�*�8(��8��`��>g7��'(w7-�Z7�<!��V�)Q_7	�TB�i�k7�O��Tz��z@��N�;���8��1��BZ7����]�'�*8�Fe7���Zi�86r�7�W7�DԶg�T7�Ym�H�k��U��`�^�X�L���28����3��a������І7�-y����Khķ b�Pp�8v?��v����� 7��7���7�:�8$�7h��8�Qy�^j�7�e�R18o��- �+��7R9�7�J~�(�2��U8��D�.8���8H7��8��4D�7����~縎�����8\�����8 O�86�9|�7b	�8c��Z��7NW��D�W8�	�5bO��E��7�4�7A�]8xS���z�8�������8#�]�*O�8��z88������T��k~����7�;��v8z�������D���8�P�8�������Uv�8Ѓ
�<��8�Y�8�9^8����������V]�8n=����8(;�7*̢7��7Ԓ��s���
���7�r�8��8��\�[=�7�v���ڸn���r�7��3�L��8~}�%���8a8�@긦q����Y�9�Ȉ��m�8�9̠ 7$��7�2�{W68;��@��8t��7��8�r��g*`8��8 3s4Ֆ��!�8�B�8N��7D��՘�ŉ�8�t8Xie7<۸
)���ȹ�lU7yޞ8B�o8H_�8�U긐�	�Z��ػ�9��81�9�������8���7�O�?��7��H7��8n��B��7�N}��B�7� �7�k䶯O��i]Z�B���B�8�'�7V�۸��ٸ�,�7T�8*� �rw�7���7�y�8a۸�KZ��M�����88È8\�8��O�\�����8�1�o˸�����9���7��÷C��458HN7����������7.[�8�_�7��9��8�8��(27�ݻ��t������)ַpԵ�P�9�_�(�]8��5��7V�9R� 8F���kڸVa�7��9��8��38L���M9�����a{8�67�G�7	�׸v�8�&�7��뷩4]�"�e8�̃�Iu۸��7S��8&M18�<�7�(�TV�!|�7[Ʒ����3[7���7��O��ce��/[��u�7tI��:28L=z8��7
�7�L��$֓��hܸ�T)6�����۶7h&���8t���U�8�暸4T�8��48̇��!�16�y��A��7Q���6���:��8:�9>M��v�7�����W"�X��2@ո~���7�H�8��6"}�����Q���3j�`�8�G�8�� 7ж�=�y8�8��|�O�S����x��L̸�27@ȵ8�}3��䵷�ඤT���L����ܱ7��~��M�v�{8���828,�^8�+18������� ��B��~&�7��薕8�2�(8���4��8N�8Շ�8?+��`�9������7�m��Q��7H�8^J�8����Y�24�S��7 !7������ �@�7���8X4�78-�7@��8����^�7�ʐ8a/�Nu縼�7.���冸{��ڷ�7`��8�1�8�:�8�8�H�h~ܶ�d9y�~8���h&׸�����^7��9�u�7z%�8���8�3��8~X�8����̷���8z�8p
7��W��8 ��8 �7�D�7�/8oiq�ƛ�8�����[8���Y��8��7��\,8X���6��zy�8Mr9"1�8��7�8`%�rٸM��58��7�x��<۸D-ٸz��Z�n���9
��5�^8İ�8�8���߷`��8���z>�C��8���8��7�Z8Hx&��X�8D��7Q�8|@��vp18�>�R�7�︪��RP8b3�7�M����8b��8��^8~A�7i-8_-8��7o�8�\����8ȴ8�������f9��8�J�{��7Ֆ8��7M9�X7�<��p`����T��D�7�@ܸ'� 9^w�8������
7<0�7Dk�dF� ��L��8����V�86��8�r��n��8���g�3^9��ڸ�M������&��8����7���R��z~��*������_8���8\cn�0v!��G�7.�|��q�4Q�7�쾸�Q8�V�5��H��8�����X��|���b7�	�����%Ir�IX�7v��8$���"�7T�87�U굟_���縌�5�UH8��N6�,�6�8��880�ʸ���7��7 �}�
��7~ŶXx�8_v8�8͸Ar�68���0V 6#��7���8!�3� v�8Np63�����]�(��6��T�7��m7Y�y8��ԷZ�6�^��*}���N8��2���8XF�7K��7���5L��}�6��"��u�F>q8*]���e�8�b��&�8d�]8�,8j��5kJ�8BM�7��C82j8>_��
�7��\��n�6��踌7���^�ZN%6�՚��K�8L�8"��p�����7˱����9���z�'��胷V���-�7�8�F� �·Z���M85�7�t3�����_�7��6�3�8@m8%T���ˌ���8�l�7�f7��7EP�8��(8)5�7��|8DY���7����J6d�7-��;�t8[�7oV���ϸf^����7�?5ܓ�����7 �P�hw��.�E7г�8$Z��'�8O�ֶsG8�]�7�f7oG��s��7V�.�t��7�d��7��8��a��,^8D �1U��Nί��/�8t�q��f8/�7^\*8�E7�Ci�4'b�fO=������:m8D�� 6���y�8�rN8��Z��88�8��7@��8	T'��]�7\�θ
\t���F7& �7$�Z8 ߇8BrضR����>8�ȗ8�[R8
Ԗ8�8���6���6��8��7	 ��8��8{!�8a�7�W����7��8�38�z�����81�8Q�Z�ܭ}���	���7�/8�
���8P�08��ѶZsa7̽8:G78b�K8;� �7���ԏO7b7���7��Aڿ��<c���H�Ȣz7�m��C8^v�8 oh6˨8�9�6�=/8Bj�8�հ�(o�8g����ͦ8�<����58C_�X޾����6`��8�?�7���8��8��b8W������&�8�л���6�*��8�J����u���*8ܞ`5�n�8�Ow7-�8d�>������B����շ�A8B7>c'87tA���1�7��8@68{ʝ��i�6��3����8�8�	��p����7��2�����b�7n.M7uFθX88h���������8��7�b��P �8�)8��8���&�u��Ey�F�$��F��Q���x�����7a�Ḣj�8�B~�u��7`2'�<�7�_�����7��x�Z�7~I���c����72{^�p\����Ӷނ�|)�f4$8��<���z�w�8zh��[��� ���A��ġ����{����0���X��1��\�����<8�7c0 7�L7aI�7Ζ���𷙞�6Z>i��̳80Q� �ڸ��׸#�	���N8��h8��8����܋��W�6Ơ�"eQ�y� 8��$84�8/�?8��f8�M�7��M�����P���D�8T8A�o8��6
"e8~0
7��7*ռ8ej�Y'�7 "�2<^�7+p��(��8@CF4�)����0�m{�8�y;8��37䂷B��7���7ꂶ7��� �w5��b8I�зQ�����7���� .�\T�8���8��B�y����J6�ڳ��"[8�c8z�����8h���"8��8� ��\���^N�7�f����8�(���6�Y8D�g��-��V��L��8x��{ķl�=�l׸؞�8;� �jٻ7���7n��¿��8�8n��7R1}6R�q������8�A�RS87}�˶��6�/��Cd8��7C�u8#\k7� �7`�����Z���r�\76���G��,$�6�1��_�޶2>:��M�����58��6�8J8XW�7��38�P4��_-6�7 �Z�<�b���G��ܧ8Gqv8��;���̷R�8�K��s�6�\��|���8JΧ��5��V<B����Y �΅L��N7HDH�,�8Ы��w8|M�I�Q�
�P7'	8�@8h�8�(����I7��U�S���8�]�ul�6q�P����8r8֎L��8v&����O�f7�^��0P7�p7/B7����6S7���7q}8�����N����8�1�7��O�ި8Z����7�I�yĔ���8o�H�'�J�@`�MSQ78���U��U�4�K7���~ 8bW��դ��CO�%*8��8���7�D��'U�ϧ8S���i8HQ7�<7�%�m�V7j/�7�0��P�k�E78.��bO7������5ܔ�7��L�(&8?�8ȦF��b(7<��!�L7Bk 8J�8��R�V��.��&�I�������@%86�T7`<M7�`7L�Q��|�7@7�'Y�:.T7�L��C�7�&��F������K7�U868�8g�Q��8`�W7sES7��P��1P7QE����`���Q7CO7�qO���=�6y8���)R��0�N�-��B��7�rN7�>B7�&�7�� �K��-W7�K8b���)L������?�8�S8����b
��R��P��T7q����8�c�}�74BD��R�x��;�p7��M7}﷙�L7��8����Y7eW�v�F7 �8<�8��8nJ7�O7@�8q8�rZ�/�[� F7jwM7q��ʬ�EpT�T�8�8�P��^8@��N�,��z����$�d����R7Ld�7bn���M7�
�pC7����`S7�@"���7��Z7"l8e׷�M��8V_K�?�S�(��fB�<V��T�Չ8�HQ7�=8�F7��hD7���7DzP7P��'�]�U�ַ/N���8��8�U]�A ��FR���8wdP��@R7�S�n�����1 M7�8A O�g�K����T+8,�Q7�N�w�J7%շ��M7�LR��J�7z�D7�&80�P7�d8c��7ejK7��8�*��Kf75C7�<7�5P��\Y�e�67DF�d��5?�ӷ8,�8�8�����M7��U7�B����8~�8��L7,S7��S78��9���88\#��8Q7�jW7?(O���8��X7w������Z7�d@7,��61%�I�F7�Q8؃���X7Ѣ8��O7�.�X�27L7�vQ7B�O7�8�4�H��V�8��8%8Aܗ7��7ʙ�a��58�6T7� 82�T�PAM7�8��6ʲ�1�M��4 8�wR�����J��O	8�R��;82�.��S7i�8��82�7�<P7WN��d86�XF?�N?8�q��[�Os;7�p��c�mm��K;7�>8A�
��_�g/�6�ݘ7ۂ���8 Q�Ѩ8��ijK7!t8��S�B�Fr�F�8��V�� �7�
Y7�S7�$N7�I8l5��;�l_�<9����U���8(��� _7{R7OEU���@�PO7�80Y����lC7��85�������K7:�O7������|��*2��Z@��_�[����D7��|7��P��O�`�s�O��8g��6��S7����<R7�U7'�N�T�Q��JB�s���/N7����
8~�M�p�N�)MQ7BX���8 |�xp�D9��p���8)��$<��|���L�V���L7���#޷�c8*8�@Q7����N7��ȶN��x�ȼ����Q7�X������
D7ʐ8ђV�{ZW7������R�a�j'8@j7�WX��}8^Ms7,AF7&3Y7�WN7g�R7�"O7z�K7�P��o8 8�.����T~8
8�8��6oJ�����`8�[8M�P������I�9�Y�W��H�Fn�t�S7�
U���8����BM7���}ډ7���XI���7��8�u7�Z6�ቊ�<1�0�﷜�o����E��8���H���_�7^r8qA18R�7�s_8��8-����Ƨ���/8*v8:�w� g�6%7b8~|\8Xh�7HAX���_�Q��8(��7&!3�d�a8�N�8��_�HԈ�H�67�6�7����fz�7�ʅ7�|·���8����L18��~�8�7 �7�_�74ʐ89{�8HQ�7�_'緎>�8&�X8���ʁb����Ò�7/�38�%�슐8���7��8�j�
W8�Q�7Cҏ��N��8q�7T����~7hV2�^8�T9n� �6:�/8���8Ԥ��{~7�W�85��A�/8ӷL/8�Fs7CΆ7(��j�6:��	��7X�v7<�\8@����:74��xy7J�08V��>q�8����_*�7p�׵j2a��H-�]�C�@�l��V6�68�%E��>Y8p�"�`����f��<��l;y8�`�XI�7�ߏ�>搸���`O8j+�8�Uh7��71=/��ꀷ�,����Z����7G�����`.8`?�ԣ_8@օ��з �_����N�8P��6�ݎ�o%+8�<?8lKv7`R����L���;�����sOY� ���+17��07��]8�N������l8^�6�]8w�8��-8��\�䜬7~H�7�����8�6`�8PCf7�z7���8�~z���18ಪ6�X����6qI���j��~�y���7��7���#_8+
��&�7z8`����7�����<~���v7��`8JE��$���_䷗I�8 ��6ĝ^�D$	���-��q"��\U8��Z��8N[7&^M�^A7#`8 [���w�J�ܷ@}����47d���#�8[%/���^��P:7�G8��ٷ�8�?����O߷��7+�7ס�8������d�������
�8Ď8L�1�,�X8���6�^���K�8���6�%��Jg2���18h�*���ܷ��{��;b8�÷7��%�O��O�ٷ(�`�6��7N_������78:���l �7�K���D�&��7M�7����֗8�(38�hv8�� �K�
�$ �7r�e��}7a����Jc8\a�7�}�8P/��G7Y8�gڷ���6�xU��$�'��8�����2�Q�7�&�8𙔷�*[� �C6�Z8��w7���Jr��^e5�p�6�M��E�s8�u��q��xn;8p�6�
�71�a�ܰb��~2�I�8�ܡ����v ��bp67�6�A��7d'G7AWȷ�
Y�m��8(�ط2I 8���6��� �b�����wY8A8̒�lW/7�7���~`�9]�7Z�j7Td8���7��0uV�qU��"�1�0F�7c�\� �`8�-�����A���a�Pe_8��f8�"ӷ�͑�0��6I�8����fÇ7&_8�ys7����GP�x�86���q�8������@��፷8���t�d8Z��2�6�|nG�@j���_�>�`8���80�6;4N8.�@��x2��1�@j~7�v��yx6��/��q-�p�67��L!�0ɐ8#U[8�F	�9(����b8��������7��77��7�v	�z]B����6�*)7|*'�b�;8yP෶�8KX_8��8p-5�ژ�� 72� ��V�7p;_8���#�T8@ˏ6C�8��8�`� ��6Ni��,9�8~��80�^8`
P��햷J�t��Q(��0�<AT7&dT8�ߏ8"�X8��986Q�xe|7@`_�/E�	8�e=7>�8�a+�+��� ö Ǧ��Y��T8�	8�˶�A�6t�_8t&��8�^8p��6�-\8\����5:�������7��R8�!�5�S�6DM�8��2��sa�W,䷰���`@���0l������`��]}7�,`�����AQ8`b�6�.��;|{�಄8z�*7q8.+8��-�<uc8*����O8����Ь�����6�7`8��87��8x�=�ވ08�T28��X�x���<��7����U�\����8��r7�Jy��.۷�=$���#8�f8��#8����K8J�9��B&8�� 8�t&�?4#8��#8�&�)���@"� �#8Ad��$8V�8��#�A#��#8S%8�J%���!8�L!�4�$8bk!�d�#8� 8�f#�e�$�����d%�8�0�ނ!�ȿ!8�����%��O򷜔&8�3&�>N#�$�uZ$��8�/#8X@!8�d#�\"��8��"8��$8��"���!8t�#8Xg%��H#�C8$8�Z!8��!�l�8a&8��"8��#���8I\��"�(��7 s�7^'#84�$��z#8);"��a#8 j"8"�!8`T!�X���$8�"!���#���#��@�7%��N%8 �#��,#8r�)���83�"8��'8(�)O&8yz!���%8��&���'8^}�k%���#8�� ���#8�7#8��#���$8P)�7k"8����� ���'���%�ՙ"8p^$8i�(8�%�"���8�s&8�&�Ԧ8V7��i��7��8�G&8 �,8{�$8��8EW#�%I%�{�#�b%���%�($8Y�!8��&8{�!�Q���$8�"��V#��<�h��8�$�jv&� 0&��f$8��"��9 8`�8�z�7��%���!8��8�]������ ���#8�!�0��7%8ͥ$8H�%���'���!8*���� ��Ĩ7$m!8�}$87��%8� ��#8tA��3&�)�#8��"8Z�"��#8�R&8` 8�� 8�8�O&��%8Z&�A�!�
�%��"8N|#8�!'8th$8���5�)%�߂#8��$8}.$8��!�_'8�#8x�#���#8�i̷t6"8��>�7��%�6�"��$�Ѡ#�)&��@6�Ś�6n�8�u �v&��SķN�$���8^�#�4'$8�#��0"8v=8�v%�*�"8���z#�D�"�F %��_8K�&8uz&��n"�� �/��2�$8�e%��80A#�a%�W<$8+7&�h�%�O$8�� ��C'�<��7�E%8<W#���&8��"�R�"���%8�"8�%8��$8Őc��+�ƌ8$i&��M#��"8�� 8��%��\����,� 8�T$��b$8�$8��#8�#8��$8O"�� #�j�88*o$8�8ü&�Ѿ"�zC&8&8q�%8*&�s��73� 83�8J;#8N�+�z�%8�*#�R�%�I!��%8n4�6n������W8���($8C����7� %8_��p��&�a!�#A$8 �����&8{�&���%��� ��0$�&8fO81�"���$8;z%8Q�8�o��k#�2��7�I'�,"�g�"���#���%�ט$8�h%8�$8d�%�>�"8�"�Q�$8�� �
Y���"��$8̚#8��$8��!8`^#���*��Z"8!��/���&818#��3!��$8.�"�z"'8i�$�:�&83p8�7"��]!8LS8>�'�QC8�d%�ݼ8Qa$�c*'��$��"��� ���!8�����?�#8�
8�� 8�k$��|$8�K%8�%ö^�U$8��$� �"�\=%8�1#8��%8�(&�G}"8Z�!�{��,^!�"s!��2&8��8��"8H�%�tD"�!'�
P�S}"���'��!�I����$��5'8�@!�+�"��$#8����&8E��V�#�̥8D"���!8NT��J%�b28��$�m�$8��!���$��y&��y&8�#8 !8��#8�+�]�#87"8��,��e&8��8�J�b$�7�ߵ�8pn"8y�"8Z��Y�ܷ���B�$8�0��:#���ۢ$�>!8��%�b�*8�x��AX*��#8ys$�w�$8�}�3 8# %8�^�%$��#�DF%8N���O8?.%��#��:"�>�%8��%��"��K%8[�#8�W!��T%8�$�3��k$8�
%�
�"8��t�&8�o��jq%���"��C&8	�#���#�,v#��8&��L&8��$8K#�="�j�$��Q=8[Q�����8p�67T�8P��8��7~��7��7����8 z�>F��.|8Xh]��/b7���Q=8lh��lBh7�p�7�l�����8 x��������7�o�7�Q���8�==���y7��8ؼr7{y6���%�=<=��Fʷɳ���w6FQ�8��F��ݜ�1{7�Dp�>�����@��"�7�u�8H<q7<ߝ�t7.�o��Ã�����LP��\��8�+��P`v7<98��u7��� �i���=�j1�7����A�8���N�П8Z��R+���r?8�����8�R��k?�֏7ր����l�?�F�,��7�g6��&6~���Hn�7R�C����7�ـ7��|��8�p>8��}8���p��7�.�8$��7�a���^�8�������v��u7>ʓ�+YG��Eu7�~07\7<���x�c��0B8��`7'��8�x7���8`;�8�?�7���L�I�Β38��7Ěk7Z�x���8>"�8�՞8������8K���+e��BН�f:�7�#��]�=8�n�8�
W7�88/v7g���#q��6���8v+�8.a=8�3��T�7�k�7Vi�8Pʀ����8l箷 Hx�ʁ7x3��̞8�J8��:�B�����B]�7��z�́7�t�7�맷�1<�r�$8mǝ�j7�1�7��_���;8�η`In��(�6���[���f�8(Vv�e@8A>����48<B�8)	'��>� �q7897˷<��V8�����O8�_���}70p��۞�N����3������焷20���x7冞��t|7���J����"���}}7	Z��s����{7� ��X���:8,d�7Еw�oڜ8�ň��k�8��Q6��<8�3�7��˟��$68�F��h�Q7H�u7�:��z;��4�8��74I>8BN1��|�����8w��vs:��П8pw�l�x�x7��7��������8�*=�̨����7��7�2=8|Fo����r��pÞ�pQK6�f�7�}��ݴ7h܈�(rz����6�u7X)y7��y7�x7��!���8�Xu7�$��\������>�V��7��8��7{}>8@�}76��� -m��r^�xI7)�(8�Ԃ7j�8|ڎ7�(7�~��7��v�77�P�y7�y7�r�7��7J�A8�������J|8���<��b��!`88���@ā�7�I��&C7��3�}b���Jl7���74/�8(u�3R;��ma7�3��|ϊ����8�����on7�6<���/7us78���7�i�8 h��^Qη$=8��q7OV$8H�i�P�����������M7�!8�o�8��=7�
�8�8�7�v�8�3�8��:���y��-��xvR�2������3# �Tś8`n]�H�a��=9�/�f�L?8 p��V�8b�7 F8Hͅ7�D;8�e{7��8�a�����7���8(r}7�br7�C�8���B߃8�՛8��=8^񄷔I�8P5���Q>�|���'�8M�O8 �*��O8*�380�n7	��7���S�:8�Q�7��<����&�����8���4=����@$;�v"W�R8��<8Hs�#���Rg���z7�.V�ۙ����c��%�7,q�8P>�4X<� ���������w�,�8j�ڷ<ٞ���7�dz7��=��F��p�7dV=��"���BA�Ny7<g����	8eT����u�@ew�{�58ԇ�8X;>���8�z7�G=��2�� u��1�7���"�·(�v����� �7�VZ���y�^�A�8��/�t�;7��m7��h7v�8�,85]=8�/^70q��ퟸ<8=O8x8�7�.>8Uշ�_�7�����G�7��8����r��X�n�QP=��8��~�0zs��<�H�8��8�88"��8(s�7�Uȴ�w�8�x�80���7T���6���ϝ8��q7P�}�j=80�v7�<��j�K�mx7�f/��H\�������8`q#�hE7<1�8@�S� �v�H/7@�$��k��U8��g����j�P��7q����I��(�·k��8�L,���{����8\��8Xr�7@]�Ff7��˷���+?8]\K8���V���"�8]�G����8��7� )8��ha�hw8��A7 }K4��a8(����:>�T{!8D��6?Cj8n��7�!�8���%�28�Vz7\2L�{É8܇:���;�cm!���7��}7�8u�,������cf8Up�=���p �7���80���c���8x+��fR����
z�7=B��b�P8O�}8�p��PC�%6R�٢�7����V��8�ũ�-K��q� �(��84sƶ9�㷸�7TP�8�ȓ8M�7VF7�‸G�8�k��D��8H�������p_E����6dJE�a:8�	�����7�h���?87"i8t��͖b8����<�!7�T 8J|������+����8���7@z�7���8n�������$���71�7Z�1��ӷdR�8���=�u8�o���e��ѷ��A6'$���<���)8�3�7!�n8\��8U%83 ����Z������ 8xg��ģ�2�8j�+8��8&�7�ퟷ���8q��8�M!7��61�8 �g�`�v��뇸r�t8���e�&���8�#�7]�N8r��H�жԗ8ťK��e��4G�8���6�1�����R�X8D�6)DW���$��dܷ��p����7*�)� ��8�8tU8�,�l���8�w��q����n�[1����"��8�)��;��7iD8NĜ8�7♶�����܃��(8��8��]�د���j��"8*@��ϝ���7CШ��AK8a���z{�8s$�k$8���|��7��f7��:8�荷8F��`��Kr8��18��|8�`7d�>r8�ф��d�8� ��O��7�?��ھ8�ͱ8�[e6�N�7[��
�����7<�6@M�7��S8tV
�٨K8M0��%8�~�8���ʝ�7޹�8�@&��L�8�P8n�I��ٶ�2�18�y�^ʕ7!��8�!�wv��3�������YZ7HC�7�����Y)8�|j8�Y5�pٷDH)7r�70�8	���S�7x���I������֊�=���1t8�L�6�ER��	���u��a'�me7���6$ηf��0�����7&��aH���4�	��0�m8@@m�?�H8��8���8\}��d(7���7�7��U���0865���G8�q8�^�T� ��8A�74F�6�m97�#S�,�C7D�;�7L7(8"�7�8s��O���߼8@�^�ὃ�<N+�&�8���7`�f��y8�!8�g�8��8S�8����,�Ƕ�2��E8
��r&�7Gjѷ�ʤ7j�78(��7x��T�|�ҷ�4����h8R�>8�,2���8��48_�N�R�@7�8�8�e��h�87 �k4r$�7��'�^���2�{8��c�����z�7����y;8Y��x�7Lґ7�y`8��ȶ$�7�{���L�7t]�8���f6y�\�H���8�G�|���b[�7�g8 s^��(q8�w8�8��.���;��l�7Ҝз7$�8�zq8�&�7K�e8=EX��T����7����6��6�ő8E�7�l�8n^8h��8��82��8-I��ǵ�7K�8=���98�?˷˿�8��38r[�χ]8C�E�v`8�D�8Vxӷ/38��U��X<8C��8R�8��2��q���~�����>ك8lᚸ)*ŷc?�8��c8"aI�ZՊ�$�7N��8 }6!x��(�^��g4���M8�'o7���8�wc���7�~8D��8~��7�°���8}QC�h��6��8gh�`�<6��[���ط������۷�/7}8Xs7D�\�":�77����_���F8���8p�%�跾7�I�7�>W�M���x8�� �
�8�d8��p���8�E��D�7r�c�h6Df8��8FXַ.w�7>��7��V8>7H㋶���4h8j�%8�08�#8����I8���d�`��ٚ#8���l8�� 	8�b��򃊸n��7\�b8��i���82ˋ�r�%8�䇸��7�o$8��8��76܌�hF��v$8*�#8�p(�=,�� ����7Yu�8��7�lg8�%8�f��b�#�����Hkj8��8�7.�$8l&��g]�����7��j��ɋ8&�鷧��qi��#�ا���7�~��i���7X��7���7���TH8�Y����7V+����8V���Xi8\E��ho�8Ԋ�����xh��i8�$��$�S9�ô�8�kk����7��]����>(g8U�����&�3�7��8t3%8�t��xk8g�8�D8Ri���]��"�,Eh8��!8��c8
i����T��7H��7C�"8�j8q$�����7`J���������K��7*Oh�L3�8�:�7,�7��%8�&����f8���7�tf8/�j�T��8�[78�5�7}@f��%8{��'�s\�7�Mh�?�g�� �����8JX�7�w�H�$81H��n%8����U�7��8��g���k�l�����8p_締��7�r$8zy�7��7�$�f!� %8�ډ8��i��&�5��76�'8m#&������%�珉8�!����8Q6&8"6��J�7l�8� 1�7��8�?%�~%���7�w�|k8��86:�8�d�7g��=��7�Ch8�h8��h���k8Caf�tc&�������j88�i8����{h����7*ag8j���m�7x�28�|8oi����P�m���j���l8��"��ߊ8��%��l8j#��k8��m8q�l8�X�:G��1f�b�8����<�$��h��l�7�&8]�$�Vz 8����p��7gi���u���H��G��"���d��<�7�&8��g���#��K�L1��!���Ő ����7v��JY&84+&881������V��7�r�7ŋ�>ku�"o#��緟 8;��ꊸ]�d8ᡊ����ZE�8W���d8+�]&��j8�A�8�	�7b���]&�t_
�m{j8�~��Hi��̋8j+i8&�8�9��1�k�u��8u.c83�l81-���kh�&��\���t`g8�*�8qf�O����J�'8��8��[8�.���j8cg&�(�����N`p�Q%8���'����8�5�8K�$��m�*�8cb8�k��'8I��a�m�v$8�w�<r��)��7	���j8��d���@m�f���%���\ �7i��7�/y�8'���<c8�*��F�7�ȉ8�M8z����#8������g8"�8��煍8�r#8W�k8n׉�g>Z8���V�76o%8���7-*j8�!�7��h8m�8d	�8�j8�� ���98tp���$8�c8b�8B�j�O]n8�{l8���<U�	y�7~3$�n4 8�{귩�AT��=�8�L`8]Ng8��8�;��%|8ɐ���7E\���oi8�i8�g8o#,�߶"�^��7�A�7M?��跦3�7N�b�q��7j�i�$�Jj%�TD�y���X��"87�f��I߷���7f�'8 O�7{n%8dj�Q���t�&��]p����8qV�8�g8\�"�~��8L�����&8/2#���m82%�8���tL�8LO�8�8t�鷐�﷩84�d�&0�7�"�_����7V��7U�U2%8^��7���8x�8�Ԋ�O�l��*�7�b 8>l���$�v�8t�&8
3����7/��8� �7��8�����%8:���vO89~�8@�!����1�7��p8=o�7���e�7�$����7�;��&�����i8/zg��T�7�k��#j8�[8gcn���$�C�%8����2m8^$�|ˉ8�!!��m�H�'8�T�����7wA���6*8/�86�i��U8����r�7|3���7�Il����wy&�#H7ws���74E������D7�<��N78�� J 7|H��x��|	7��7 �� 7&���/72l���7��	7��7Y�7�'��� ���7���C7Ą �nA�����7��7z�7X72U7�	�g���� �g�7wJ�6^7{6770 �_� �j�7fp�� 7Du�	�2��������B7`M�G��~l7Ke7��7,<�w�7���7����7|���7����7�T��l��t�gY7����C���78J��7��������7ީ� J��N7�7��7[����7@7��7���P�ix���7@�7�7������U�&7	7B�6E�6�����7z��tU���^i���7h��t��6��7��7Ge
7���(7�7�[7G �X7r�7+�7�����7��J��
I7��f������7��x���#7g�����{�7� ���7s&�6|���h��x���J�6���7T~�6 �7� 7^��R:� �7�$7����Z�dj7�&7��Ȝ��1��� 7q�_���7W7���p�7*�7���n57�72�
��� ���7�[�U9�6OZ�6���68�7���77���6��7�B �;07�B�������4r���7�78�������7c7�0��9�7�P7�7������{�(1��37.p�FR7�9�g�7��j7l�6��7D��)��J���R72������Ћ���7pA7���U7�>�<l��c��z��'��������
��\�6G7-^�Ɲ��s��% ������P�7~�$�70�7F���/��"7�}	7d%	�\�������Y7l��Zv�H��6D��C���M7���^� 7X��L4�`7���6��73T�f7 �<��� 7q$����;7�d7&�7�5�f��]7:� 7F�7p� �N����I� �J�7�'7�� �����+�S�7PY7�B���#7>����7Zq��V������;�7����v���	7��7X�� �̏7�i�6H���� 7��� ��w%7L���f �|��ab74�:- 7����xv �4��k��4�7ӕ��ڎ��7�!�κ�6@E�=7P7��7EK
���	7����� 7g�6���7�7v�7 8	7�;�:�7*}��<7��7�`7���6@�7(r7�:7�7�W7�i��h 7Gq��7T2�6�� 7 Y�@�7r�7Qq������7(���/7���� ��H�?��6��7��7��7���VM 7��Ez76�3;7���6�7���oQ��7,.7Ѧ��l��%7����
7]_	��6��������l�n�7�@�����l�6�o7@�7�{77����(���5�7�g 7�	7X��T��L�;��t�	7ɶ��C7
h 7;����7�97b7f�����@e7���4X7��������	7��7����7�r7�p7�7}�~��+U7@�7�P�Α�N�72V7���ۤ7�67+�7T�7�=�B�7�$���7�7�G���X.7���6 �7�����7�v ��J7����l���/7���0I7�����7 �7�������674)���7�d��i7���z���&7^�<o7�R�f��6�B7`� �ˉ7��U7�h�U 72�^t�������_�K7�̶��F7B��7카7�J?��t�7Z�@�L1�7��;��@7��C7��A�����˲7�A�u~B7-2���?�7�C��D�ݮ<��|G��j�7y2I7�����H7x^���c�7�B7�Ĳ7�C�<���
�^����ݠ���9�7IvB7���7�P��Bt����<�%4���
�75ĳ7t���Ō@7����$ F7��C7HE7l!?79��7=�;�|<�7��E7-hB���?��@����A7L[��-E7t[B�V׸7�ɱ�η7j緷�;7b���l�>7M3E7j�?7]���� �7D7]�7�Q���7�uC�+�7X]�7~C�8z�7��7,����&?�E�A�I�:7�����z?��p���ʹ7��E7���76^���kI�cB���>7e;76�7��>�D�C��a���<�켲7�i�9�7^�|7�}�7vD�7�u��4�A7������m�Q�E��E����7��:�M�>��ѳ�-z�7��B����⛲�a,B7~p��6��77�SI�uC7�X�7)�A7hI���E7�r�7�����e�7�(E7�:�p-�7�{����C�M�:7`��76��7M�=�}B7Q�B�|ɱ�TA��������7�ZF7�7B�KC�Ҕ�7���7/�@��D��UI7d8�7➮7}��� D7@J7;�C�ڽ����>7������lM>7��?����b%�7�MD7��C����7�G�̧G�Č����C���71�B���B��Ĵ���]72���n��7��708G7��F7=�D�48��'ZB7}�;7��=��,C��x?75�I���A��ϵ�8��7��E7�7�@7���&4�7�:�;�7-����H7�Ե���C�:ڴ���D7ں?7��D7"q��H�7��7ݵ7r�@�������D7nK8�A�A7or;7��O7��B7�F7iG7��7�@F7掴��u���>74��7�9D7���7�C7=D7��@�z�7�ٱ��_V�.س7�=@7D�u�?�"̴7���7���7�l@7�)�����7��7�^��A7u:7澵�&W�7v���N<�7��C7�j����C��#H�ǽE7<C�7��O7�(�����7�G�7�I�G5G������mE7�޳7��C��bF���@�O�<7��>7|@7��7����@�V!�7�cF7a�@7�F�ڣ���3�7��F�?O�7�E��NG7ϝD7��D7�8@7����~�7��70���^۳��dC7�g7 G���_9��E7F�@���7��7~[G�GJ7�5I7��7�g����>7巷
�B7&aC7�?7 TG7�7��?�V�76bD7�}C��>�7ҳ9�lK�7՜�����g:A��n�7"����.�7���5�E�(C�7b�P�⡷�@�=�l/�7鵷��7�B�ꅯ�R���:�����	p>��𵷰3��b�C���7(��dܶ7�q��o_4������7��I��9����A7e�G7_?����7�&���8?7<I;7j�;7�?����?��@E�������;7����u�D7w�C���J7�;����C�u�B�:�I7��7U�F�_�D�̍|7d�7�v��u#:7b:���)B7WTE7 �7�7���7��7݉@���7�O@7.˰�aH���?��S��p�7>"�7�ߨ7��D7Mз��7@�Z��Ft�7�7��F7�l�7l\B�n_�7�I�����$j�7���>㵷�?7S�>7�fE�f�7|�B��F�7��o7vrJ�%����M�7dnI����Z�����<��H7`f�75�@���C��߰7��D7+�C��?���7E��Z����C��,N�
~F7�I��iB7ڶ��F�;�7A �7�;���g���굷��H7b����6�7�D��1F7���7Hw��޶�7ܜA���>7�ڵ�����\��7�B7jH?���E7Jȴ�QԲ7��D��&<7
Ĵ7�m���[�7�OE�J<?7P�:�Q��iڳ7a�E�bPC7�ܲ���A7,����C7��N75�r7",~���/<��x��/r&.^� /ʞ���E/ȓ_-p9�������/ο�-��n�:1�/!�N/�M쭽��ϼ*.jD�.x�� �*�<�z疯�KN���.ݭ�<�/t!�/(��-�܀/�ͮ���.h�.)�/����R/��D/;�/�f��z��������h��Vx-���.�v�ʇ�`{ݬ�$������ϯ��A/���ܛ�/�'���u�.↮��4��f���.G��.��R. ���X�.x�-�:M.R�گ���.���,9r����/:/�.��.]����-�����Y=0��"�Y���10�7���L�� /4���s��/s�/^�Z/?�s���>/]31/��o�ׯ��/I]�/���T9�P���ï4/V�v.u�/ Q�+�_V��j��Ï�?�/<�".#������6�-���/�0T0��xR/3kY���1���,�0`/\:��9��4��.�]����+x�¯��P�e���/g~]���ڮS*�܆/��Ɂ��Zp�.9�����G/R��.���i�/�ܮ�����K�J�- 2����"�/��/jJd.�D���ɭ��h_���3/��]/8*��\?/Eq/�n6/$��#�.�R�.����L��U1�.�k�.�M:��w�������'.\j/�l/����{�/�����Bq��0�BQ�`������/�/J}�/�T���Լ/���e��4K����/戞�`�*�g ������/'�!0b$�/�����a%���/�Pw-ղ�/��!/$�-�� �a/�A�/�T�v�$��n�8��-10'V���n"0��e/��q�m��/�t����/�+*/��=��;��=�/�}.Y�I�B�୏���8*/���Y0Z/��/8�6-0�4/~Ư0q���/�@����M+��e/�j�/�p�W7���c"�� {/�T���4>������/�J��(�~��S�/��6/_20˄o/���._
/P������/:B��'�/\J�.~PK/𨨭���/4ޟ�F��.�]D��Ǣ�"3/vѯ��/�/ޯ�e��� ���0�M�HL ���V����/R�A�F��/;��S�T.��ǯ"C1/��֮j���e�M�s�������/�F��Fz/쬴/@�F��pB��S���8��� /@���4�.����h`+.��'�~%!/b�]�t���o�/oO���s���[�/����+�/Ì�*��.��\/��/�5 %�N}/,����&Įay��?�/a`����>}�/�/t�f�Ȯ���/̂�/��/
��.��0��/0�E.�j�/�V	�LU���L�.bMn�h�.0S��(�/89����0���.��=,��/-{�/v��.oe�.Lx�-D�
0��/.���4M��}����.�b0�ϧ������-}�(/��D���@/���.��/���$/Rs������p�--��ή�=}/]ůn�Ϯ�jY�Ƞ/ę9����/r�m/�g."�/4����Qʰ�:��/3sV/�!]/��)���/��A/'j�/Օ</yy�	�m��e��w�u/W�-����e�p��8(��FlŮ���/)���/�ݯ�@����ْ/��/����Y{�/�*.Yz����կ�j�/Ւv��s��u�/�>���P�.�a60�<⯡�%0W({�� .��..��/B��.\��i�}��R���*�/�&��j;/�B��f�I��f�.�ә�G��/i3�.�}20��h/���/���R��/,E�/pj�-~����A���x�Z/WC[�R��t�q/,ow/�����<� 6�.Qo����+�,��\Ѳ��r5/�!���/fr���/�r�8� .D����,@ ��;.�dw�/������.V�G.s\���l?� ��Dl�����Uڭ@�g/4Nf���}/^Ǯs�c��\����Э4��-\T�V}�.�S/>ࢯ��u�c�58��4�]5��A58s�58n)5�8�58Y�68�5�k08�6��Q581�58��6�k�4�m�6���4� E6�y(5�Ak38�>6���88� 68�U6��6�X�28]!78�C78647�S78�G88�@68�#6��)7�c�5�}a58�4��;68N+78�T7�0c6���38��78�k1�;A6���6�O�4���68q6�NX78uH5���48v�88�58��5���7��P68�5���6��06���48rX7�
G6�_�68xJ78e�58d�68e�58-	58/�58��78P�68��48M�5�{�6�H18��78�6�J�589�6��W5���5�9�3�r7�2�68X�4���48��4���6�EX7��5��68V�7���48R�38�27�`O3��&68��58��68�58/J68��48x�7��$6��68;�78��5��O58�68,=6�$l6��678�P5��3�Fn6��T5�B�6���48��6�RJ6�4�5���6���58ܚ6��'7�!�68��68B�5���6�*6���48�/68��6�P�78�M4�d~58�78f�68�)7�M�5�� 5���4�G�58D>68e�68d�38�78���6��R78X�6��X6��P58�b68@6��78:681�78Y�78��6��*6�_�78A/68�S68�l88I7��6���58yL68�558FE7�:�68�b5�*07���68_+68_�28�S6��5��6���6�A5���18_y5�Vq68S68�96�T�5��/8�j�6� 58I68f�5�?N68d	48<�584�5�\�5�Ȥ68�6��6�9�78�75���58M78Dw4�L�48��58ۄ4��L78��6��668)'68�u6���68�f78zr78�-8�+�5���58�88$\78.7��R68\�6�t�5�tg5���58��48]378�'78�F78�26��a58�.78��5���5���58*�78��6���28٨78�7�?68~6���5��68�68��88<�6���38��48}�4�sJ58�7�v�48�d38��78Ef7�=Q68s6�[&68�F6�!�58�b6� %88)
4�6X68��58�e58�<6���7���68��48 �68y*6��q3��68/W6��z6��88�6�0�48�k48�48Z6���4�K�4��u68Cf68�7�Y{5��:5���6��7��68dQ5���68�~58L78!c78#�38[�48�_6��a��5���68�<7���58�h7���48En5��\68N�38߳5��958�58�5�|�58۲48�R58ä5� `88�68`�68�^7���5�l*68@/68��6�֋6���5��78�v5��A18��48g�5�V�5�c�4��c5���58�i38<�8��868L5�r5878F668�r5��5�A7�W�6��5�
P6��28G'7�7H6�868�6���58��78N�58�5�$�6�/5��5���58�d7��`8��<6���7�68`T38��38	�5��6��a3��`4��6��{48r�68"s4���58��4���6���4�6�s�4���6��7�.�6��E6���58S28y�5��L68��5�!I78��4��68�O68��28�(48�*78.]6��g8��4�.F38��5��48�Z58�h58�6�k�5��?48K�48�48�/68n-6��_6�ٻ5��5�j8���6��68P�68��5�l�48�58a�5���5�6d7��6�fA68"46�+�4��t6���48v�68{�78*�6�
�48��78G58B�7�z�68q5�97��Y6�L6��Y38�#78Y�5�G58�B68j5�r58��68�o78H84���6��&7��[58�78!,4� �5�o5��+4��68%68�F68�68��5�j58�6���6�I�58�u2�k6��78M�48�78K�6���48�U68k�5���68�~6��58o'58e�3�ێ68$�58�w78�68dp58��68�.58ϡ5�,p48���6"L���}8,�{�C{��=�7�� �H>�����(÷�����z�^�7>����eK8��N�s�t8��$���R8F�\�3�~8{_#8�%8#%}8�{#8ꖌ7��#8@�U��׷�dL��[�7��}���~8-tO8�0�"��Bt�4B/���7��$�J}8Aw���s�Q8��!��!�Rڏ��7��R8$w|��%O���~� 2�@{��9d8I�7~���}8��z8\�8�z~�sz~8Ew)�T���`S�L�%��l�7_��y�R��18n��7��~� ��������#8�	S�����MQ8��}� |8���7S@�7`~8�t!��iQ������Q�.�S8�a$7��~8�����M8��!8x@�7�jR�W�}8�h�.��aJ~�{/}���}�A���c4��S8е|8�!S���P8x-�7Φ�767T�n(8!�|8d4�7(.T8f������P8�1"8
�f�{8a�|83��7��Q8#8&y{8W=�7p&�5N-�7=n&8��8��7�1U�T��2\8v�|�J�7�#8�JM7C
{���G8��7w�|8T�T8W:�1�}��}�7ʠ��PK��8��(�@q8�z8N�Q��z�&�L8�#�!}�f��7IJ8}R8�y 8êS����7]� ��ؐ7vaO�Nâ��_"8��T�~����>8v�U��}8�\8"z�7�ER�"��דK��~8`�>6�XƷS�{8"�z�m�{8>��l����K�m}8{�7��8��
��u�R�|8�����P�$Ւ7�*|8U�r8�F|�>�~8O*|8I��'��7�~��|���O��L8//U����7�8S�#�|8�b�7���Ј�����|�́|�ʱK���T8�}�­R��M��}8lx!8�<#8�KL8@�8�oR�@��U�r��Ue�et��끷ğO��8�]߷v�M��R�$��7�)#86{�i�}�a�|8��7,=�K6O8��7�/S���|�����7dlq�qu#�Xl�7�Y8�ذ��uO���K8��#8�|��Q87:\�$����T{�\�7�C�6��T8ڋ�>-�7�T�� 8�	ො֐7�C{��#8P��8�R8Rb����7�Q8�|跸98"V�"x���{���!��~8�t߷�.�x|Z�8}S8Qn8}+ 8��|8V�P��c|8AT���U��}�Jy��_&8�Z����
8 ��7��]8{�P�"BG��]�7L�{8\P���PP8�R�k�n�L�Q8T'|����7��!�%��q�7:�{7�jL�,K|�1�y��g�7\.��~8�2~�֟|�h�Z8m'��}8�bV�0m}8�( 8�X�y�J�8�7���7/v8���6��u�s�S8}f!8�z8!�R�l%8�7�.�8�Q8�=|8^~8�~8�~8��L8�NʷHrz8@�Q�Nj8B��D�$8������M��~8u�|8��N����7�a���t#��S8ybs�`%�7 〶(��6TU���38�d8��M��H<8悟7�x8�vv���~8ь~8I'~8L$"8�""8�E}8�O}8��G���7��L8��}��'��\*{��N#�@�S��IK�5�R�?��$r$8 }��l}�6��/̷!6|8��"���L����74�7�$v��dS86��/IP8��S�FJ�7Vg|���7���|/ 8�A}8_�Y8�!8�N$8� 8&�S8�S���D�7�v�7Ԡ"8`|8!2"���7�}8�{8%�L�v#��VK8��$8Y�O8��Q�y�~��~O8�TR8J�7��!8�_S8�T�8��8��O'8�ˏ�={"8���s�S8��o���L8V�"8�8��#��ǉ�=����	P85k�7�O|8L�#8�}8�`S��P��1M8 �|�!lx8K�}�E�8PϘ��zv��%��^䷷h|�T�M8��7��T8�f�7�=x��N8Q�R�Fn��jYT� z(8��T8¶|�Q�!�N!o���鷖�~���9x�z? �DJR���A8�*r�z/t8��r�,Zr�EM��x��768���7�P;���7�1s�����V�7�q8��r��!s8Lr��[s8E~r���r89os8�<r8x�s8?������-zq8�)t��� 8~r�]����Gs���q8�@s8��8zc�7>��7��5�ze���ts��ws8H��7b��7~+s8A2s�%�r����7Q3��.�s8�r�؞r�y�r���%���u��kj8�P��8>u�ƍr8eq8�9t8�s��s8��r�֭�7��s��n�7�0���0�7��p�gr8�u��S�r�c�^��7�.����s�t��r8�s�l=s8�P���$�$�s8�Qs���r�C�7A�8~ls81�$�*�s8�w�7�yr8Wq�����x�t���r8<[#8���7r���r�z�q��*�7q�(8|s8B�q86^s���r8w��������s�H����r80����s8��7^��7Es8�����7~�s8�7s8
 ��#�r8PAq8p�t8�����98����x���1r8� ���d���n�ݽt85@t�gH��z�s89��z7s�?�o8���r	s8Fq8�s�a�q��[��}��7�o��9r8e�7Z�o8*,s8��s�I�q���r85��7�ur�5��- q8Q�r8����|�s�
I��G��7����y�q�x�7�q8�r���7��Q8��r��r8��s8t����q����7�r��r8��+8�$�7�r8u6n�Bs8�[�7��7��q��t8Q5�������iI���p�v�s8�k�72�r�9���Yt8A_n8H�r�Wxs8��s8��7a�����s�Xs�A&s�!�r8��s�[�G8RSq��ss8����e#�7���7���7щr���p���o��>q8"s�os�q>q��s8W�q86o����l8�@���q�1�r���t�cr�@�q�{�?�\s���7�a�7�p���s�����l��rs�'�q���r83���^d�78Zr8�����q�]��7��7�1��R:r�_Os�}�� qt8]M7�}wp���n8X�����r���t8~r����7z�t�97+�q�.8O}r8h�7l����Sq�54��)��7;�����s�Q�r8%r8�2r8�q��N����s8 S�7@
s80;p��o��Ir��bt��r8�4�7�H�b�r��3��ױs8�r8�2��\�s8�lt��Or8�s�B�s���s���r���q86t������?8��r8Lt�x�n���Q8j�l8��q�V�q8��m�ENm��_s8��r�����0gt�29�7����&?8�@r�W�r��fs��'�)�r�*�s81s�gs�8�q8�%s�IYk8�s�ƙs8O�p8@�7�Gt�B;8����]�o8z78R�p��r8�>s8�r8n�r���r8�����s8"�q8g~s8@�r80Qs8�ur8Uar82��7(q8=�s�W8��r�~�r8�9�7�@�7��r���q8A�s85r����g�7�r���o8\~n�l���1+��-8Ө�7Ss8XHp8B�r��%r8�j��w-q8:$u��-q8��r8�pr8|���_h��Os8�s8�p�bI����r8>�l����7�ss�.*r�!u���s�F�p��s�0s8*kr��o�#��7��8K u8��7yr�������os�i�s8Z��7�Ks8�q�����6r�s���4��7�����Lt8�{s87����r83Ur8��r8z:s�����98+��
�t8b�p�_���c,r8s�s8JLs���7Jbr8gr8|nr86�r���r�_�t8�r8����r�����t8+�s8Y��~.�7��s8B��7fNr88�q���r8�n=���q8H�r8�W��6jq�~o�7��7(�q8���`&r8�E���Rr8�s���r��Ms8}�q��8r8s���s8^��7��q���r�1�7O�s��r8�t��>�t8�����&s���q8�=t�6��7�zs���r8Ĵn8X�q����72�r��,�7�As���7��r���q�#Pr�3�8�wŸ_��8׸����O1ȸr��8����J8i��
_�8ڞ�d8I�v�8q�{8G���ɯ�8*�d�3��8l��;��8���85g87�8jƎ�<����8	VI����8�_���G���߳�h�8iM�89�8��b8O��8ʅ���Ԝ��Rh��8ߖ�8�Q�8�Û8��i��뎸�_�8+LM�vX�8�5���~���.�������T���Ӝ8"Ҫ��BJ����8�ޝ8N��8�"��HH�8�����t�8S���e8�>���R�8��{8�8Ί}�o���?�H�ف8�֬�һ�����d�J8��F��Ĺ8�Gw�=/ĸxW�8=�l�\k��By�8�Ud8|X�8�Jd��I8�0�8t	�8�����^��+��*�I8E/�8�3m8ޖH�,7��x���tT�8l6�8厹8|F8`T���/�8� ɸ�O�� -��_ȸ㣞8/����8�G�8o�8չ8�ai��Dd8�5�8#GG8>Ɏ��U�81z�8=�8 g��8Ɖ����٨�8��g�|�M��K�R�I8�I^��.�����8�X��������8	Ǹ/�8���8'�G�3{H��G��,�8�꨸�Ϸ8��8/¹8�r�8f���6ǝ8��f8����/�7I�8�8�֩��`J�=��lDf8�����0ȸ�\�8���8����V�8Ъ�8
��� �8��8�_����Թ�89LǸ�PH8�|�8���8���8�|��9�8<g8Y�8�g��3�8�m��
����Ͱ�NX�����84��8	jt�R~�$G�8B̂8���Z�8�|8uB�83��EX��_B�a����8�����I8I2���EF8�к�w�8}8*я8�����#��#����G8�ٸ� ����+~�=��8uʪ8��Ǹ#{�8�e�DkW��D�<�G��]��泛�����lc��P�8���8��d��"��A�����a��񹸾k����8K`��;n�8|��8v�����b��8�\�8����F�8�ȸ�����8�<���
|�*b8�oi�K{���JH8᷸�B�8�칸ɄǸ���8�G8�@�8њ��ⷷ�%�ɸ)u8�d����H���g8�J8�~8V��]ҏ�0Y�8Ym�8ڱ�8�|���H��d��\ӎ��D8F��8��i��C������؈�8/>�8�ߊV8 O���,F8���P���ۛ�PH��2�8Y:��S���\�8�Ԁ8u˸��ub����8&C8\e�?��8$?�4s���8�۝�����5R���Q�8|����	�8�⪸�R���5\�M��d�S�8�`�� y����8���u8�����8��8��8��Ƹ+��8�Kɸ�}8+��8� ����8vf�8�=I8[���(έ8虸�2�8-F�8?��81F8>f�84�C8��8��8Gw8@�����8����2��8b��8�M�8����H8�J8Q������ۛ8f�ȸ���8�)������d՚�W��8��T8
_�8*.�8i%��4h8�쯸�o�8�{����K8bF�8tM8�S�Ƹ���8���8�����?Ǹ ��8'�<�ݟ8��I�ȸ����������D����[լ8Q�B�󫵸2�8,��8ř�8hK�8��������Sa��/�E�G�K8�I8v7i8͘���T���흸�[�����8*j���a�8`8�l��X��8��e8y�G80睸&��n��8�_���q�8o��wgS�dV�8p֝8����:�8���8�e8��8�����w��s�8¹8_Ѐ��׫���8o�8�H��87��8v|�8��f8�����*�8�����$�8���8
%Ǹ�9f�
�8
g8]��8�Dɸ�[�8"�Ǹ��8J�F�+�M���j8n�L��8R�G��n�8�p�8�D�޾��t��8D2��g�8������I8�ͷ�o⁸���8Y>H��׺8#��O��8���8��~� �8"��BO�8^����8�eL������r��i�6����/�0{��wJ.�0@!�,���(�
���Q/��� ���|��/U�/�/9l/���/07-X�2��c/�V>�e͵/��6�����ȋ/��.d���j/�S���bS. ��.�5�.�>�.�󮴎
/#\�//�/�'�/!��o�+���0/��Y�'-��T�:9���ݰ�K9�.]$8/6�.�}��j��/�� ��k�-_J���,�f1�R�d.P>-����h'.R:N�//�/�k�/�!/z����X/;/x�/0��@��-���.~N���*߭o��.A]%/�_w�Hխ�
;����@L�/�w\�?���"X/#q(�v���1 �$�@.�/09@/��1/千/�j[/,.j�$$4�ӿ�/��t/(��-�Q�.|qy�k�V�Y�B�2��/�H0U�,�b%����L�H���0�/��9.R�D�۽�S�0�tկ���/@�Z,#�.*</焯'r�/.qH/P'߮8	�R�U/t�A/O(/M�P.Z[�.S,��+��/(�_.H��.h�*/�(�-
p/@�Q,`x��L����UI�|��.D�8���/�:Y��s/���0�-�?6/j�/��@.���t�t����/��b�$ �*\��'0�_N�~��^��/�f&0&�/Q��/�p���T'/����n���/6Q�/8�J/��-�8Շ/�ſ/�gV/bg��ӽ���.�qA.<��P�����.�%�`ơ.�9�/�Ţ-����� �����W��▆�b���s���b.�V/j񕯙?0���/��/\�.�<�N�4/����$/��m/����.|��-�p�.RDs/�@�?�N/�/W:c/�������.ǽ.�`׮�d�/�I��. ����,Hgk������/�/�m�."��/���вT��� �3�.�i�/x^�/�����_/��Ȯ�����.��®�	���׮��.xE����*���5�t�0�b@/�k�X&��]�-\��9�@��:Ѯ����>!�~{�/�/^�̮�( ��8�/`Rޭ�0K���9�x{�/&>̯�X㯊i�/w�Ү�_���ɯ�X୒+����/�2����K�/�#��(֦������/��#/��h�/q�/2[��~[/�Ԙ��^��"�/�<�.!�m�4�p�-S0/�g�/:��/r(�/����&.ԯP"�.�aC��v�ؔ����/,�z��0G������-�F��R5�/ QC��""�����Z,���.%K�/�}��q����.�2�H^�/�z�/phf-b΋��/���8/���.P���+b/�)/k&�/�S0� .B<��|�	y�/��ꭢ��.7#��%���R.���/d�.�|/�&/��0S��!0�Q��s�/�>r�4�/8��.���.\�/*8�/�2�/�5����Y.6Z5/��2-E��/'�B/�e/�{��u���b.��/���.$��p�~A/���.aY/�8/3�E/{x	0�FO�
�������m��ut���/���K����.�g讈(���ɵ.�6/���-H߮�f>/�B0�V�.p�%.A�*���-'�>$���M�/@Ӎ,�����ʯGy�`��.X�c.J��/0p�/���/&u�H�@��aˮ�e2�a��/;�/��{�����V	�/(�X.��Ȭ2@�.��.m׊/J�}q/®���.�%��yM�9"E/�6��g/�+Я��q/�/�H0r{���N.�m��50���~ �29��K
0XԵ-���/p��-��:�J����%����^.C����l�/��{��&?/��/��/H���y���U����	0��/j���.ﮆi$���/�u/.j�u��&.s��F��/�*��8ƣ�Ti/`;{/�ي.�٥���I0r�.l{Ϯ�eK/��?/��5��rį*Ʈ�G����ɯ�����/�_.\`�-IL�`���:��m/z�����/�蛮.��Z�֯~D��s8|���88<
8,��4t8v���8L<��o8F�8(|�$���L8>��D8H����8J������}�N�h8t�8�����8rZ�
:8��8V48���j���?���������8��8��86�����}��8�8H��H�8B���8��8��8zJ8��8���\%8<N8^��B�����ܝ8 ��8f�*f8� ��&8���8����8��8�;8���L8�86�8����80�� �8�d8���D{8�t8X��b���\�ZA8�,�^��z��r�8�8��8�H����R�v�8p8�F8H�����t/����h�8�&���8�,8�848V����8#����������8n��X�����8���4:����jD8�\�JA8��8����O8ҁ8ر8����88�/8:E�0�8�8tw��^8��r��2�8��8¹8�|���8X�����l�(4��8F�8`��>��R�8
8ğ�h���[8�[8��8j���8��8�1���ƃ8Z-��V���8�$�,���B8jz8,���8�e���֩�ho�bF8���A���pX8R��ة8!8��8�8Z��V�X�8��8H������8T����|��w80�8db8�98�#���8~��8>z�XH8Lp������8h�8rk8�����8n�8е8d[��^� �8�4��r8P�88 h8N�8�8N�8�82��v'��8x8r�8:U8��8��8����D8ؓ�H��^�8�h8HC�"G�;8DQ8�n8��8���:[8(]8TC��j8��8^Z�lg8��|]8�78ަ�J`�����~8:?8��8����V8,8�)���֍��d8��8$�8��\���58ܵ8�d8z8H������8�38�q8n��*A���8����8@e���8T�8��8��8�]���8��8nU�8��
�8��8������8C�ޮ8�8����8Ƭ8��8�z��8lC�b�8F�8�O8�?8��8���\8��8�m�t�8���X�8��`��P���8���Ƈ8������4�8�&�F��vX�P�8���,
8���,��F��<�د��\�1���V�6t8hI�d�8���(��Ȁ��8,�2O���8�J8���6v8b��/8�8.�8J���J�"�����<�8����8���^�8�J�X����tY8��8�&����f8v�8���-8R���8�8�@8ھ8��8�84��B�8�8�����r�R���8�8Lc8�R8�	���
���8��8<d8��8~
��8�j��H��.8L��h?����U8�8t���8�;��8��8�I����N�8����7�԰�Θ��Y8چ8D
�D���68�u85�*��Z�8أ������v����8\F�t�8�O�<��f=8xw8H[��4������8����88�/�T8~�8��8�)��=8���:�o8��82��N�8p&�\�8L��z88D��v	8����8^��	�^8���8x86l�2�8���&(8E8q8 �ֲ(ŀ�{��bGt��Dj���[�b�f��s�3������wF�2�� �@�>�L�:2�І���&��x�2��2����2�3|�e��o3�D�H�ͱ�S�:��2�g��3�Ҭ��m���_2�'33��2�S�0�l�2a�r3/3��
�y[;����M�3��426�_�ui����#���3�"'�ˏ=�<R'�a����(�2��G�ڶW�� Բ}�J��>_��zȲ�~E2�JO�ى?2���2\4�1/�2�z���B�1�W2��3�&�2�3��2��W33}l3��2�&�1(����e粡�[��*3m�$�o��X��1�]2%mC3g��3�ײZM�3M3J��.u3� ���`�2 �讂P_2-R���71O�1U�2�;O���3�uW3RW�2^�L����2N��2nī���2޺4����4hl1HO���e1G�2����U����2�:>��)�2B4a2�]Y���23p]��V3�>�2>02�β�o�2X���� �	��1�1d�83�>!�+�h�@P�2��G2�3�I�]Բ��X2$��2���0н��n���%�l��1��2i���2�3\��1�"�1g�1��
����?X�D��=���筱<"3�V531k�2�������ff�.@2x��2p����q�2���P��2�3e�K3�3Gs1�E���'���_3���2ʗ�2t���A���-3tf11hֻ��Z�2G��EAܱ��q1�L�1�����1 d���~���1@��2�!2�Y߲D|2�we��DB�$ {2��&2�=�xl�1V��2B�52Y�ϲ��زq�����j��lE����2"��2g~�2\/�JD�2?+�VறC0䲯�3(ـ�jŵ1-O+�b2Ա��p1���M{�2��0�-��W�޲`y�3x2����Y�f�i��0�2;��3�2���2 ��/�{���,����2�:�
�X�g�3h3�Z��uu�2\�ǲ-R��>[2xi�OK���B�2�3�����u{���>2�p2�����|�2��2����r��2�ң��U&3�ΰ���Բ�ӲB8'��Y5�!�˰�w51q#�|K2 j�2R�~2)(^3���22�1�22�S�-83H$3�(3��1�����s�F-�1ȉ�2�1�0��3�+�����3�#
3�;3�3�1<�2	l�a�F�J��?�y3�]+3�Ų^�r2DYl2��[��s�Xʛ2�����[�.�r��R3ӻ�3Lq27~2��3i4��^��5W��J�2�2S�8&S�~@A���3 (�,l��3��ò=�'�Բ�'�0Ġ~1$�l2�C���1�83XI��9V_��`Ĳf%��3셲���2Y�x����[�7���2��9��2(*w��,1�{(3��ر$uѱ^?r��/Ĳ�Ň2��?3<N3�3�5���,2R7,20��V��2�3gv3�U��'A�4�2=s��ĭ�2A�3nO��(�#�6���Ĵk�Q6y1�)��:���ܱ�ȟ2H��2�M �<�s2�ߡ2J녲P]����1�}3O�=2���v}���>�2*1���^3��в~�2�:2�2��3�+3::P2�~�2�'�'�	����2 �����P���Ų5d�2���2���=����Y��X�-��_�5�3 e�����3`�2m����
��ɲ�%�2�F�2݌2&���i?̲�������2Ț72�_3��D33z5S�D[A1�3���2L�²B�����0;?3*^E�rۉ3�~3 �2`���T3R�����2����hM�1`��18�2��ɲ���A~�2E�?�G��7<�2�Ւ��p�1�-g����b�2�N3�)��<�2h~�2��P��g�2�}&�l�2���80�34�P1M��X��1��s3��L~߲��r�m`j2���3 ��EF3����È��8x2��1)<2F3z��2ڝ\2�����]+��D,8l6 ��S�6��	7�>,8i�*�q7T��<	7(U���7P�6������R*8 �����)8\���17�z��-��+��%
�#�*8�i7�$-�\�7�J��{7�]
7dV7�� ��k����Ē)��{��"7H�7��+8���X)�2�+��W�V�+8�r+8��X'7�v��p7	,8�7|V7|7��ԭ-8Ĥ7�L�8��D��T7�c�2o-8<+�\�7�`*�0:7��,���7�M*��`�6��7X�7�:��|%*8��7��7(R�PL7�`
�},8ʪ)8���u+80�	7(��:t*���D9)8��	��i �@�*�z*8�17p}7��@��4W,�t7X��6�k7t�+���-�`w�8��`��6h�,���+8J7@R72�+8�b�x�7��
���Tx	����SB-8��+�\�
��(���+8x���.�
���+8LZ+�07\X*8H#��J,84�7l#7�[��\�7p�)8��*���	7�M7P�
�Zk,8���Hn���17\�	7��7�+�@�)8T���)�����z ��Z7|	7l�
�v-,��
7���6�+���
�^6+8$�7	7d>,��7r�+80&���+�܏7��*����,�7���������7`
7_Y*� z*8؟��-���`�� 7�?��t�-�P<.�d,8@G���)8o.8@�7�68���+���7�J7�X��ؼ�6������s�,��1+8(D7��7��+8�,�؟
7�`��7X���7�0,�D����+�xu7�"7Q+8 l��7�7�}7�A���-��^.8 ����r-8���6�N 7 ��6�C�6�7`�,8��7��*���R�)8"7 77�*8��7��
7D ��7Hy �����7D/7��-��
�0�7��6�G+8�>�6d��h7`7��(�vw,8|�7����z7T��DC7�;,8�I*�� �vh-���7�q�6�,88��7�V�6T`,����������6U*8����>*�b�(7d�7|�7@�+8���`����E7��7�A,8�e�Լ
�|+8����7�� ���	7��7p}7�}7l�)��7�,8;n������7b)8Ҥ+����p�7����6��7 ����>7��6�"+8T�)��7��*���*8$~7(R7|�7��+8Hu�p7P�7���S,8���`7$+ ���(��-�"q,8^�X4-8������*�Ć7�6	�-�0��|�7FA,�D� 7�d�h��\�
�<)	�T���.����)�(
��S� V7�� ���7��)���(�@�
��:,8|��/	��h7��*8 L
��t-8������7�^74F7�P�$T�h��lH�̵,8V�)�L�7T���6�����X���Y,8N�+8XT	�����6)8>�*8&I,����6|x�|+
7V�,8LE7��)8���6�e7��*��?7H��6���$�
��%��f-� �*8\27�B7x�7,�	����+�l�7��7t� 7��*8)��e*8p��0a����*8�+�l�+��4�`%7� �6O�s�,8p�H�)8H	7$O�L8�J1+8��*��l,��*�|����7�F7�*�D��DK7�R-8�c�����=.8�Q)��)�L��Z+���7����87��+��,�z,-8�\)8ē��Q+�#�*���*8n�p�)8�����7ȕ7fs*�$�7X���7,s �c��x�7�t+8��\� 7�-��,78������6���6���p�
7���7�,�����7p9,��f
7lS-���7��,��7��)8x�7�h=�?=8�?���<8�=8e?8�"<�c>8��<��Q98��=��=8�[;8?�<���=��k;81�<��<8�Z=���<8�<���=�>�>�<�@=89�:86;��n=8��=�N�=8��;8n=8�|;��%=���=��;�q�;�F<8�N=8x�;8A@>��t<���=�t=�>x<8$�;8v'>�e�;8*�<�ul=8��;80N<8Ws=8!=8L�=�~�>8�=8S<�V�<�M=���>8��>�Bb=85�>�44<8>�<�=8��<��<8�~;�R�<8H�=8<8�>�x�<8
,=8Ѻ<8�s<�F�<8�5>���=8Mx:8!�=�g�>8��<8*<���;�Mf:���88��<���<���=��[<8z�:8�n<8��;���;�#�=�&�=8X;8q�:80�>���<���=�V{:���;8*=���=8��;8ȷ=8�;84�<�S�<8�Y:��/<��d;���;���;8��:�\�<�X�<��=8�F<��r=��(=��=8��=���<8M<8�=���<8�;8V�<8�=�>8��>8c�;��z=8�h<8��=���=8�;�\�:�d;85(>8t�;8q�=�6�98NW=�Lt9��>�A�>�_E>8=8C;���;���;8m�;8�:��@>���=8�V;8�}<8�<�S=8�J=8��<�l�<�,�>8�T<�8�=��<8�<�g�<���;8�X<8V�=��<8*�;�F�<�lc;�L=�`,78Tk=���;�Vt=�:�;8��>���;8.>8c�98>�<8.�<��3>�%�;8�o;8��;�<�h�;8��<�<��v=��e=8P<8�<8G'=8T�<���>8 �=��:8@'>���<8\=�@W9�<���;8&%:8�d:8q�;���=8�=8��<8=�=��E;�U2=8(�7�h�>8�5;8;8<8_=8�}<8�>8�<89:��J=�x�;8��=8`!>8�n:8��;8�,;84C>�h�=8��=��G;���;8�<8�,>���=�2�<8#:8V<8�	;8�6<��#=8^�;8S`:�TL=8{�<8%D=���<8�;�)�<8�b=8߈=�=��<�s�=8��:8a�=8E3>��<8�;8��;�&�<� !;��2<8&=8�H:���>�w>>��98�:8��=8F�=8��:�&�=���;8{�<8֖<8g;���=��;8��<�ê=8^];��f=8h�=8�|;8��;8��<���=8�I>8�<�^1>�.b=8�88%�>��^7���<8�j<�D�681b;8Em;���=8N|;8�=8'X>��>8u�=�I=8�T=8��;8��=8�:8��=�#�=8��=8�A<���=894�v8=8}k=�i�:��W=���=8�i<�k�<8��8���:��y=8=��X<�Jg<�H6=8T;���98+�<��S;�֩=�+n<��>���:�l�=�XG=�v�=�:r:8t�;���<8��<��'6��<�l?8��=�Q�=���<8�P;8�)>�{�=8r�:���;8��98Gf98@�<���=���;�;p:���<8�N=��>8��<��;8��<��D=�=�;�m�<8,�98��:�_�=�w<8FE;8�=��38�B>���;8�y=8��;8}>8�:8@t<8��<��:8��78.�=���<���>�}�=�J�;8�U;8N=8<�;8�=��=��=���<8��<8ic=8'�<8Q�=�+=8d>�g�=���<8i�=���=���9��=8f-;8��>���<8�=���:8��=8}<��b=�:�<8ܿ=�?>�e�<���<�G<8I>8�1=���=�x|;8�>8Ka>���;�E*=8Ұ<��=��1=��s=��<8a�=�
n<8y;��<�P�>8s'=8;�:�h<�F)>�T�:8��=�tJ>8~�:�!�;8��:8�=��!=8<�=�.�;82�=���:�I;8�7>8�=�2=<8��<�|�=8�?�O�78�D=8&t>�V;8��;��9>8=�4�8�j:8�;�B<8+�=�&�>8͡<��1>8N�;8I�<8��S/eQ.$	��D7Ӯ.���®X���f�Y/�i���!����.���.5Ѕ��h\��s�/B�/Y/�R�bE[/�����>g�.�������6:�.1Ԗ/���-R���U/,��/
)/$욯X��/���/���/�n�dVO.;$K.�ƨ/A��.�Z�/.��.�h��w��������#/ /./�/k_�.L?���ë/�Z����/q[.��E/z��-�G��?z��Q���R�"=�.�����m/w7�.���婃--����E/-��Z�/��z�dgJ���G/�az/[�Ю�ᆭнI/�a*�f
�� .06v+-�L��74/<�&�3O(�2��/�D7��D���K/�(_.�9\���/�`/�F�.ǆ��0�T1/O�,���/yݒ��
̯\��.�؁/�}�.���.`�L,�舮����ʁ�-߿y�-.~�n/� ��q��T��/��/�ȳ��YC,�Ń- ~^.�/����Q��.���/��,�"B�f�."������.Tn﮿���յ7�[ʘ-�6y/�~<��_/5M|��E�Q�X/?����9��d{��Je�����J~�c��#�,�F�.|_�.�l/rwg���t��W��%�.�)�-�kʭy���+V!/߲<�\<�.	}����+�Ⴛ��'ůx�9�������t/�B�/��-A�@��3�/ H�+^��-�p/D��2 #�%S�.��M���E��Ϯyy�^U.��n�V!�.��[.N�D�	�M˓/7/�G��p��o)ӯ�"�/���/���-��.:��.(�x��Hy�	�(�J�/��/	�#/}/��p�28#/)��,ە."B/˪��yj�{h��>	.�4���-�ڮ0���S�����殎��-��=/�\F/f�.?Z�/B�-�f���®$CE/��1/���/BS���k.n�T�j�y/D�.f����J�.̠/>�-/�|��7�/$���6�1.��ܭ�Î�&��.��/��n��?��r�.����Hg��;�/m9�HlS���~.�ܓ/��Y.��:�v�J�,7�Qv��n���ۤ.*)�����/U�|��r�|���/u\V�:��[�9-�/}>��#I�H������/#V\/�%/-�s��k\- ������-tO�.5�/ l�.C�������m'�ПL-*E�.��/"aQ��Z����Ag/������	�t���򸳯۠ �g�s��>[/p�^�F/�e�/�����;,�5�-c[S/���)�z�Hb������i��� u/�#�(�&/.eA�L�	�+�2/ޥ9��Q%�k-�a��5�-	�[/�u��'����M��P�/cj4/+�����.��ٯf�0����%���.(�G�5/z�/�)3.��/V�d .�t����t�/M�/�
خ�dA.��/�d�.Uq.�A�͑/��k�P��/�/�h����/X�q-"��.���.�//�lJ/X8-/�L:/��������c/���.��\/oK���r����2ϕ�nn��K.0Bމ/X.*/�.��-/�˥���x�*�0��r/�1.)��-�	=/Ș$�S
$������E6/�!8�S�.� �:�IY� ��-X��,:}%�lq�j懮�/ }-Wyj.O�ϯ$����%K/�M� \(/��$���-Th�x6y-Ά���̒."N�-\В.8�����N�� �/���^���R�(/.�jC��0��b5//r��8j/[2/���/��ٮM>�/V6I/�a���{�._��.Z�e/�Aح=K�.�20������.��.梆/V+�-��Ү��P/���.�M/�����\-]�0���/2��-&/0-�.j�"�Ak��k>�������.2YJ���/������/��I��}w����.����KW/Ё�x7�/��/ʓ��ni���6.p �f^��*��-��
���Wa9/�U/�Ю��"5/�0��G?����Z�y/�:��4��- �e�vZG��}⮌���hҁ7,샷lu{��{�7�h�7��7P��7�m������h�����7����� }�ǁ���{7>G����|����7�^�����D�7�>�����Da}��P�d�z�t��7��t7�v�7�Sx�d̓7\���!���0��Ё�J���7�}7nN��̇~7��7�I�7��~��ր7���7�?�7x��7;�7�i��NT�7 �����78q��Ҟ��Rց7���7���� ���h~����7�}�g{7�7��{�4�y7�������j̀7`ꀷHv|7�*}�\~78���H*��*��� �~76W���,�7LO�7�ր7�}|7��7�b���}�>샷�J�7ȁ���P���V��R�7�����X���Lx�|5�7�l7����h�74�������^��JA����{��J�7N؀7���|+�h��$��7{����|��:��d����+�7숁���~7���>�7��~�L}7�C���L}�0s~��L|�|���<�7 ����|�lj7�'���@��(̂��߀���~��s��Ԉ�7�7L`�>y���5\�n��7V����ڂ7r���{�7p���Ԃ�J��7��7��y��������7��7� �j�7X(�70�z7��|���|7Hy{7vk�7R΀7<�~7�2�7�1�7�����V~7�&���%�7�v�7��F���z7l6}7H�7�����%���7��~��~�4/{��x���Ls���7�܃7��76��7@V|7���X��7�+�� �7�T��ޡ�7�V~7상7b〷Ο�7��7~�0�{�
5��l�7�]�7��7�������p`��3�����7�փ��.�7K��\+��Z�7(�{7����h�7P7u7T7�i|�d�����譀7\)�7�^~7���7zn���Հ��؂7X-�7d�7ꯂ7|��7�F�7��}���y���~�Дx�0������7�8|7���I�7l�~��������76��h|�7P���0���@�7����8�7�j�7�$��&���j^���7���7J3�����7$}v��7�7
E�7�}7(~�7�n�7�����[���<z�d�7\�7�-�7p�}�֏�����F���8x~�Յ7`�y����7H�7��7X���p 7�y7��7f���=�7�d7�L�7�L�7�Ѐ�(��7lx��P�|7�|��;�7�A���ς7n!�7���7R<��pf}7���7΂����7��{�|�|�4���\V�7@�}7}�����y7�z��w��K��jk���_�7��78�|74�|7�Yy��)��&Ձ�Xrw� ���|��7 K�7�΄��I~��o�7�����Q�7��~�x2�7�N~� O�7\�|7��7� ��`<7ܵ~7��7��y�@��� k}7g{7����\����}74�}�|Gz7�倷��y7�u7�u�������}��_��H�|7(���X�~��m�7�o�7<ς7��{7T�s�P7x��H�����7�����7x%y��U{����p�7����W�7dt7�a�74O�72���ʅ�p��hz|�j9�7`�k�H6~7��������:~��8��:���|�7�܁�@��7��7�Ɂ76B��(�~�!�7|��7��7,D����7Bł��~7������h7Dp���́7�؁��Qz�6���zp�7���7ĝ��P�}7��7���7�P<}7��7��7�7*��7��~��f����}�H�|7v<�7�~���{7����4<�7��|��&���'����x7x��`��N��7D7��y�ʭ��'p�����3��0��� u7p7}7�ك70�7x�|���h�7w��7�b|�X�}7�ڀ7�����~��"��Z���S}70D{7Dxl�|�7�Q��rP��@�y�4ԁ7�+}� \�7�Ճ�xD��概7�H��,�}7@x���7$��7���7@���TB�7L'}7lo�7�����W��J���Ю7�|z7�i~��7%� 7��#�a��7!�޷�3巘�$�>S"7�x緧�7��۷�s�7�|᷏��_��7%��7'�y��7B�+��7��ݷ�7��&7U�"7Y�7�u$�|߷��7��޷�%�7mA�Y�ᷫt��7c��7��7A 7���7�p߷+9��1!���7�#7� 7���7� ��!�T��7z�߷Ld�7:N䷉���්c������7т"�V��5}�7��7���7	�n�7]j!��~)7�6��-#7�p���$7��߷��&7����q߷�޷���7� �S޷-�߷W��7to巜��7���� �w��7�=!�i`ݷ��7��$7*�7Ve�P�7G�77��iS�$4�<��7~��71�7�O�w����۷�%7$"7���7>��7����!7 )��u߷0o�f,�=[�7�@߷���7���7�]�7�d�7��"��7�z�7<��7�0 ��G�7)b!7]�7H2&��\'70߷�,��=�7},��߷`޷k��7�M߷�%'��z7]�ܷ�F�#��7�/�k��7I��755޷K�䷫���7M�!�S��7�9"7fc�7S�7E{޷>�޷�r�7s�!7�
�dܷ��7���7����oݷ��ܷ�%7[6߷x��#_�7i!7���R$7�Q�7i��i)�7	��7��޷�!��q'7A%��2�7�Y�7�1�7��7��ط���7.� 7z7�&�5�7����� ��"��r�&�7�u 7A^��P෼��7sR�7Zݷ~<�7g��78J#7�#�&���ݷ��V�&7a���D�7�'ෑ�7�{ⷀ@%7rF�7��7�$�G�A�����7���~�A߷��7<�"7�"����7��(�_�MNܷD��jz�'�㷯V'�c)��740�7`j!�U������F�hv޷�=�&��7���Z�7�\�7�z޷�߷<%7A�7����߷�� ��B�;��7�����;,#7R�!��ܷ�O�7�"߷�=�7��߷ա���(7�4�7Y�7��ⷥJڷ>P��B�7��ܷ��޷�7l�7H�7=j���9j�7X@(71��7�ܷN'߷�kᷩ� ��%�7�]�7b9�+��t�!�B��7>=�7����{�7^�淹R�7]�{Cᷖ ޷�l�<#7��ݷ���鯡7�r�7���*���a'7�f�7�ݷ�%�7x�ݷ~ݷ�j�7af޷�pݷR�#�17��㷚�7A'�
�߶�-�߷2�71�7��޷C����7hg(�g"�7��ᷓ��7Ƌ&7��"7���-��76�X]�7��$7�Y߷�N�7�Q$7��7��X?7Q޷���7�!�7~A�7	��72l�7��7�$7�?�7�r�7Bw��7t���7�<7���7���͐�7R��7x�߷ �!�n��7e����7�ݷ��۷�ݷd��7Z��71��7Wi�7�����7z�QJ�7.�I��7DC�7u��78"��V�V��70��78�����7��ٷ�v�78>�)����ݷ��$��Xݷ�(ܷ �)7\�޷_��<��7���7b��7�57%�$�q�޷�!�7n�OE�7\F�7#7�ݷ@�޷��ݷ�B!�n:�7��"�>=�7a��7A�#�.�7�)%7�#�7��hy����7Z&��%�7��r`���7C`�7���Ge(7TA'7��7,��7��߷k��(j7��7���>)�<��7�6�7%�%�=� 7-�7���7)�$7�q߷��7"�/'7ж7�r#��y#��7�5%7��"7V �i�7.+�YS�7��᷉~ܷ�H"7I%ݷ_�7g���/�7���7D�ܷ�l&�e��7ɞⷕ$)7��߷a��7�Fܷ̗��;�7xF߷e��7��!7���7d�ܷ^�79R���7�޷ª 7K᷾��zݷ�n6��'8�wJ�&DO8��I8���Vh�8Ԧж.�q80�5+n8�zP8��p�6�p8�CC�.�'8�dO�hU+8��J�|8M8eDP��*�b�)�yXK��t���zo�(�P(L8�e8��G8�*p�,�L8�O��H��*K8Ϋ�8�rm8胜��n��((8��L�gI�8��8�K�̇,8�&8[om8)�o��1P���J8��(8��K8f���0J8�s*�����:�P8��N���F�)O���L8oM�9X&8h�8�L8�8PYp���8%J8�K+�z1s�w2M8}��;m8�����jL8��M8��I���M8��M�0팸�Ɋ��DK�ܑ*8�K8��o8�ow8�aM��`۷��N��l8w(�@2���Ao��L8�M�3��7t6�8b�K8�2Q8Z�M8�N�8>��7�^F��O��K8�<)�&��No�=aO8�@���J� o�b�J��!o88+r8�M�/�����8��K���K������L��S$���O��]���77n�����1M�������8E�:8�N��rJ8s<���,�@�T��L8�	?��ߊ���K���K���K8�nM8|�o���8;|)8a�I��B�8��=��cL�]SK8G�H8��F�f��8bJ8�{m�v+�G~N������L8�o�p�8 Gr��a,8l�k8��'�	�K8���8�Ġ�d�M8*qM�*N��Qm���L8@[�8�(8pM��i�7S\q8�M���M8?sM�Ǆ�8�׉8�+8�rI�`����͇���G7.C8�N��Ҋ8�eM8
Qm�TIL���>��HK8,�L�P2Q�]�8����0�K8�J8�h)8�#�B�L8"%��L8;�M��Il�0F�8\q8zC�8�O8�M8t(8��K��]M8��G8A=L8�qK��&����7J��6���M8=iK8ԪN8�cN8��F80�϶�M8�	�8�*k8>�&8�LL8t�p������O8�O82�H�l�p�(�r8�lK�X3s���M8�1�8�!q8�q��&K8�Y*8*Tp�5/N�$�����F8�%�e狸��J8��I��M8fIr8�7L8�0ɷ�ͨ7��L��)�8��o���J8�Ǉ�6�r8Y�r��YK8B<'��eL��L�5�J8*��?zL�>"�8"�K�	.N8�D8�'K8�)8�^M�z�j8��/7��L8(Y��<�L�W!M��:��]�K�9�K8��K��K8�6L88@L8�M8��(�)�N8�8���
/�yNM�SrM8L&8۰&�o�L���P8*I�ߠK8B�:8iWJ�5 N8�s�8*8�y�8Fp�4�6�/&8��H8��O8�V`��/(8��O���M8�WM8X�O�l�(8y�O���K8��K��"(��8�U*8�=�6:h���E�J�D7��C8��L��Q*���J�r�N8V�*��Wl��gL�I&N���J��?M���K��M�g�*�?�o8}�J���I8��ѷ�N8P$)����8�Cm8��&8ѱL��N��9K8D䉸:�s8�''8��K�g�A81,p�n1j��l7v�l8�JM�WkI���&8(�Io���C��O8ԸI�@>I��J�����X��N;K���N�_3!8nH��6�)��K8�il8%�J8:u'8�5K8��'8
M8(�M8�(���K8>N8nu8��[8�?L���8P>$8o��7p�3�K8f�M�&-p8�a*��8N8n�l��EM8�n��9�m8�$���K���M��b��Ȟ(�c�*�,�L�<K8��r��\6v@��7�L��+8�Dn�L�J�v�L���'8G�8Fv'���(��-P�YK8?L8�N,��:M�	2n��Ӊ�0�K���K��І�uV�8�)�@Dp8��&���N8
Q����4<�*� �'�>���v�,8��n8�J�88�&�$4���I��Ɋ�"�L���N8ЉK8��*���O8�F�l�O8�K���i8��N8��(8:�p85~O8>(�tbo��UN�D a��M8��G�9lN8��o8ywN8^T(�:\P�7
O8���8^K82z�8a�L8��8�G8(�'8�O8TO6��,0��0X%1g4�0�'�0�a0�՜�@]:.�QV��H1�44���|1@J�-@u�XW�������15+�0�_���D�D��0|��/C �*1� N�-��h/>��/�2��j^0���0�,��@�h�,� ��u%19&y0{�0>���G61�����[��|�8�ʰ�A��/�/�0@_a��=0�\1��1Q�1�1�0)�0<�����/X1 ����kڰ��������e0P�$/��/%�0����0� 1n10��Ȱ ����{�#�h�Ԃ�ƺ��r�/m 0$��0���0����g���g�0�/ĩ����Y����0\9u0j��/?>1/�c���:1��0�˓1İo���\��uR0�2��Jo1	���W0֨�0~���uְ����m�:8N1X敯�B)����4�j�c�0�0���q���v/���0~#�0Zy&��I>���0���h�5��'�xUݯ�b
�e���1��+10�-1��p.(�/����|{R��/��~���/h��/UɰaVb��m�0��r0�\�M�>0�kg�hf�/,T�0/��@�.���=�ް�\�0�'�0�P��֦��	J1lߛ���/�f:W�N20��/�,/��z ���41v�d0��V�fI)��|�1�(S�a��7����t$1d?a1V�31��/Hܝ��?���0(�����U���Ѭ�B�.���)0FM(1��w�w�p0B�0�̰/ɰ�N�������q���(�0V	�/F_�0����j1��b1H@�0��0މ1T_���g�0�Ji�7�r�0���-T��[50����$��0�J	1c��0p��H�C�,�Q�m�
1��,3��0���0o��0�J�_��2��0l�7/o�0�"1�;D1v�1 �1 %1�o0;�4�����Jl�0��6��	���ӯn�11�ӑ1��Z�-�0�C����"G��+o�0�<V� ���&�[���޳��!0���/鰅㈰��D1������/���Dװ$|�1���/M$���Q��]O�d�#1�>���!0Z�(��旱2Ӟ����08�2/�)Ȱi8�0�ǣ0�&r�lg�0��4/�
�0������ް�@W1y1��#0H)�Y �0��-��b-0��B�J�0^0�"����"0.%R�~��1���ڮ-0����ư��ǰ��@��h�/�1�j�/�0(ƨ���1��`��l�0G�13ph0k!�0�?Q/�?M�[�$/��K��C�l�/�h1
��0����wo��~�HO(0:vװ�@,�������������0��1�;1�ӥ0�=0��A� eK.�+.1��'0���XΏ�@Z#�����ʅP1[謰�τ/��m0p��1�0/���0��0y E1M�5�`0��010�/�큰-=��c1�C30@�`-$�. oE����:e���0D(�0�m�0����a.�ʭ��*�w�����#1�c�/�0��7��9��`�0Z���������0.�-1 �X���X��[�0u������@�Z0D��0�LR0�0�A�.�ư�4g���0t?�
l�/P׮v���3۰����"Q��0q,21hů�Dt����/>��/ߓ�0�uq����0
���`1�H�4C<1<7�/�	0�u��)71���*��0��J0[=�/�c1��2���o�9 �0G� 1E6ưlD�/���vo��mw/ƾy0�m�0��ݰ��1I���&�$��X�0~���1 eU.\ê/ ! �	H��j����D��t=/���2���ݰ\컰t��/��a�pkV�>?0v��0�0?.z�0�Ys1�0��E����0�|�􀨰k[������h�Ԩ�/�ݢ0�yJ�J�0]����Ձ�Y�/��.1��U1�ީ�`�0.b��d�0�2�I `��t[��;//A1�:�T͡�I��1�61����Ba�����0(VT0��-<�u���'0�D��ג8�����8��*h�S�ь8Rc��8�4�Ŋ8�������8��8i��8����8���8��8	�8`8�����.8����58���y�F��38��8�>8tI8c�8Q�v�������8׿8�8(8��������8�����8��������u�����8]B����� 8�8��8��|�8���#f8�l�U8I��M�8C���8N�����3�D�8����l�����8T��]8(K����8a��t���8
f8��8V��4�8�K8y�8��?��n��aC8�,858�;�F��X����8E�8*G8��8���28�/�iF��^������8��
�8:�8M8p[8H3��:8�{8��8�����8��8$C8��?�8��������8N���c�_I��F8���2��8BA�E���8�;�181%8���������8��P.8��8��8�86�����H8	8=�bp�S8�a8֩�gY��D�z�8�u�����8)I8���	�8��8l���8��8������l8��z�8�8��8�D8ا�0Y8	�8[8c5��I8���������I�@�85280��ٱ� �8�$8�l��V8�8�O8��������Z1�[�8���K8���Ct8���J8��8��8������&�b+8�Y��;�+j���8�8(��o<89��w�%B�����h���������:�8�8�P���0��ڧ��4�L�2�8�����8�A8(c�G(���8I�8<��9��?�������8��M��~�8"��G%��38�j�M�8D[�c���8�\8�a8H��������O�8>�'��\8\Q8ն8�_�֩���8B8��8����h�Sb������8�-8������&/��8�
8����80���{8���zH�7/�y���8.������~85�8 �����;48��8���M78��Y���8�E������-�8���!�8�h����m�7�`��
O8���ZC��8���w' 8����8yq8��8����E8x#���8��8qg���8N*8f�8� ���8M���J8��8G�8�P8��8��8FC8}�8�(8�Y���8�����8�8�8b����8!�8�������.8���8�C�2\�����o8�@8��8�#8g����8c���8��{�8��8�%8@N�u���8mj8$��\]�ͤ8(��	8��8��Z����vg��'�D8���t��\*8�Q8fQ8��8� �0,�j�����F�8l;85M8h��/f����37��68����X8�=8���N8(�8�
8�`�E��8Q����8b��s����8�8����K8��8��8|�8��������8�38k��|E���8��8-���8;�8�H8zX8�>�k�8�"��8=�8@���V�o�8�8:8�:���8����8A��@�`;8��M�8���`�8ڛ8������8�����8�T���8 ��2����8�?��U8;��v�8,8����8~���8�_�W�8J�����*�����A�7
m�ڈt8U|t8�z7p��.�v8{�s���j8�m�T�o8"�p8��n���q�l��7�u��5�7��t�,.p8VIn��ӏ��d��o�n�<ހ7^vr8���>�o8��o���m8��p8e�k8o�q�ƫt�dpm������o��On8x�t8�b�7t�m�8���(8����p�x�y7��7"hp�hq8�<n�҉p8'�7�t8os8�"s8tIs��>�7��s8Xmp�~�n��p��j8��o�xa~7?��L�u8L���9�s8�ʊ��Uq8�����o8!�t8
p8�~r�ܧ�7��q8��u8�sq��p8�&q�(E�7P��7F+s�`�7��q8�q��a��zv���7@fr��cq�49��,z�7�yl8��q89r��ep��9��`om8��o8�p8Д���ꊷ-�q�%�n�w�p8�����7�kk8�.v8�3�7
s���l8l%u��ar��kr��ir����7F����q�U=o���7�s�����Sp�T�7 _��)mq8,U�7�p�hO�7xUs8ޖr8�s�u�t8���7즁���p8՛q8.�r�h��77�t��!o�]eq8]�n8�jp8�����Kz7T�r�$߀��^r��ws���r8p8�)v���}�Ws8�s8��z���q���7��t8}Dq8<�����o8�jy7�wn������q8����qs���p8Z�n�n��p89�q8�1��x�7��n�J�p���o�~tp�צl8�l��	��<	��8�y7h�r���7L8�74�q8��t8SRs��Un8�vp8�jt��w��p8��q��m�$��p��7��s8�'p8�w�70@��P8t8�q��p8rLq�Zs8 ����l������n8�n8(|7�q�N�t8�?p8�o8�ir�h:���t7c�l���~7�Mu8\�m8�r8�m8{7p8�Ս7��t88#���vq����7}�u8��s8(x7�Ir8DDn8��s��Cv8Ԭu��t�2�q8�.q8�Ȉ� Ju��Ss8�op8�.�7 rn8Fu�2Xr8g�p8H�u��2�7ֆq8pt���r8��o��q8�̀7�	���Vq�Pڄ�qRr8+8p8t��7pCp��u8Ml8t����dp�Lt���o8Ȭ7f n������Tt�!�p8]	p8�-t8�_�7�zq��7r� #m8l�q8 �7bbp�#�s��
�7�q��Ru8��m�&�p8��t8�go8lm8܍���,r8,��7>N��Wo�8Yn8Ȱ�7p���\�k�d�l8��t�g0j8�	q8F�t�bys8��n8��78+����o8���TՇ7}'t8Jq8��w8<�7�
n��i8
*r8�eu�À7m���s8<.p����(����7`�q��O�7�Fp�T��&�q8@�m������nr�l�n8t����j8p�m��s���o��o��q��k��m��8�o��Fo�P8u8_lo�vq8�	��Lȁ�p�컀7�vp�Arr��<t8�_�7"�p�@A�7.zq��}l8��n8��k8.ct�۹r��5q�.�q��v�7젉��p8��q�s8��q���t���o�0��7�'�7��r���p���7xP}7���q�h83 q���t8��~7F\v8졊7�im8�q8�!��Z]m8�Xk8��r�f}p��6q�\@��`;�7��u8��r8؊p8 <s�zVp��-}�x�o8�r8V�n8�7u�`�y7ϧu���q����7@p����y���o���q8h�p8_�p�� �7v�t��y7�o8�'r�NFq�܆�7��������5��Ho�2m8=�q8<���t#s���o8��7Y�p��}r��74儷�扷��n�0+����s8��n���p8`1~�4n���]�7ȩ�7@�o��7������<;�7��q����7Y�q��4r8�n8􏊷V.q8߼v��Mp8��q���k�~cl8Ȏ�7�p���r8tك�-�s8��r�l'm8E�o8|�n�1/s8��t�N�r8��TEk���q8 Ԋ���q8x����o84�����r8M�7N�r8j[���b�8�]��T$�8D�8��8�����8�ָK��8�����;�84%�8J�ָ��ָ�ن8y�ָ���87��Vq�8t�ָ�;ָC׸����:��8���8�S��	2�8↸���8���8���8�}Ը`ָhZָKʇ���Ѹ���89��8���8�7ָ�>��p�ָ�톸���8�݆84d����8�_׸��8V�8�k�8�b�8���8hָ=��8�G�8=DԸ�Ը��ָ�l�8���[�8��ո�a�8�
����8�Q����8��ָ���8���8��8��ո�e�8���8!�8�+��:=�8|���j��8�]�8�|ָ���8N��8��ո�����׸�L�8�?ָpK׸5�ո
	�8�d�8��8|׆��ׇ�t���$e�88��8���8;��vp׸Sո�>��x�8����;�8T}�8H&�8�`�8�rָi��8�����#ָrU�� ׸��8����ո�ָiÆ8��ָ9�ոFԸ�r�8M��*�8�{�8?ո���8���8.#�8�vָ�D�8~ͱ8�nԸy��8.�8�ָq�8�Ӆ�����2�8��8�Y�8I�����8�jָ�Ӹ�����Cָ���8�i�8x3׸?������8sS�8�Ը��ָ6��8ڎ8�&�8XMԸ�T�83��8E׸���+�8�Q3׸VQ�8^8��V�ָ^�8�,�8*�ָT��8�߈��؇�n�ָflո��8`|���j���eָ@=�8Gø;�8�X�8J�8S�8��� 1�����8!k�8fiָtc��Cr�8HcָD9ո.L���v�8���8��8�M�8��׸��8��Ǹ���89ن�&;�8+����4��Ԝ���{�82m�8�ȅ8ḟ�vf�8�v�8ጆ8ͷָP������8Χ����8���8-�8�-�8�)�8ܯ�8.��8��8�@���׸�1�8���8L?�85˅8��8���8��ָ~��8t�ո\�ָn8��8�LָʩָȢ�8]م84\�8l�8K�ָf��8gR�8��Ҹ'��8�H�8�m��f}�80������8��8�7�����*�׸�v�8!�8ю8��ո��8�8�jָ/.׸/&�� އ8)i�8DFո��ָ�ָ��8�8�1�8�6�8F���P�ϸ�8C��8�N�8�\ָ/�ո*)�82�ָ�Ň8z�����8��8��8�.�8�2ָh1�8���8�F��>G��tІ8���8��ָc�ϸ���8�M���e�8�9�8D�׸8:�8�>�8�'�8�'�����8`ָ̚�8���83��8��83��8:�ָ��84�8]��Kׇ8(�ϸ��8�hҸ�x������i&�8�׸���8�H���=Ѹc�8��������<�ո���8����X�8ICָ ���Q�ԸJSԸV����(ոk{ָǸ+Kָ�Ά8���De�8x�׸�Tи|χ��7�8�ոV�ո���83�81�ָ^��8"Ը���8��8)��8S�ָ\8ָ��ո������8��ָ8��8hNʸ$��8껆�s����ָ�%�8��8[�ָ�ָ���8���8��Ӹ8��8�卸 E�89@�8ȿ�8���8��8TW�8i����8ì�8�ƌ��*��
�Ӹ~������8-Ї8���8z��8́������+b׸�t�8��8$(�8:�8/0ָ��8׸��%x�8�u׸ֈ��.����J�8RV�85�ָxc�8όָ���8���85�ո���y^�8F׸��ո�׸T�ո�2�8�E�8l6��֠ոܝ�8��8��׸����$�8G��|>����ָ��ָ�*�8��ԸU�8;����҆�<!�8���8��Ѹ㥆���ո(��8�׸6�8�oԸ
܆8݅8�)ָ��8Q���L�8~f������.��8�|�8�ָa�8n�׸$��8N熸��8_%�8J���ד�8��ָ��8�����Ҹ|�8G���/�8�P��Dp�8�C�����8U!�8���8�G����<{͸�����"�~=8D��7�.�0k���.�(�a7�97����X�b���=8����)�7��6O�7 Æ7 �6$.8HH��S1%8�!8�º6Pj�7�l�����,��7ޛ���J�������7�BT8��7߽�~�z�6��T;�78M�7�:��&���Ga�� �8j���)o8�=���7X8%#���w!�؄S7b���7V#�8��95�ܓ��O8��;7��Q�I0���48����膸�jF8�k�8@{�6�ty7�����8T�V���5
����X7�15��&� ��7p蓸���5��7�@��֣8BE�8<J#8^���v(��Eq8 &�7�;����p�0��6�N����8N�8 �)�N�緰�=��\8��8�z7�H��K�8�)����7{��8��8e!�8�Ǎ������^�8�� I�7�{�8z���Љ�XO�%��6󕸱�8T�7�o8�}�8Z�{���`7<��7�^�����8b�89Lg�\�=8����8��8��a8���7�v8 �7}.8B�7�8봙���58p�'���8P}:8p�79�X�l	V8J��80"#�L38\�+��A7|�7d�8Nj+�ޜ8���7շp����U��k�7.�7@�8�&�8�+7tԷ���8�Wj8�Ŧ���7 T�6���
���P�˷l���<��������.8h���������7h��@��W� 6;4hI�8_'k����|ȷ҃8| ����k��%�� ��������!�h�7�4�6	�8`�F�n������|U�����<_�7�l�8��
�y�����Z5��ظYL�8'7�81���8$|G�|�Ʒ�r�7(���K8�Ɋ�ˆ7���7�`�8��w8�+\���O���27����{��
�e�-8�%�� }:�D�&��8���8>�L�0�X7�"ն�x�6Ȭ�7�7�8 Y�5�w��m����!/��I8���0^�7`'D���7���6���L�l��ȫ�nuR����8H_�6��0S:���8h������7���p�6 �̴Ό�88e8����u���y<8�"A8६6a�8Xu8�1����O���(�Պk��[�7��T8�)}8"n_�z��70$�'��8p]R7�ߢ7hQ���8�lf�b��8dk?7|R�7ĩ��~��l�J7o�W8.�B���]���#8(�8��!8�O8�08#{8Ї�6>�(8&�ڸx�73��8K�E8�h$6b`8]�7"��}���B5��1���_8��8`80�Z���7��7v��x�q� �6q��F94�L�7M/�Ħ0�BO�7 � 7;�����Ѷh��7�G����#���������C��o���D�R=+8rG��.h�7d��8�
7Py7^�q�x�i7�.�8�Է�I��� 8�K�����7�$���8�J�{y���y8*��(D{7�����'����W7���8 �������	�&+7�08��h��ݬ8K&8r��j喷����8�Lx8�go8x
��L8�6P7P��6�7@�L8xJ�7*���F�#������r#8�����=#��1�`1���08>��s-y�w��8�,�7���\��������^��s� ���8�7ݷ�^l�yu�8(죸22�7������g89�ַ
,>�Z��8�78���8^����'���8䠷�876���38����nٶ�Ed�6S�8�靸"?���k�8a¨8>����7F���F*�7&�z8r,Ʒ���7V-����7.gϷ0�72��8�{��v�����~� ��6����	�j8�P�8�Β����|g7��x�$�8}8�8�A�8Wm��U�8�N|�%���X.�7�̍��鬸)8�"8D(�8�{d7ı��=���x���,�:���ڷ����X#з��_��w�7[�y8Н���X��Ch�8�$	8���7D�8��7�^�����7<���ʜ�7��L8 P�()]7�u�80��8�+���0���0�4�-�Rs�7��7�O�7��˷��38��f��U.8@�U7�<�7�g�8̷�N�@~e��BX7���8���8�q�7�4.8nc.8r�2���Bз�,f�V0�P��7��Q�O.8f��7~��7�rY7��ɷ�x�7�=c7`lk7�|���8�8@;z��d72s׷^5���5��:��8��`7(Sk��d7��K���X�u���H�\7�Y88��7>��7�5�����7 �4�fǷ��8��-���O�(�U�z�÷�(�7��̷�C�7�Ƿ��7���7(Qa���0�� 28HYL7a����k���m���ķ��䶞��8A�8��1�[-8<��7���7T\�7R�ɷpY�7hWS�v��7`wηH�V7@��7��V7�wU��P8�A�8@�d��-�8rη������8���7���7�P[7�W�Tj7�K�7��7�f��~C�7jt�����:�6�[�8����(a�70�^��{�8�Z28`#[��ɷ`��7p%c��'� [�6r��7���8d��7X,%8BE�7\�˷�Y����c����7��8bĥ��A�8���e��eʷ�(�7���7��Ƿb`Ʒ�`��p�7�\7XIͷh-8&ۤ���ʷ� X7�i,8�V-�(y(�h�M7�0���-6 Ʒ�����7dNȷ(��89J����ɷ�Lj8@�\7X�ķ��ܷyA�8�*�7�Ƿ���7�Ȥ8���8x6Q�~�#8��S7�j7ބ��/�6�ҷ�ْ7`$ķ,�7�ŷ��7��$�0�X7X�]7��38�%˷�.̷`��73<�8D��7�R��zg˷��R7���7 "T�f��7��b�K4�
��7�.�5�*0�
V�7$�׷/B��D��7RF7E�뷈ya7-�6�ї8:��7��.�\7��߷aĤ���H��{�7�·��ɷt�Ƿ�J7��ȷ 	^7��x6+Ӧ8�/�8ȗf�Z�18��˷�eҷ4��8��Ƿ���7�RH��wU7�18P�L7F��8^z�7F��8<�·���0��7x�\�d��8��^7��Y7���8�ե��c�7��e7��>7C����P7ʩķP$�7(�7��f�H�W��a1�(�Y7*x�7(n[�@`�8҄�8؃b�8DL7�7����~K7<·��Y��XǷ �U7��)�Aiq8����Ŷ���8��J7�᥸8�M�/�h���q8|<ηN!$8ЦU7�T�*�÷`�-� �T7h~W�,�÷\�ƷXa�7�A:7���7r��7���7(�`7P�ķ��d��e-8~+���7�e���7g��8�Ƿ��·�`���������7��7��a��j8`#��!����W7��7�+8X�T7�28T�0��08��Y7��8������Ƿ���6���7u�,���ݷ^l�����7�\�7:�5��K7�Ҧ8m18�|Z7KQ28��ɷ
�7�Y���Aq7��_� Y������5�7$<��@�7���7<�ķ�(����˷�T7���7*ʷ��`��/�7�X÷���7d�ķ.��7ED�8��7�÷>9�7غ\7��Y78�A7PзJ�.8P�h����7���7� ���:�7����Ds�7���8VF�pmT�h��7@�R7*Q�7�n�� ķh�Ƿ6i�7
w�7P,l7F�̷"X���Q�7(Y7�,8��F7�r�7�%�� ��7�tS7jB8���7G�8M/��~��F��8��1�@K̷����l�7H˷S���ķH~_78����ڤ8x�V��g58�C�xW7"��7J.��.�8�ҷ�h���E�'|�8��N7.|�7��7
¡�HBd7��08WS��)�8�%S�(�\��xQ�T�Ϸ:"�r̷�ķ�W_�JS�7V�ȷq�H+_7^ˣ8d���o��J,8�e�74D38�2�7$4Ƿ�C�����8�:Q7��7�}8��*8����XG�7�ƷRϤ8��8����CN��gǷ�We�=�x��Bŷ�÷f;�7�ʷ�ʹ��$ͷ።8b��`�8�kƷ,���	S��Ʒ@m6�\緔=�7 �t4��7��� ��D08��18��8x9�����v8�>�8�ո\�!8�f�8�����^,6_���2��8�*�P����ȅ8 B0�ɀ�8 �6�+�����8�$��# 8�"8��7���}|˸ =;��˸8*�80� ���7V�8"�r8h���8�g 8 /6v��.@��5˜�, 9,P�����7���TT���偸*��8�J[6ܞ�8G��8��A���7U&3�x/���Ŵ8P�8a傸�i��,EӸS$|��4������@�c7�3ϸ�X�6Xtϸ@QN��͊8(�8<��7�z�� �c6H"������<O���b�8�h�+�����8��8�ˆ�����\�9�y9�����
8��9`(ն���D��7d���=��������8<�������,��74N�8nAʸv��������*�7`��ɑ�8�7:K}8ą�8ȵ����6�Q����7���z��8P��78��:�9�3޸`�5�Pخ�G�ո�\I��e66��E�$#�8$�7s=ӸG�1��ڊ8��8�ָ8�r6 11�6�%8��� x%6��,8�?�8�ָă��&�28@���P9�6v)8��淀�7\s�8��>;���O9�O9p}�8�����������6gI��� � N6�٤��ޤ8eE���Y-�;(8Q����C�5$9|����C�6�����l�i��8v���Я6�Ox�7.)��F�8Yڡ8ؤ �J�8I���Н7�b8��7GvҸ�_)�B8,�r�8�w�5,9�;%�@��� ���x�8�? ����8��8�I&�t}�x-��l�8 ��7��.8D&9��� w`�U+�8ǂ�������k�7|(%�,z�8r[m�V@�8 �"��=&����7|�7-��`?J6E������$�� 406xA���1�8��8��&8�}ո�h����8(����8�M7U��-Π���� �6!��8�8� PO� N6J4����8���{�'��V!8P��ŏ��C�7Ư��,��8�Q_�u1�8T�踀�6��7+�)80����ɂ�L"�ʪ��h"�7��8PF�7�� ����8��&�仠8��,8��)8��8`Z6Myָ���1��x81)�����v284�8��/���#���0����8؛�7�8!c��@&Ը�$�/A��G�ָ`��6�K947�7>?���!�� {��H�׸��X����b�$��7*6��7�U�8�O9�>������^8���8�÷8A*8�˯� ��7J�T��0R�z\&�Ԍ�7$4��`e8� 6x׸��V�l�18@n����7\�8��"8��#�(��7�c�8`�M6��7lL�8��8�38��8�͸�pU�@�5bM,8��7��8�J�;���s��$�8������8���7�W�8`=�8,�ָXU7�" �������8ך�����6�_����8C$*8J��8��7�d�8��8��t5Pv%��뷰r�7?��-&��D$���
�l��8�	)�H��J�����&�@��2��8#f089�8{Ƅ� Ӹ�p�П!8���8\��V��8jq%8��U6���6 gi��{�8�ф7�8��/ۂ���߷�Ӏ86�8�B��'$�8��8 [�7���8+�;85LԸs=�8R9���8��ﵘ��r��Fт�@K��o�7�۸����4�@�5�#�7t��7[�%8�PI8nR����)���T6@T��Ł�@SR6�m���U�8��%��n���N�7������B�8l�8?a�8�������N� 8�I��`ո@��5e9��P���O҇8 �h�v� 8���8��ٸ��"����kC�8��c(�%��8�Ӡ5�ƹ8��6�a�����@���u58V_��O���)9���8�o�8�9�6@H16���8�,͸�ԙ7݇�8����ո����6�0��t�8�ւ84ָh)�7�q��f���7E�7�e�8|.V4���+�跺R�8�M�7�7�sp8L��70��7[/�8��7��7&��7��8c��^���S#᷽+�7���8��귡s��^����~|8K��8�g�8���7�D��D��8)6�7ٸ��%|���5߷.ɭ��,��.竸�B�`{緤��8�852�����F۫�Ľ���&鷃����P�������7k�4)�8}��n.귤;�7p��7��7���8Y�����8�z�8f��8l�7�Q�7�����/�8t����総6������8i��7�U�8���7��7悭�B������7���8����.89h���ά8���8ZW�j��]:�8�$�����7���|
��%��N޷?���� ��8>��Y���K�7�R���\��m��8���t�I8�(�8�H$�8$���䷘��B��]o8.��8\��76�鷁$�8ì8�H��t�8;\�8t�s8_���	��.���+�r?�m��7�_緄����8��C�7�!�����7o��7���7ny�6�΢��Z�8���v���i��%*�8��8V�շ�y�7�H�8)P�7A~��/X�8숮8�淯��7��7:w�G���o�O��8i�8��8B��D���i��7ݹ�����7=�;8��8������귀o�7Y����2�7����y���	��8��7P�7�)鷨I�7�s�8A��0��7��8⬚8���8���7pϬ��z締�8!��7����U��7��7��r8��g�7_K�}������`D�����J��tX�8$��87����8h-�7������쬸5#����7���7d3�7�^�8~᮸� �7��8 �8��80f��#���޷8!�8y�������ޮ8 ��Sӭ���7�o�8��7ý�8�䮸��S�8�p�7�ͪ85�8����<�8��.x�8ǐ8�~�78J5y��������8s��7�n��j���yo��$��8����7MU�7�٫8�k��yP�����7�r �hp�8��7��7���8J���2�D�����q�7T>�:F�7z�6��8� ����7Yo����r/�L���%�7�������8*����8�:����7��p8ن�8�S�r��WI�8�ܬ8�O��o��f����l�d��8�E����7�M�7��ﷆ1{7> �����N}�8�Sط�H�8E�7����Sի�)�8\�����j��7�/�1��8�l�7�b���)�:ߝ��p��������s�7�8�[���D񷗧�#/��[��s�귯��8c$ѷu�8���7���7��6/��ѳ�7^�8���C�8t-�7�P�8���8Rw�I���[��J����_-�g"8;�7��7�d�8_��7���8�I��[�8�38��7I�������r�7i��7.�����F��7U��S��7��8ф��N��<��֟8Q��7\W�7듯8ʫ������¬�D뷳J�8|�8���7���7����`�8����SB�8j��8	��iA��G��7�&�7hɫ8������ݷ�X
�4]���z귕\8`�󷖮�7���8�y�WW�78��7�ެ8�8��8���*��7�I�7Ϭ���뷠�߷���8�m�7S[�8�B��8>�7��8�x�7�u�7 5�7�㩸��7_�緢��7ѧ��*﷌���|f������7��X��������̪���7qY�7w��7�0�8��8h�G��7����"���R�7<�0C�8Z��7Z&��}w�8�췣H�8̅�	����7B�߷Փ�7M��7���Nڨ�r�7���G�88_�7���7���7�譸���7�Q�7�
���٫8&�8]�����7�
�8�R�8M~�8�g��
<�8�P��8i�ܷ���8���'�p����H8K#��]��8���8n��8�
ȸ��?�,ˇ����8#a��=�7�˿7q-�8Q9�2�8���/��7�g븿8����m8ј䷲]��̏7���3e�\�ϸ_m�8�7w��V'O8�}�6�XP� ��\58h��7�jK7�ķHU�8pk7d�9��	��lM?��)#7��A8��$��o�7I6�8���8?��y�8(�ŷZ��8Q��8Kf9���8�0��Y;D�ը��>��6���6��8bs�8�" 8��Z7�6�����R��8C��8�9����̆��8��8F%28��8�k7Dצ�+���$�,�&�9j�:��$�� ���L��+9 yb�@ݷ�8�\���P��6��8�u���c�(�Z8cC�7d��8 {13�X���������YN��-�7b�8/Qθ�*���`8��8z��r|8���ϟ踐���u��8�H⸀�����6ׅ8����=8�X8�p�7#�L289�۷��.����p]�������Z8ˈ�8 =�7���
�
��ٕ���^���`2���I������8�c�5�g��l���KM8�{����83\���[��J��8����+>ָ@E�~g��Dy�����7�S����۸J���|�7t��6�Q縠k���A��
��8/x��.�8�Φ8x��~̸��28�M��,�8�9��8�gq7
�Ǹ�r48�쫸!�8�Iӷy��8᱌8E8�{﷚�N6�D���Tu�(��8����me�8���8, �b�8�	�88]8B9p78n��6��5s�ݷƮp79�8^9��8�U!7��9 د�� 
�{�U���g���8��߸$m3��F��Ƕ7�÷�l9&8w7������0s8�vǷyW7@�8V��8��	9��&��J�8<8�8��9��98{��n��8�@��t~���F<�vH߸�.<8������8��&8�%��0n8ؽ��X�8i��8rL��@�����9R&�6�38��V��챸���7t8�n�78c88������u��8��98��$^8�R�@��7$K�mB��<����ɸ�Go���9p;X8_:�8�۠�l�����;���;8{H��U67߽�e�8<BP6�9�ĸub�8�6n�
m���t���P8m�ҷ�.�7/�9����/E���9Gj�8P8���7��N��ء���57-������]�j8�`����8ׇ�B�d�.���N8���<�N��������O��{#�jjS8Ƈ 9���8|\�8�̌�����$�2�ʶ�38rظ��38��s���8X?�8@�b7����K�{7����8��m���8(��7�x�8S��8�)븒������80`�7�u׸蔋������8�'ݸH�8���7{�6���8��� k��ָ6������E��wԷ���8��8P����7X;�8�r�8�t�Y�縪=�s08u(��$)��QJ8؟9c�97�ڼ�9��n<�
���uK�8P�>810�8P�3��l�7������8+��8��7����8�!v�  1���0����7���8Aܽ8��M8%��6�K����8��d8ԑ�����7
�8e�η���:۷	�9﨣�zL��4K��y������ ��8�m7�����?���8j8�A����8�%88s���@�8*��7d�9��6�J�8�$�L�9��6�>��g�j���I����RB8��L7Ŀ4��ԍ�9(8��Ӹ(�92�{�Y����X�8g*��x<9B��|��\�9�$�S8�:{6�N�7^���h��7H�9�98��f�TK8���be�7�/�8��5��O��4`��<���B��8�	98�M�����82��ܟv�p�Ը�������ے�8���V(7�n�7dv9@���0>7� ���z����8�4�����иT9���NE�k��6� ��z:(�\���ɝ8���5	�g���u8��w8��7򁊷�t�3����p�����6o7&d58�%���ț7j@a����7b<�.K�7��r��}q8�
�7�(��v���҂�78Mt��u�[+f8EGs8p�7�o���7�M[8L�;��"\��I��![�7%^o8D\�7��k8FBp8(�Z�]�d���l8�'m8�n8O�n�,x8)2k���s8~�q8�L���n$8Lה��䒷��t� �v�%�l��0t8��p��o� i���!r8���7��8T�n��r8��v�h^n��r8Y98��`�);�7m�]�,2y8�
o�m&��yП79<m���5M���|!v8���æ����v�l�v��A��V�7L�^8.�A�N@o8R͓�.R�אu8l�q�.�7�ȳ���j�z����\�������a������7��x�m�Y��᠞��q�īw�[u�����#��������{�K��7q�78�p��p8M�u7;�M�u�o�p��7[Fu����a�o��7@�d�Tݓ7�]r����7G��>�77zo��J�7F8޷D�7~Ō7�ju8��7s9 8.�e�m׈�
�7.��77�Zѷ��o8̜v��3q�K�t8�%6ffm�	�a7�Y7c�5�JE�D��7��o8E�����7#\s���d89pm�%�h8O���-e8l�q8��q7��n8�%�7�
��R��7Qw8��r8F�w8�ۙ7�O7Z�o�>	R8�#m��H��*=p�'��7�dr8	�e���ҷ.��bw���B8�^��e�q8i�t�K��gjs��g8�on�xdp8���7��n8&�i84�n���6�]v��%k�Xt8�Q�7�o���k�V�_�]Fw��n8��q8po8U*�3�7l�K8��7v t87b
8j�w8_��ܜ�7.`s��q8��Ts�n�{q8��s8��7_�r8��7�+8:yh���s8�ʈ�H�m�r'o8�r�"ql8���7��.8�=�7�d�]��7y�u84�Ϊ�7,R�7���s��;n�q�T7 ���MO�7�㙷���l�}N��{bu8�o8o����Γ��"r��Hc�7#m8�r8q<q�x�v8��n�'Gj8k��6F��7�ͷ/�7dzn�`������7�o8���7LM?7 c�7�+�7�z��Xn8�,p8rLl8���N����Wp��vs8<d�7����V�w��7̣�7�S8�h8�u8�ѕ��l��P�T���o8݀��d�7���r8�?o8&8x�Cq8<꛷ɤs��%l�.�o� �h8s�p8��p��֤7��o8h�7�n�>y8�u8�i���#���l8�����!y�҈�7g�+8��7W&���P��Lt��;q���^8_$��𸋷�t�7`L��k��7��g80���>����q�J����n8�2u8�����p��`����s8��m8�-�78u8hb8V{w8�1{��ˊ���Z��!�7 �r�-��7����tg��.n� ����7LՎ7�,�7|'r8��l8�	�7MÍ7}��l�l8�/�����7�]p��Ӝ��t��+�7Jq��r8��t�ADi8%�p8��l���o�lo�l�t�{��7f
m8���7~⓷L"���g*j8RWt�B�l�b�r��J{83 ����h8�-w���q�@އ7X*����x8v�o���C8 ��7�'y8����$,w6��k�G���`�3�38T s�Bm8 	x�7ur8"�H�B[t8GB���@p8���mʕ�lr��l��7m8*���Ep���7xcr��9��C��>ѐ�>�s83����"t��e�����7߄l�n�p�^����~r8O�r��+�7u�7���7�ƌ7��>7�_����s8��m8�u8)0���p�7���74�>�c�j84�\8�Ր7bU7�v���\n�r�7��l�9�r8Qv��r��C������ƌ7�Lr�ב08�r��"�t8-�v�����*q8�QU�7.�7��n�b��7��s8sGw8��p��!s8.q8�	���ʍ��7`�o��@�7�R���(t��uu8;xU�	�8��8Wc�8� 8���8�z���l�8�6��B�8aK8QN��$����8Bk�8$�8�i�8��v8/+��^�8@l�7�9��ZJ[6���8�B�8�ϒ��S��<���+��8���8�U��\�j8�U	�ށ��o���M���U
�MI8�������87Й�yX���Z���h�8����� ��x8����m���x8� 8�d�7?O�8���8<��8B?�7E�8�f����7���TO�8Ǔ��fz8���7��8b�4M!��9 <8}�8B��8���b��%��8�^8.� �������18T������7H���t6�8@�8�d
8��D2��Cf8�����=8���8yB8���8q
�����	8hВ�`G8 !��#�8߮	8�����c�������?`80��8u-�8^i�8X4�8�������7�m�8a�����	�c��89虸������8���8ȵ�c����Z���	�2�8D^�8y>��)� ����82+�����������080�8C=	��u�8H�7wՓ8fِ7#�8��8^��I�8�������M����ޘ8&o8[#��n{����84��8~k8�c��0�8���f�7'O6���8I�8	��ő����pI���6������9�80闸�������z���<��c����ᐸ�6�b��Nt�8+��7��5���7��
���(;��w1��ㇸ��7K3��n89싸�F8�;�8�.���ژ8���J�8Ʋ8�,���|�����8�S8���x���e��d}
�(� ��@�,��8���8י�(���{
8�28Ź�8Y�7�����gY�7雓�oC��}��8�	[8a��7�v81w�8��8��8�ۙ�(��:�����:bK8�T�8ꌊ�>8`:�8�j�7CK��1���
�z.F8���8D�8T�8]���!�0	��T����?���Џ8U.���8�	�'W
8��7E�8�����!��@$����7�9�����8j��8��F���l�8�?��
&�8�m8w��8�^���>��J�8Қ8(��˺�8�ך��K�8[�*��ٔ8!f
�\F��l���6�8��8�ܮ�읙�)��8����8|���q'���p/�T?�$�8��8����rl��$���	?Է��8z��P�
�V������?���I�8�X��P8� �T�8:�����!��7)��	��8���T8㓸vǒ�����ϊ8GS�7V#8���8��8�B8��8)��7*}�6Gf�x��8�}���� 8���������
8��q8�P��q��7�D8����U�7�.����8|J8�g�8@�8Ӓ�d)���9	�pV 8�-8N��җ8�ȑ�9&���Ó8���o���a8�X�8�#�813�7"� �G���7ܸ�7K� 8h�8:��Wˍ���	8��7��
�L��u�7����6 ��b�8d/�����8dԛ�lU���8
��8{��8(a��-��p������c8u�Y�8�h�������8&���H���Ә��(��_�8��8�	�X
8�n��b���18 |�5G���t�8��8/���r;
8k��7�������Y��P�08�f�7b=�8�u�7q�����8&c��pƒ�Zx8t3,8����A8 g�<ד8�	� ���u����7mᑸzÙ��o�ɍ����8IA�8�o�8�8��8g����83ʑ8	S�8Q�l� ��8�������_�#�g�����84�p]�8�
p8x���
8��s/��j8`��8o���
�����s��\���8�:8h2��A��:'>8���7o5���,�c����	8
� �o�8?Y���[��ݚ��6�������8U���7����8JY�Uc�.9���0���	��1����88 Y����l�@����F8#�8�M�8l����쑸Tp�@EڵP[���n�x�˸W7�8n�����5��8hh��f�8 �88�D��� �0{h7fJ�8�Ґ���6��68�L��γu8���7��8ᵸ�FO8�Z �}�8�����*8t�5�RW8�+6 A�5��8/�и n8�Ʒ�֏������8��o�|�$����,���g7��Js��^7ND�����7�+8��̵�`28 �`�xo�����q�1�8���8�����@Ԇ�x�U��8P������@a8`:� 9W� n�5�@W7�$7hVոE�����8�*�8v��7Tsl���8�R)���6�N�5rY�8�2x��658t
�8�0�柸�zI�� v�6h<�8��r8���8Տ8�B�8ڠѸ���5NRk8h�[�ԡ9�<��7 α��OY8���8A������8����׊(8�"]7Q�ɸv��`�8���l^�4:�D�e7 u>�;�8��`7�*�8�9�8ȼ�7��i��(�'*��6�p8�=^7��r��o�rY���8��7��8�y���ͷ8����I�8�Cϸ �8'����87�8�p�o�̡�8�v7�θ\P�8�~�8���4���8�t�84��7�68����.
w8�Vb� ;���M:�p��8ڴ�B��,��7�w�8 �� ��5��h�@_��@e��7 ��50���W��8�W��֣t8��������Lw���>8�F78=�8@U�5�M=��f˸�o�s}̸��s8 f���mθ����l�XS���W���.&�̊�8���I����öR���t� ��g��8�8�L�7�"58&����]98�jt8�Qt8�p��ep8�i����Ѹ*ˑ8hq�7"��8���XNq8�µ �ɵ@|õ@�Ѹ�������H���$�ʸ<��8�߶�*.8�Q7a"�8�6m8h��� ܔ3"����C����8EW8�@�k8�N���o���8��m8?����8|8ϸR�8k�s8�m��6U�� �8�:��$U���8����"��/`o8g�L���8)���l��8���84t7Tޔ8�~m8�fo�l�j�����J�5��8��
6F�����6$�89�-8�9�zI�B�6��D�8��0���8pwQ7@"�5��0�N�8�� �
,l���l��8B� �> ���{7V�88�t8(�88yU���E�8Ft8"'���Yr8(6����5���8[��85p�>�и@�5t��� ��8f=�8�Ҹ����鶸���+y����5:�n8�Cv8�T�N��79z�8����lw7�u�������(8��8F�p�A(��'48�8�ٷ�F�����wa��t(68@�6�X��HNs�u��8L��8 9V5���ض 8Q��� ���8bs�  �̸\�%øCxǷأ8��8@r������t8�E�8F2t��L	��1�5��8�#88��08 #s6
�7p��ٕ�p���v��8,�x8���8�5�8�_9�8^��5��8<�7�Sٷ4��8An(�����/�+�������8��8,��8pOɶn+1���ѸX`Ҹ��o88�(��-|�� n7��Y� w�ܯ�7���8Ep8p4����7�8GY�8K18�������ɫ8�h{6�Y5��и�aU7����8i����5([���H�6�q�j'*8�33�v� ��o�2#�����8,�m7j�8[�6�7�8���(ep���8d5�8��n7pȴ8�浸Jy��껩8䦣�@��8���~��7����Y4��xe~���y�>p�T�a�S2�8 Y7�����M8U8 �`��6k@�� ����/�׆�8WH88T<p�����J���j4��	-�Jr�T�8��8&6w8��6Է8$�����8�]Ӹg���t�y�I���U7b�8�
6������;�i8��m8,��7�l8:�8��6R3�8@��5�ZV�4�����6�؂��0�60��w�6��7j� �n�`8�l��}�`7��7�7�B�S)����ҷ;ׂ8Xζ\܃8}ǝ���8\�ַ�뒶	5�8��]��!8
Hɷƭ��@%�8����8D7��^�-l�7%⋷ų$�6)�6.���p�7z�8�+��Ƴ�#�88��7�!����5��I �7iqD���ַK�߷��C�����Hi���i��3}ʷT�5��6�Ir���G�P�7e�8���7��6e�6�18��5�c���q7{����RL�'��7��B8��_�j�ѷX�7&�׷�A�7(58�ذ8�bV5�7�#�����8���7�������vd���^8��78͞��jҷ$1�78�79�˷����Е7�A��%�]q��FMB�;���NSJ�W��72!ط�+�7�8߭��'�8�ט7_�����D���7���7��8nT_��v71�N8|��7C�8�mϷ��u6Rh�7��ѷ�ڷ��8Q���·9F8�6�5�����HD�8��8�	8��8�ZF�9����@8�E�$ڷూ�����-�7�#8.܏�ى�7��6!�&6WG������1��8�S���ϓ� ���^�;7���7�|�7����Ϸf *�
5�7��g8iKG�ɬ�0�8��^1��L:���n�L��A9_���7-M�8�o-8Q�7��<8n�$:�����T֝8��8o�_��蛸��7��7z����·$r�7�]�������.t���^��J�7/�8ȹX7�ꙸR3����6�n���+����8R�[�^G0���?8v��7$-*�ʊR�u0���-���d�����<8��7�6F8b�7j)\7����r��8�ڑ�-�ڷw�)�'��e��7v,�7K[�7;�0�e8�o�7�J*7I�#8a���T�j���7~��/�J���7��8`q�7=�E8������7��8k�6��6k�T�H�:~�8	�7T8�'�8�m8ZP�8�>Ƿ��8��ڷ>��75��E��^�{�E7%dH��h�7����{��\:8���7'\h8��r8L�7�R.��H�8���7`I �J�.��M�8:-�7��`7tGD��D���~����8c������7W�x�`7A/6:~��7e��6�f�5��$)3̑�7�%��u����1�����7*�h��ӷ���϶�1-8ƀv�*;�8&�r7��ڷ+�7�B8�] 8}3�7z�8FA�7h�d����7	��7�bJ���8y��7+�c�Q�98Eط*��y�8��8�
A�cg8��
��s�8��ʵ3�<z+8-S8����s;�����W����v����7m�8
�_7�ȷ����7T��7xM6�;8K�7��F8��j7g~)�oE�m�綈��8�8�5jĤ���#8C.k���C�Cķw����=��=�8����yI�:j�6D�ʷ���7��h84���ie8�	s�Xǰ7�d�8�j8Vk������y�8F��7m5�8kg����S��ꚸ}8Uۜ��X�7!�ѷ��}7������7����RH��qU�����7T�e������Z<����8ӭ��>����I·��U���Z��*�7V�7�؃�}�c8�F�8��~�2�^��eI��a��i�y7N��7>��7��8å��3�c8��}�v.$8��7�vb73���� ��u�	�5�t���;8������7������%���8\�U�iꊷ�8Y���9c6i��7�l�<J7}���88gn[8X��7w��5�^���H�7�����o�8�e80�ַi:�7��8<���+5�/�����]���18������4�d"�4C�8%�7�v46
�ҷD��8��8��ַ1���ͷ�|8W�!8jL��K��yַ3�6p럶ȣ��7�8�y��R��6A��7��Ƿ�w��ڜ}6��Էϡ8�嬵r�Ƿ�h���Z����7¥c��1�6�ɷ�2&���'��k2e}g�O���q=��*!17%�14T"����1֔��&���`�C�<2�A�.>���8>�/��$2w�41�-�0.�y1ˣ�+8�����1�l1�"U26)�a��F=2́�7���1�02��22:�<2��-2�m2񪇰ч�0��1B��1�Pi�?�1ߙ�1̌2����'1�^�1��'��2�1��;�p�n�f�c�t�u�퉸�i9�1�=�1 ��/	Yv�AR�0��2ayI�$�M1�0m�D@ �21�1<"�1CN	�����6�k��0jޗ1W�2��*���̱���1�~�V$��q�Z2�Sձ�Vh1�3��:�\;�1�H�J��1�)81���T��1�];2�U�1��I���ܱ��0��]1��401�1�,1h
B1��#1Z{F2v:�k���&-�5�Q�B�32,R(�5��1�7��|��d �<rB1�|
1�? 1P�2�R2eX1��ذ��2��k�#�!1�T�1PjC2ڣ��q� 1��H1�H�`�1q2�1�X6���Ѱ�9����0�R�14ӱCԱ�\�I�1/����2�(17��0�n���1�g�!����s�1N	�2��0�:!0��˱�\�1��02���z}H�D�����1o�2.K�1���. %1���@�1[*12��1�V1
[�1�52��0�ؚ10����'�r
ϰ�A"2�0A�d]��$#2ԩa1t���˱�;1<��� �*�1�ı+����!�T����{����2d'�s��xO�1�쎰����e�1��2���gұ�Fѱ"���×����1��1.���0-Ǳ����}o�:$ѱ48���<�j۱7�N2��1���}��PG���f1�|��f2� ޱ� �� �0��*z2Z[� �N�|7űs�2t"�������2Vy2�1ӯɱ82�v���we�?�1�8[�9���1G2������1Og�,����[ϱ�����M�	QݰL��	�Z�A17�0�{�1���1(�;�ұı&Ţ0��ұ"F�1�귱�*ʯI֌0��J���Q:�1���ۖ1Y� � x0LO71��б�{�1��0�C2m�:1BE���H�1��b�w�2x���:������'�1d*\�����T��1���>��1���:&1k	�.g1#�g�=M��~��1�pK1c��1��1d'2]��1BE�� �1V4�1�9��7J2���������̱S������K�s��1�v#����.|�0�2��������>�}��Vl1߫�1�t���1	����*1æ'2)�񉱴v豘�����2��1�/����1݉C�2<��f_�HJ/1��۰���k;2/���s�s��ۋ���İ"��1{>����I0	ܖ�&�p�&�����<�2��0�1^�+��S������2����ة�^Da�A2(2"�V1	���&ۙ1�1+2�x֮���1?]�0�ӯ���	2�2>��0a�	2�2����F2��1�I��y�U2ž2�X������9�0�Ű�q7��1���71���0�;���np1���Nئ�ڵﱜ�12^T��`�h1G] ���t�ذd�R����<aU1�e1���1?��1
�1%{K��}}���1X�t�_2���7�2��I1Zt��#��0����]2c�����F����5T�0��1��\��닱	۱2A���P�1����ֶ1ȓ2��ᱪ̱��6�h���1@�?1��2s�#��A11nxޱ��1=�(���1��1O/`0�T2j�C���/�Y�[W�1s�1�H�1�������X���� ��1���1�t�1&��1V��V��/�L2y�°M=!��yұ[�11x�1	"E�`�1��2��s�K4�.���U��yŶ���"��4��V�	�t[�1ƙ��kB�1n�}���ɱ��5߿�����5��˵�c���;��T�5k�̵�&��]�е֑е��5��5�5%��51�����5�ݶ�ao��?/5���5�׵$Ծ��xе0 ����5ġ�56��5�d�5򷱵ޠ�X���^�5J��5`.�5�ۭ���5���5�{�5]j�5��l������5���5�*ɵN�5r�õyR�5�������Ut�5����監����nz��5S�����]㤵4�������5�������M̥5<���@��M�5���5nFյb!˵�7%�&��'�5�y����|�`��58��5�)�5�<�)��5����<�4�������L��Q���V�5/-�4���5>�y5>'��@�5�)���E^5I������� ��st�ڷ������ ��056"�5`�۵����*��Pș5���pР5i�ҵ�	`5���iS����s5ֱ��(�5W��5�ߵ�t�5.��5�{5��c5���5"롵j6A�3p�5�묵$���i5,�6�5�5V�52�õ1�ĵm�5V�5s��5�D�5����(�5��5��w5�%q5����g�5���=����5��5���5���޵�ŵ:kõܜɵM�66���h�5_L������^�5j36W�����5Ok62@�5��5�4R5����x��椯5���5��	�i!�5�k�5���5A��5v ������e�5˃�5Yܘ5Spε����n�5�v�5�����c��]�~��j�G�/�Gw�5p�5��ӵ�ޠ5�v�5����6^6������56��~@�5#f�5|���u��5�J��4U����Qq�5���5����{���ĵ@�b����5���5��\�\�5�5m��B����ٵ}x�5r���F�Nq�����5�r�5ƛ˵u�5�{����5�Z���wv�{�55Cϵ���������1�5���5�d�5�����6V�(ŵƈ5r�n4���5�$�)�5, ��X�5�dǵ�^�5j��59L�*s�5 յ��53>�5|B�5<���pɵL��	H�^��5پ�����5�_��QA�5F��55�5�{��*5}��5��6h>���v�58zI5�=ɵ�G6����5QΦ5R�5�?ܵf'�5U�s���5?F�5g��5v]�5��5�CB52s��l�5���}5qh�5�m�5s�C������5��:Ρ�y0ԵW�5��5o۠5=p�5�۳��.�5Mɵ��5n��5��5�(�5)T�5�`յ�o�������z�5s��5�x�5�%���&�5̋��nN�9�5���5�ŵ)Õ��╵h���~���5����CE���j�5�6�=t�5�ԭ5�o��z�_D�������k�5�K���Xص5����a�5�N���u�5���5�>�5X��5�}�5�%�5�is5y�ѵ������5�56:��!��5ǵ�孵�Bµ�^�56��5�5���=n5��5�5��5�?�4�9ȵ�#�5KIڵ�ކ3˰�5�v�5ܻ����5c�5󃹵E���ꤥ���5�۶�4t��4s�5*��5^��5�;���EĴ!��2p��`�������쎵\�5�5
!ڵ
��Gֵ�5">|�=��5�g���5{��5�@��`�ɵ2�5��5?ܵ�Lߵ��ȵ@鄵���5eSԵH|�5ۿ�l��/��5vG���$�5c�5:���Ĝ5��5��׵���55m�5D�۵L릵�D��?A�^Kg�;��5ec��.��5�4ε�~�3 ����_y�ю5�g��1ݵ@Ҟ5`�~�DV�5�����{�5���5/�����5���<��uH�5-S�5�嵽�5ka5~��5�Ј4�f%4ᲵLJ�5!L�5W��5����T��5 �5S��}�ٵ�~�5u6�ϩ5^����B�5�7�5�4W5����4��5?h�ߡ�5bu6乍5%aQ��6��W��5���5=�5�����Ƶ�W�tJN�[+�`a�51�����Ϥ���'���pAq�[����7������V(��d{�7�x�6�27�ƶ2ߧ7���(�6��8��7x�����8�̞7�m7�(�6�� ��7��ST8�47�t�6<��(.�7����R��7�Z�6f�7����_�6ڎ���8p�*����+7h]���8P.˶��8������@�7��8{��Dh!7��8P 7PN�6��$�<9/����d~���8䰜7���������7�"���7W������.��r\�7�x8� ����79����7�ͪ7��7`�����x�W��z!�$
70�60���0��d��7EB844�7:�6�r�6�੷�X׶ �7��p�S�6�K8~����u8�ت�j�8D57:��7�h�Ŷ�����2�6P�����t7�ф���5�y�7~���}�7�537`��6(�$�Hτ�����z̶H6�7��6P�׶<47x��,d�� �8�!��83�6��赼��7�s����6 �(74~����,���� w7$<��9�����D88�ݷ�.����1ʶ����x��6L�7 $47>�7𾛷0��7(i�D\�����8���0:7�)'7�5�6��϶P[���J�6���7�^I7T��(=8�D�������6�՘� <�d�7�k߶���6�<�����7�-8Do&7$	78RY�����2��l<$7���7 �Ŷ �)7F%�������57 �6;�8��7�d�60n�7���70�47p�,��톶����?F7��8iF�Ϥ��������ዷH���h����|�6����7Ρ�7�ĶH�����&7�-7Z��7P��6P���V8��T��g����$l8X�6�����������Z8�w�6��8T�
�2ǟ7T/���O7�N�7�>�=�8�����7�"8D]27�Eж�i�l(2��A�a58�M���M����d1!7ON7�C�7\A7%%8�����6��7DFI7P�8����`05�M�8�)�$!�D&7V��7$7x
�6��6H�708�0����7�����7����g����70�����8('�6@Ͷ�6��7�%ٶ�G�7(��6p&���5��m��5�h�#7
�7�6�7���h}�7���n۟��@�6����7S8��7�))��W�6l�.�XG+��`�7�t�7�8�֞7�&��yy8h�%�X��7��!7����l8�*�7�6�78��6�I7 +�6H���!�7����LǛ�����Y�E�8@�
6�v�7l%7�f�7T��7l@m��}�z��7 �����6(��6x��6h%ж>x�7��S)7p6�p�ݶ0���|x`66·��7�?57l�)�؜�6���6x�6
�7�����v����7(�77�/,7�h�6i�>V�7!���h��@ђ6��8�;�6j�8ؐ�6�>����3���7�!7�����7y��������L7����j���#�	����$׶���7`�߶4��N��7�v�6l�-7���7@�ն$�� 	�6�m���ݡ��/7��Ը!�����බ�m#�5�*W�7�17t/����7�	ö(�/7b/���7`����x��7x#׶��6➠���7@7h�k��k�hӵ�o�8TҠ� �57@�{7�r8�Φ6����
�X9�7X��6w4�7bA�7З���>6���6^W���4�60�ܶ�)7���h~�6[J�T�����7�7��%������6���Ѷݭ6����`7.���
�,%��0��d*7�2�7���F�����6�j�N�7�J/7���C(8�����8�
�6Q��Z�7��8ȣ8���7�C˶�84L�7�ܱ7p�Sʶ�����7x�6�o8�.���7����A{��(��gr�6z!��]�Z�.V̷��ͷi��8�n6�ȷ�f�7��R�K�Z6�˙����8k&��Ŀ8�ηe���8�7��17�������8�d׷�/��h���q��YΖ��/��rM�8�Ǖ8����QĖ��:���-�8�@�62>���A�8׹�8�f6�:�7��7m6�8�P����Ϸ�U���t�7��7�w̷qѷ�U��7O��bG����8��F�Z�8�C�8'�6���8�7���f�6���8a���Rk�8�t�8c޴�r��7�4�8�����8�8W���&]p6�8��8�3�7�8������6Ɍ�7t!J�b�5���8ԩ����r62��6����^Y8�Ӻ6�Z�7���8})�������~�(�ӷv䌷R��8ږ8��7��88i�8�T��Mo+�8�8N]��4�ķ\��8�`��3�8��ַ|,�8���㶓8H�������]�8�e����6�����7��QÖ�+x�8�5���k���C%��i�8�Q�����k:�8�����62�8�d��֓�8�ｸ:D8p]��]ݖ��������ٓ�@K6�|��F�O7��8W{�6��8��8����+���G�8��8�o�7��6Y`6u�6T?������R�ѷ+��8�ƷfS�8a�p�J�ķ	��8eD���"373,���^~�L{�����1��)	����z8�T��"��6�ֽ8Ԁ��V��6�ۆ8Κ����\���g�8x:�7�0{8
E�8Zߒ8�	��a��8:��8 ����q�8����{T�8 ��&��7<��7[0��/Ѽ8�q�6��w6��8���,��Q޼���6�3��;�8�N����j6�#c8|��������6� �7���7�4˷��ķ�ҷua�8�g��aý8GF�6G��8`5�8���8��8�Ҽ�t��7����w���8؟η'�08r�7��7�5ɷ�í����74���N�����8B�89Zg�B�7�Ȱ�������A<7<���퓸B��8�����B�8�ȶ8Jwx�^W�7�U˷���7��8O�7���8��6x�6շ��~A˷Dk�6��8>���lɔ87������8���6��7d��8U�8��8�qշ�$�8����A)��G^ҷ���a�7X�ʷ���7�?��e�&6ڿ78J_7"�W?�6�e����ķ�-�6�J�7�Ⱦ��Q��N��7����`ϗ��շ��8���7pO&����6����Ow�8�>�6Jз�1�7M��yi�7i[�n岸=��8k�7~�ŷ���7�������wQ�8I@�����$�Ւ�Z���b��8�8��7/�з�Q�7��4@9�8��76O�7���k��6,c��I���s"�8�ݓ�	��N�շ��8�l��>�ʷ\lJ��󂶙��К��nT��ݗ�Wd7�D�8�yз㎽8�\ȷT��7l�8�x�8�Ә�w��8E��7����j����ѷ�qw�\��7��78@����ڼ6���8JOe6W��8�i�8���7�U��R�Ʒ>��x3�8��7�a��q��8M����p��8���8�뼸���8�ɾ8#?�紖�sW�6nm�8]Xͷn���k�8�,���&��A_8�η
��8~��8?Ҿ����
g8+�n6���7�Lg6�V[�e�ҷ��Ʒ��8dc���q��e^���׿8�e��\��0m�8�f�7 0�8{�&8>��8a$�8}+ͷ�3���8W�u�8[�̷Õ8�7H+�67��6tf�7��7�6kY��eW8��8�ض8�s��e�����69�8���6���ά�7q'���a6�Ͽ�:�������n�����7�Cͷ�8j@ڶ�>��Y1�8�c�8�Ɠ�"��8�$+�a�����8�8־7���6h�÷u3G6�8�8�����	��m"�7�;��M0�8�]8ʀ6�S{6m<̷J��8LẸ|ғ��\��"��6����Ż�������Ϸ
Kp8�E��(}����7�>ʷ恊6I�޸Q��@�6��8���8�l�7�sd�*����8u��n��5)�P߸�[���<޷�gz����8��A9��ø̞e8 ���u��P494NA9�C9H�[�����Q�E����88���E�����8�;Z8'�8¤n8	!6�������јC9�z0���2a��A�9B���u�68*��@L�����`	9	�ոPl82���J�8�v8[v?�V�v��8�8��7_�9 B�I����7+ݸ,P���7��E��Z8Vρ��i8SF�8�y
8�Y��.�o� EԶ���[��h��8�Y��̭B�M쥸b��8���z�u85��8uO߸d�u��A9�eB9 ��f�B9���ݯ8�x8��8��W8t�8a�9�K���c�8T�9�l޸H��8���8�Y�T�8�b�7 =��}9 g8Y9*!49K�A9D�D9�@��X�7��޸�nA9�bO8x��8 �嶀�K7��7��߸_�9�Nf8 9C�8�9Y�9&�y���8*a�8 #b����84�c�^�@9
څ�4�x8��z��=9VB�@�l8D�q8`#9Lƥ��N�8��e8��q��_�` o���86�{�sj���9��8����e8'b�8ٛ�7<�?�>x�ô]�w�8��8��%���9��?���׸�4
� �5Gc�8š�<Z������V�t����8�&v8���7���76Q_�6��6�r߸v$����8�"���D��z���Z��V��n�=9/��� HԳ���H�з���,�左�*�@��6��7��A9kf�8���6�(ȷޖ��8
8�Ú7Y�x��3�6��A�Т\��x`8ʘv87�
9�/�7�h����t�<�4<���d�7�幸��8�F�2�7X�Y8��ַt�|����8�5�7~�?��ặ�]��t�j�6���Tݸ`�8dr�8��s8D.�7�KѸ(�]�@�����8��7�,�8��O��D޸�/�}h#939�V�Z�e8�z��#����A9��	9�	�8�B�<��7 ��6H!��y����D����88B�y*�8N���7H%�7,�8��G6�c�8Pd��x;�8�>���Z:9���70��7h�p�.�D9ˊ	��66�Ƿ^_9��7Z޸���H�L�6Y��Vt 8M&9/������f��/�8�
V8�C��Ne�p%շ��]8�|����'6���˲�8A��q	�ۦB9���*�@9G�F6��9��⸁\n8�"`�h$d���5���8u�8���8nw_8��?�ൻ�r]	���X��
9ҵB92�ƵB�9_l89�>������9"J`8N����Z	9@��64��8ܶ�7�q�@Q06���N���ߎ0�`��7`���ӝ��џ8�	9��	�ثƸ<�7(�r��Ԣ6�O�6R�:�H'D9j �8{X�����`f��(s��@�y����i>9<�y�I	�jE� r8 x�6|�[����L�9��z8����2z8. k��~�7f8!9&�8Q�q8��P�4�޸~���{騸��8b�6R�o8��o8>��8a�C��Cb��j��%��8O��7g�8���� ���8/�C(s89����{�� A�|�8'L_8��R7=<�8����NIb8�`˷�;�6��l���j�*��8�S�JY/�.k�8���7���$g��:n	���{�7U�8�&�8:����{��	5�����u�7�$<�n��a��8�|�x�X���R���8��7N��8�����P7�8lF�5��9��ͷ��A9�?9�����|A8 2_�D��7o�7`��2f�8W�9��⸐�y8�e>8?�� W8�7߸�ϸ��	9Ȑ���(@9F�8�vq8��B9
��7R,B9�����9A�X�7b�9�A�4@9 f�H��7	��h���۶�v�7Z��c�8Z<m���bc8�@�򽸾3���7��u8��`�zz8 �d�W��8��7\ٶ�hv�6�E�8�N߸�-�8i`��3�������.7ԭ� �,9P[��u�9���4੸I�8�7�z�7޷�Cf���5�Q����(6d{¸�{18�7茸��������Ʋ7�gD7�T7ڃz��3�e˔8�8��~|!9l89$.�7�6�E�7&��j�8c�9���4�;����87��=��2#G�=}�8�D���N�8��B8���fvi8P���
i�B�-8�Iw��+����R6I�8���6�}�6@䮸j����1��ܺ���v8�t38q?�8����a8Z��k��8\ �7v�a8�<}��(�8��$9f��4�����6_���jb9t���̨շP/���7�'�8p��N�j8��18��8�j��j�68`��6���8������8&�>8��7x248T��7P�*�Ǉ9B�8�8H<׷uϔ� 2G����ɍ��i�8�O�8d��T�64��7��`8�o7ё8�OV��:���E�8'L9@ES8$n�8ɯ���̓��X7��8����>9�@�85>9D�鸼"�^wh�1�����D�"w��� 8�$��t��8P5ɸ ��7���8�
-��p��`�6�m�5Ya�8��`81�˸+�E���7(�ȷ�I7|e��n:�3��/�K8� �����7,��8x�V7&.�p��7l5�7���7F�9�z�7Xٱ7�W��`Է�G��\�7���טּ�z9 ����m.8��6��3��[�8��8��8ik�8]0���9~x��?8H��8
�F8�4580�϶m��~'��~>���7b�48�j����9�@�8���7 ��7(d�8f9�l)8L688�>7��8Z��T8��J�R��A��8�b76�g��h8��<8�j��Zu8�&2� ��8�`��0��r�8�8�H�t7Z=&����@t��7�詸�!%8�%��a�8�#�5F�\�sՠ���#�<�ŷ�@�����6֘9؎47��7/��8���8����<�7��+�d\��t�뷀ͷpS<�~��8(L�7d�F��e|7���86�%Ց��b�<��7B鞸���Y����w��l���8��9}�?�^���� 91Eиj�V���̸�q>8�
��% 98ߴ8h�E�d�޷Ќ:��a~7�9p�r7i'��Q����8��9J��8%��8j[���xF��.9��9j�9�Rʸ��&9X��nƢ8�U�H�	�D[���ID8��8l��T<8��@��Ը:b�8��C���ָ씇7�C��A�7���7(�\�F�8�}��P]��|3���̹�ʰ!�v�#�� ����$Y9$�øx>.�0}����8��4��e�������1��:���;WA���B9���8)��XF��06��t�M8h~շ���7���5F�+�LŮ���!�B����=8�9]�7�'淜�9���8# r�@�)8�Z귲
 8�=Է�]f�h�P7O����l����7��9` �x_��A&� �9,_����9�h���m�X��7ٺ8�A͸W��H�8dR8�ue8&�<8�|�7�2�5)~8��8���7@,��ݗ8��9�h����9��~8%u�8N{��N8��e8��\�)ਸpw�7W��81鸪�86~7�+8%�}�#9�棸٧���~�6�s�8���6�d�8�Ҡ�|����< �J�8ɸV�8j�9@$Q�f���,x ���@7�=9cԿ�RW8	��8;�8 2�6�7q��8��959ޝ
� ��4�hJ�������>y
8Y���xb�������97�
�7 �k6��7]�8���\��7�˖6Ԯ�7�o���W�"���
S��B���7����.�88(�7���8,�!�H@e��?�8`�p���޷������8}�ʸܞ�8@p�xx�8���8??��7~�8�^¸��88�T�p��6�$�7F�9lɾ��y��Q���&��t�8�`�8�� �Y�9=�9�J�76"H8�`f8~�]7���7'e�D���e�dlG���S�?-`86�R��ga8j�X8�Hb8�'8l���a8�f�ɴ_��.���L7I�L8��L7�c�gKY�d8Fh^8�B8�Oc7�&��d���]�_^b8A=Z7�!-8Gd���A7vR7ɴ\���]�>D\8��f8M[8�hd��W�4�r���a�^��	T8�T��sN�xH7/a��Ae���P��.��C]��.�m�X7s�c�J_8WO7��`��e8�LX���a��3L7?}X7�$c�Ib��d��437�\S7�-8Ɋ[��:x���\���T7N7�d8��I���B7t�Y��/M7��D7�d8`�X7�Ώ��D?7��e8U�Y���e8�L7GV0�.K^��f(�t"]���f��5d8[�c���e���c8��7JA`���a8�a�L�b���a���S�PMc� b��;r7j�f�0]W7��Z8�
J���c8��E7��R�\sb8ȼb7'�a��rT7��f8���Rc�ޤW7�Jf7�Q_�u{�j�A7U�b�J�Y78�a���]8\a�nId8c�e8c8��ͷZM7�e8|9a7��6X"b��6�7��a���`��Q�ycb8�|]����C|b8���7nb8T�S7�e8:�L7�d�%�e�#b�IXP�8+8~7g��@_��\_8��a8��c8����Z�c8
{c8Nc8+b8G�4�BS7^I]8N+a��#E�dZ7��C� )c83�>8�)a8VK#�C�a����7�TN�[e�L��f��)��R^L�nH��"'8�V���Q8�1�6�Ra8�dZ7�FF��o_8��B7�d�`e8n�M7�g8�Ha8��Z��,b�. l7JY7m!e��A_8.S��_Z7�ib8��d8�U��N��d��R�!U�#vY� �38T]��h��Eb���c��?!7c8ȖT��pf�I�Y��N_��Ҷhe8�}c8a\b��a��;8�wg8Jq^8�M�F�b�lWO7 9d8���y�T7%�d8�0b8�d��	�7p�^�Cf8�c��f�pm2x�T7�xF��U7@�M���_8�xG���>7�gm7��Y70�_��b8�e�]�b8�zc���a8�a���^����#n��t�kV��FZ�2�*���S7(	g8�^���X7�R7S`���b8�Za8��b���Z7�$L���Y8v�b8>�+7U78gUU���7�:e8$�T8�d�ww]8 �R7v�:�B��{Q�Od8T���{O7Sb8�R�L�\7��a���e8�^�Ahc8��X8�[%7��b��`8BT7kZ7�U8P�:7��R�y:d83b�qTL7V�[8��T7�d��+c�d8ȹg��Re�B\�i�e�Q�T7��a8��@7	�b83e8p2X7�s"�f-J7��7�c��HK��RP7Tc�5�b�'wS�1�_7��b8-]�yke8e�k��d�÷^�R�b�?]�a8�[	��;� &b8H�`8�W��dd8,"[8�pc8P0`��]�J�e8�ܷ�qf8r�b8"_�s2b8�Ga�����]�J79�W�97�e8��d���a8��P7�Q���`8�Ya���Z��a���M7��a�m�b��ua7q�y7ßc8��b��i`�b]���N�;}c8@�Y�@�b��ee�āe�XAc�emF7�M7Õ�6��^7��P�T7��/72}\�oE`�4�N���U7(
V7��b8� p���_8I7`��ld���e8їS�37�����_��^���`7� K���d86�[��b��_�����o8[7�`8څc8B�j�|�_��P� �\�K�d��V7��a83d8��7��+c8��_8G�d8(�e��)P7W�c8�;7��`8�`8Җ@7�qU��<���)�u�c8/�]�J�N��nA7pd��d8D6R7P�#_b���Z7�ZS8rIK��qN7�O�j�I�%G�y�Y8��]7i�L��z�
CU7AES��ia���_���973�c8gW`�E�8��`��f8�̖7Z����o�c�9�V7�bc8�$b���a8�h�����,�rd1Z��|Ͱ��-��l�-j�1�0+�L�$0RTW��HS1��R1,�s1{�1�r1�0��$1bL�0�7�z)�0��L��a\���;��w1#�0��i1����B��8]��m�5�W/1�j1Ͻ�B����0�5�������H�R��+�0۵ɱ����5���#��I��E/���0�̧0
؍1�^o�Z;1sō�<��0�,W��Z�0x��0��	��V�X�ݯ��㮘t�/$QP�EϰW�:0��'���q1���B��0�����,�1��00B��	��/0�	2�����Ű2�1X�����|.�y�}e�]���4��1�fc�� �\�l1���1�ł��v�����^����Ҫo0���1����
�0��1#�K��#D�X�i1�� ���7�o�� 
2��1��İX�+�꩚0�1�2O�{���p/Ծ�0�eT1���0����$�I06ڱ��@��~,�0�0&�Q�|y�����K�Ўs1���0̶ѯj1�"a���/����gs0F(��J��/���0ܦ,��+Y1���i��\b*�H�H.�~�0&]ۯrk1{{1kB���G�yR�N�?���\���1p^�.q�S00�0~�u0W�>1��0��/l8��N4�0|�ɰWP�/!h21�H��0Q/&Nc1(E���\�ԩׯ�ξ0p�1���1>�ɰ�K�0&��}k�|���5i���n0�LM�@*0D[�06��0�رb<�0p߿.�4Y1���/�����b1��.�(c��711�41x�-y�1ɂ/1<��0��:1�+��1��0�w�0�1K�1��r��1�%e0.�������� ���r��W�U�
_�0'꫰&�?�s����C1�.���|��D�M����0UZ������A1��61��Q�۱��װ<
1�S���?1&�m�>}{��ڰe&���q�X:.$oy1���0���=�/"���1����e�Nމ0�N���0cuu�����'0���	1i��1(���>��0K�W����F�/ϝ�� `�)�oA����t��֪���b�"��0��?�?�
�$D;0��1�땱�x����V�1e�1�;/y
1Lt���M�1�Cޯ�^�6�����9����-�Yа_n��mRS�j��0?��1����~\�=����_/�6�.��D���0Z�0�%V�E��-��0�hz���D1h�L1�&�f��F ��1�����V1�A1�������;�p��/���0�_+1�ѯ�ʙ00;T1f��?=���ۇ1��]��~�1��30���0�xu�L�6�ʰೱ0����K�0>��f�_<�0������/��1�M�v]�0�0ϷC�1���.p�1�P�1S�j�0�ʮH�"2�"1��Z1U�1G�15d��sj1�徱��<��i1�c4�q�/���0]�/�}01���/[R!1Z�^/�7�1������w�0/o:0rN�\ m��z�0Y(���P��</�XK16$1��"�/y�0ܡ᭰	�0[M1��گr?D0��	1<D���U1q��1_���VN��~&9��}�j��0�ޯ-�g���ʰ�C��:W�1�2!Sg���/�$�/;�0Y/0�u/����I./�Ţ�֗��8_1�4�/��ɯ^p0��1/sE�v�0EHi�X���-}����>��G��(1��ȯ	�1�O/�2!-�C�/��n�0��1���0��6�bԅ1D$T1Ep߰�%�1�sC1Yּ1���0A4$�$T�1�p��n��E�s��W�0u�I1u���\��0$�x0��.0K�/�;3�$1���P�/�W/N�#1f��0,N����0ܬ2�����08i�r�0v�$1P�	��˰���|��1�o�0Tuİ�;��@��0��3�[��\dO0�|�0򰎷n1�b�1 9��¸��Yٯ�Z��Gtw�ց��~&0|�t�\��:ð��l�I*��3>6n����#v8
�{8X�	��ld���p\G�X6·u�a8Q�8
�x�C���7�86��� �(�m8�M���d�6��9�Rϸ�钷����L3��ڞ��Nc�8K�v7�7R�Y�ύ�8p9ݸ�n�ٌ��iuf��U4���8iq8�z��ɓ87�8vc�8�8���
�t��8��l���m8=	x8V��yX�8	�i��?j8��µ�f�v8�'9j�V�<���<���p�8F��5�,�8�P�8ּ�F�84je��H��ҋj8(̓�^�8��Ƹ�8 Fv�T�k5f���P��7f����8|R�8���7�8��6�Vc���ڶ���d�8��6���j ���ʷ���8aq�����}�~��R�f�\8���� ��8�㽸̶~�|w�����6o@��F�9`�a8�Ȱ�SJ��*`ӷk��8[�͸P��5p%�5�i����8LLǸ���7���%��8 ����?�8�NM�4N���Gط����@.�54��7��ڸv�����8A$�����A���xuo����WJ���8;	f8����8S��4�\k�8#��Vj8-x���q�8Ff�����9�ZX8y����g���}�8xu�7��5:y�8�H�8��8�?��0���D��8\��8��7?ض7P�a8��޷��8����2�^�·9 ����7����8b�Ț�t�q��(���f���!��|0���C�"���(�b8�P 9{��6|�8p7�8K�޸�;7���ޓ�7@o���d 9�r8���7@�h�%��8�v�77���w�6>�O�,���<\8��b���N�b����(S7jNʸ$��8Z��� �8�:�%Nn�,��8���8�(G�B�}8�^�7�j�8�(�	��7ַc�7��7�a�8�M��;���Pu����8L1�800@7�8��i8�V9���l�b���и��N��W�6��7��8�t	8W0�7+7j&]�x9\Z���s89Ҹ�݁�׿�8ˏ8wj�7���O?�� Z�5z��	�8���79�ѷ���8�����8q�8�q�7P�8ا�8��v��Xi�D_��b��8v8�8���8c�ٷ�v��u��M�n�˸v�48�+}��b�P��8^8J8 n� m8x��7*:O7���IA�8���7B���e�8iQ8�6�Jon8����<39��ķ"<7p얷B�8�
�4-IԶ"9���˵8�9�tڷo�8ve��ZK7���d|�8~��6���X�d�.��8��ӷhW��#�Jw��	��7)��7@8��D7���ݽ�X븼W8�z9��ى6 Eb8�E��+�1�^X�8�^�����7>�j��&y8:t���^�7���8 >I7쩸��	�8)=�8��`��Y 7q8�I�$J�$֊8�?ɸ��9]�Q�>�b8;Y94O�kM�Tyx�Ӂ��t�8e��`��n;8�8Q�J��8��8��T��t8���S_L����8�`�j�8�[Ƹ�`�(4ط\9���.�8mڦ86�8���8�酸��76�G��k��7���W��8X�Ÿn����9Ǹ2�hI��)
������8���8�GU�u`ʸK���7zJ8m��8�}�75���e�9nN�Sx=7uT��v���zʸ��9Na�'ค0t�4��8�	��[��R�8���7���8�Zи��9�G�8�v�8���7���8�J������_��r2�7���7ɲ]�*�^8�+`6�f8�׆��#o�u�︹l#����A��6�Ѽ8��91o��)�d�\���f�ک���v83"�7`��7d�82x�8JX¸��e���7�-��)�8p�O7���7a�8@���W;���">|�r��8�H�8����k8�L^��(�6(d��s�7�E����82�����Ÿ�J�8���8�Dݷ�9�)�8l��8M�<n�8�:�8i��7�t���r��׺���9X38���tU�8�i�8(�7҆,�0%a��7`��5#�8���7@_5�ޞ7��7JT�7��ѷD������*��`��5 ̓6��7��$8z��L�#��dt������W׷��4jh8ε7K[8��	8P}�6t����%�78�P8`ϵ�=�6%e8���7�I�x8�}
�+�� �7�A8�tМ74��7
b���S�70ն޵��}8S��bF�8���7	=6@a�6^}�8���7ni��x� ��l8!I��"��7�J�����4BQ7T��7ݚl8�^�7�ZS�f'�8�ٶA�8��)7p�[��'48�W.�Dd28��b� a۵P�@6�ڗ8���y�8�^�I�H��K��Dw�����,���a�8X�6�h�L߿����8H5����� 37�sN8ﳸ܉������s��@��.�8b~8X�l7�݈��|�^�7�J
�)7�𴷱�y������~t8g��|�J�DIV�*p7�1�7��7�z�7@C/�eՂ��.�6P����8�o(�i8:�N8��̷FX8�Z� O�5t/��]�8����T8��7���70`%7o�3�fH���U��;T6#l�� \��V��7��07fN�7�ѷZ�&8,�74c��"�<�4��Z)�4��7�1%� ��<D�J�8��8`9K6�`�7��,�� ��7����\��L�1�6,�7tN��@]b6^70�X�8��\8~����q��+�5��{7����n���l��t���		8PjR���7��}8����Ek8�7,W5�Y�8r�7��5�>��7�g�����J���a(�h�$7��?8�vm��������8`���vJ�8he97Lb�8:�������_���ȵ�8�8�H8ʒ8v��7�X�Z#�8P��66W��`�^6����Z��&8���8�8�.s8�5�7���$\�[��yٸ4m8�4�8�P�`���7�y��(08d*&��	�8.��w̄8�b	�o�2�x?��PJ8 ������`V��Q�\�������������7l8��˷�~`�d���,�7o�V8�8�:6� a�6A7I�8h�M76G\�ȧ^��Gf�To72	3�֟��\*2�p2��H_�7|�7�EW8�8��%8��7�n�P8l�����7L�A�@
5�8|���<���ᤷ��6�M��ٝ8�=��h<x7R�78Z�S8/���v�|�߷Pr���}��8�J��"H���Y8 � 7rW�80Q�77&��V��XL����q8�U���7-�����8��8H�K���r�ڍ!8��8z<�7�g?7G�7��7yɦ���ֵ�ғ��ի8(��6�E����8\/�Н
���58���h08>"<8� ��<8}:�4���|�7��S6�����P�� 2�5����1�38����<�7���7�±�\Ʒ��8� �z�'��^�� ���X��6��v8$�/��"8 v���P`8&�{�8��6����P�L��.�+�I�j�7���5��H���S���R7�暷�I�7������,7T�帀��8$@��b8��8��4����`0�6x�H7�"��%F7��=8��j7,�P�x��{}�8p�6���874��O���G\�`�D�E�p��e���e���ڷ���,FV7��8P�N6�!�Pxηg��Ȅ�70��7��c�|u7��|���8���7��Ϸn���μ7V�!8�q(8���7L�18�[8����ޱи���7�L�7ae38Q`M�2��D*88��6��|8�(:8���8C�6������U��m�7З���7��i8D?57Γ3��I淞�����6PbL��t�7��8�ٓ�S��oȠ8�ϕ�?2�ܾ�7� �]O8hh�ܥ�7mss�|�,8�7����8�r緦��d*�\eD7*�8�8V�58^�8 �W4�U��58���8FK8�O�����%���27�	�7 ��,8b�?�k����7:��6/7�8h/�7,l8N'��{�7�l8�h�м�6,�"��/ڷ��8 /��+7����  7� ]8�6n�9׊7W�B��m�7��08p~�8٤L�>Y�\"�$��6�J8�y�.Ց8�0$�8�7�3Z����8T)8�xe8�a0��/��n]�:���8~w7@W��=V7>1%��y�8�V���T2�M�7US6a���8��K�{\�7�ȹ78b7�O÷c�8t����/�l�%8@C��>e,8��8{ƞ7��/8��q���8���7��7�O�����_C����6AX/7F�#8��8^��yWz��,5t�W7�婷,�7����I8�~[�B��6rX���F8�68Ԕ�W��8Vh�7�Q�mk>��0�7�c#��P�8�.�79���o]8v?+�o�>���6X(���܆�&�7��;7HI��[a6"b1��;��,��-�6�'8�w�l��.�g�Ͷ�&��S�g�*7��L��)�6�7b���F�^� �VT�8�qG�g�f��:y6Э�7���5�r��Ϳ����V���7��h�m�8Cծ8���$�����!���!����,Sķ:2�8�I���]6��A�ӐC8��V7�{V���8Z`�5$߰��G:�VJ���i8��'8�5��gV�r|��Y�z8m�[���;8G�P6HZ�2d�h2�7�3��l�y7�89��)\�8C
)7������v���\�B�k���6>g�&�w�oꙷ� 8�g28�N���q����]5�g8�/37��V7Քj�������������&��6*�H��7�b8�uj�Z�G����6Q#)7�98�a8C	�56K8hr�85`^�Ux�5j.��C���W�8 ���3�`�%��s%�Q�^7B������ �F��8�@�����7��18A�n8�~ɷ��5a���ρ
8V΋�ke[�G
-8'�_�|'Ÿ^,7���6�K�����I{8'_��*����8��^��߸�޹ҷ_��89�u8]'83*�8���𷴦��#��7�"�E8Vئ8��O8�f��u�5���7��9���0��3ɶ�⵶��7h%�5��-�Ɇ8��ݧ5L1�7	����렷%��Kl�)|m7u����58-Y����#��2��h 	8(u8�M����7�緙�����&�7y���:9��ƼJ��e���9�84!(���C�����hW���_�7Gq98���x�8�B8y[���t��?;��*�v�3vf�2^z8&�F8ukO���7v���M4(޻7T����6�`x��|��"�F6���8OK���8:��׍7��n8��48�Ę7h8�9 8 �6�G��BP���8�{U7���7R0�7��$����`��7"Ln6]�1co�wl�� Ƿ�8�j�>Y�7�8R8�o�6l1��CS����4K�{�P&��M�7m�4�\�7/����8򛴷ݔ�7T,�7nM97��]�0�rfa�H9�9�7�2����$������H�7f�8�q���_08�@�6#X����5�'��д�c��8�48��9~D�(Ɯ8(Ȫ6A�6��,���շ]�7Q�)��۾�V��7������Hⷰ-�8�LP�yN<�Q�8;lg7������6��8Z�!7z��hޗ�5M�e�a��럶�`�74<M8�"�59�:���>����5� �\[���;��0e7,������Ζ@�-.�8^-T�gR�7�8�F8��U70�����7�?��zт8R�e89a613�7߳��	���  8�͖�S�5�,�7Rc�7���8c�̷汨49����V��.�7ܚ8���xV�g�����&�7� U��B?��B78}18�����!�6z�[��q�6��6���
�!���$��o��8��74ll8��W8��/��t�8	��6!�8�n�����?�Y��o8W�G�8��l����7}�{�~�U���O6Ch7	ķ���8�Ⱥ8���6�� =h6 n6�8��8��{��X���8��ȶ��7 ���� �8�Ƕ����?��J�8⿾8����᫸���8���� �6.8$Mc8)�8(�{8�P�6�׶���z��8��x8�w�8J�@������8����Z����p����x�N	w��X��?��8�j�8D��8�f	7�������8@,�8r�u8h�8���6#���(Ly8�'!����m��7ȶ^�8`>��+⸸	�8��¶6N��D��7�"�t�P�x8|������8�����-m��]�7���d�8P0ݶpZ�F8�P�D����78���f��Ҷ�8�h{��6z������f��ܷ8B�~8pߛ6��8<\�8�r���Z�Q���׷��F��jBy8.8�ܻ� R�6f�8b�w���84Ļ��Ez8��� e�7�� ����N�8D����8�羸��|8�8i�8�����8���8�sV8 J��ȿv8�8�9� 3x8Fy�n����8(r�'��8t���)�6�{8�ff8�38��8"����8<���y�蚼��q��R��'m88�v�r澸����Ҽ�ij��"���8�ȸ8~{8�!|�N>u8d��ߥ6��6��w�r=�8�c��4��8<̼8�e���\q8v�8:�8�匸$|8𑩶�׸�R�8�4����"�8 <{8��8�-�|B7� Pж������s8�t�S����8�C�����6X4��d�6�37�����8ٴ�ܷ����q�  a�&�8V��8 w8p��J�t8Ҕ� �8��w�����]�8xJ|8�X}�B|��NĶv8�8���6����ݵ8�����Mw��~�����������߶���6*w��1v8��8
���v8 �����V�w�|M�8���6@qy����8�8�ϼ�B�r��W_8�N���b쵬��8�8��B���7�vv8�|���8�8p�{��[���^8@j��L�w8�W��<�{�nϹ�P�����佸� �8��8�������(8t)���?�8q���t#���t��$��X�����{�p�6�8���8��8�[�8�V�8��88!7���p8 Ϳ4����E8��U�T�$7@���b��8��8.@����rһ8 º8 �׶L�8�b�8޿y8I���R�g�@J�6Xk�� i�6C}�,��)~�8Bx�b28��y���T�@�8�j������d�Y�����|8/��8�,���i8�(�8���60��8�� 7�,;�
j�7@�~��-�8�Ӡ7��7P��^Q�A�� ��6LY��]�8"��8�ٟ���8:�8x��8 �����Az8l�8Gq\8�׬�E}�8:�8�G�8�TJ8Đ���;8ħ��t8{y��׺������6����\�����p8p8�6�u8 ��6@���� y��O8h��������.F�"�������Ò6���8�F�8�O���U��ٹ8`�ڶ�q8d�8
&��p&����6T�o�l@y��8x 7+����x���8��^8N>���8��8`�L5z8�����4�����6�Q�8����������o8����&V�_�8�ٻ6@�{�t�8�o8P��6(.��\ew8tw�7 �{�_�p��t��/��d���x���x8z��8������7�i����7�䷸���8u���r�x!~�B38葻8n[|�@V���xv�.w]���r8�X��N��r��N��8����8�H�*h�88�ɨ7^�}8j>��}8@��N��8�;8<��f�s�p��6|����7��f��з����@ �\�E���w8a����%���e8��6p�z�**�7;'��|9��������87g�8����{8�d8슰88�(�,�8�,8�8rx8��y��80��6g���:x8�D������u��U3P�ֳ�/2[�1VO� B�3���7��V[�w򢳕h��ǲ�X1�Î3�e�!抳R�2�Ѝ2Gho�~m�2B�A���׳���3��3���/�Jo3G�3�	4�]N�E�E2�3=��3��
�ej31t��tR�1�J2�@�{�2D#�3�V�����2���3�|3�Wp3e璲��#3�R3K�&�K��֩3%�32r�m2y��"�<����F�P3���3Lq�3�i�������:3H��1�d²(�[����� ��3P��34���j�C3b�x2���2��v���3#�*3�S����3._H����"��3 E��4���r�P2��3��>3K�3d߳E{����3���3���C���+3;3�"���럳��/��u���D�2`��0=|���$�p1��T�w���\��/C2hQֳ:���/�Ʋ��O3�槳����o�U���ܲ��4<�2x.3���3��J��3L�.�	z���<� Lr3 �ϱ<���F�4����64AI��6�>3�OJ��̛3֑�3�}	�r*�1��`c�p~��ؑ鲥���0�2�D��"�3ĕ4��3����] �糅>4s��4�[3Kֱ~��2_{�3^��1
��3��E2|9�3�e�jr�2�R��'����/M�W����3�8�2^�K���63���\����3Vvg��E�v�3*��3�P�3���[�^�h��>�r��2!>b35���ZD����2ٺ�2  �-g%���Q3˲�M��3^r��/���!�Y3����h`�2�[3��3:�\�N�2-s[3|��3=��S��3-�賜h2����/e��A����3��3jJ�1h[̱�|g�O����J��2l���S��<�M�#��B:�3b�T3LǲQ32���8���#�H��f�3��e�6&�$&q1�w1Y%���2�k��������b4��@�T6!�$��$[�3.��3s��|3.�R�Nh��m3�1�2@�)2H��3��ʳM�Ѳ�d�nɰ���Ӳ7Q���2M�˳�f�3\�_� ��#�F��<�v+��`��2h+D���4� �۲$Č3�T�38g�3^�3���3!�4�;�3�2�343��ĳ𵪳j5��(U�/ �2�ib����2g7X��g.���3d�Z3Ks4444�r�3]T��.{���H��3�?�z��(w�2<(���I���,3G13{��3N�g���\�0*3}����3��?��q1ʠ���X3Hš1~��a�V�3!K�3w������*3�g�2̈���%3r^23���1(䄳��3S����3�k�2��w3�W�2d~H���j�,&�3w6��C`�`چ�K5z3yw�26�3I/���p21#�3���3����3@U�@��~�K3/��m��3���3�\��J�2��p��1^3~Y{1�!�	%�2�2)���\�C2�tH�R�P����3����9�Z���;�>��3&��3j�\���]3�&���n3�(�2�4�ւ�xG�3�γ��2�	�2�S�3�Ӓ1��~���\3�$��� ���[C%3̲̱�
����GE3â3�F3�C�30�г�Ǣ�d��3���2in��,^�2k��p���_.�2.#�3��Z3b�(�,9�2D�,�
l3+�93�M]39��2'���[��kJ3�����3䉶��g3�i�.��2�3��&�Dp�2�=$��?1���4Ɠ-���x3��象�7��	3n��2 H���ɱW�ձ�}3S�53��`��@�2�����3<��2h]1��R��9���U�� ��.��ֳg��2��~3�����ñ;`�3IK��>����t�y�����3<H�1?�W3�E��u3���2����H�3�ų�Ӥ��T�3T�N1�8D��粲�\�2f��PX`���4�-�3��|���!3n�92�"v��?13���A�Ŏ���8(Q8(߃�6�������
�wε����$9��r3�7����w��W$+�c��3B:8��L�0��������7o����8$E�W9�o�8%B�y8�_8^��h=8�����8�����8(J8�
2�y\w58d8)f����4$k8�x8�g	���5����R8��v5�u���'8�8d�8��8�'�:�8PF��A
�{��6SO5m	8��8=����dµ��8�8"�8���ݓ� ��5��ߵ!Ӫ5�r;5%$��G��
5��8�K4��8�d
�ک�s&�e8	8�nQ7&�y,5���S3��51ꭵ@ˡ���87}�b�8�X�5F6u�{5J(8J$д�:�C\8�h5�}7�t�Ӳ�@8����b��,��S��E86��Ϭ�PA�5p�8����hM���d5vB
8u�L���,Ժ��/8�n8Rf�t)8�	8Fwv��?��H��gr�5����m5�	8�
�Mp�1�X��l8�	ȵ��
8��5�L5 �8�y8�8mb赦��@�2��8�l�-�	8���3��8Z�4 w���!a�<O%5���W��X}4��4~��5p��V~8�f�5b6���6�=5��8�
8�'8���5�S����5x�*6}Z 3�κ4:i� 1��`D^���G5�88 ��o����X���8i58���4F��� }8��8�ԯ�3<k5-��h/��_�4�
��1~ ���M^3�ݫ7��88�$7X�E�K��b��d��3h�'�ky8�J�h�䴺�{�u�8&�8�8(5���𥴲z�B�u5�o!��@8c���	�5M]��,�����5ʖ
8fJ���8��;����2|��z�8���:8��u�$�XZ�46�8�8q�0y54J!��)�U8S�	�*�#�q}
�
�ˁ8F	���:�
8g2����j�T�o�˫�&/�5�崗F8��8�R�5&�7�.8�)
��f�8��6h�	�࠵��^|�_n�l��H�V��8x��Q�ٵiwn�k���س6�'8��ﵲ<^�� �7'�y5sx8���Y#��X���R
6�l���)��/���:����5�J
8p 8��4c�	5m�8�^15|�5�`�,@��@�8��H��PS8�
����� �lx8s8�5��8��<��ጜ�U��5mp8��Ҷ �8��	�:~8�m8��c���58���,�Q���B	�Ʀ�~�F�]j��G?�v�3�E|5��5ߘ8�6�4:BX��m�3������Y�q@����	���е����8�.8�%����[\8�{�����0|����"8���4D�4)�5	��C8��n5��8�-8��δ2{4���4E�����@� 8]��P�.34.
88���T�m���z����5�L�5�8�h��Q8��µ�8R��o8P��''f4qs8jn8�
.6���-�53&$3���8�78�}�5���X85Q�P�8�/��9X���ʇ5Ej 7��ڵ��8���R��C&�=��887�ٳ�(�6�<
8^��l'/5��Ծ
8�8�r�4�8E����5;εw�ڶ�݄478H5Npt5"�8Z��
�7
����8xስ�-]5NR5o#���I8�Z���β7���7"Y�%a8�
��I�o�8n�15cv�5���5mf{5��8@Mb6���3-���h�!�8>���5���� �6�:�����|N6��Y� 8�����H�ٳy@8nY	8)S6�6
�R���?��/���:S6��8H����8I�8��]�/9�5`�
��G��\�
�c�	6N~���	�H0�5��56��a��� ��f�0�[~50�t�/��F�&pү���� A�-r��/���`30�ڜ0��0 Y0q�����4Q0b�0/`8�/<� 0��c��׈�E�b��ͬ���î�2�����|�?����(�/g�/�IA/�ZR��s��8�0dxȯ��0����T{̮��-�\M0n�0�]�/�\;0�6!0��@��R�0UtR0P�m�'o� $�-!��^�*0��0�v�/�Qj/�:���� �*�0f�q�$0�x�/:'���X�<i�/"Y!/�[E0pB��p=�����VH��:/M�/�6W�5�0��������F;0�0)0�"�6{��!���,�3V��1�W0�n0�e0gv�/��̯��0�@S��P�.���/����E0��ᯞ���2�]/`(�.�)��,���V� �������.k��U�Y�l3~�p ��X\�ts����0d^0�^ϰC��0"t0�x��0�=/�ڋ0�fN0�=��f��/��/����@�r-�ȯ`�j.7�3b��΄�/0�0տ	��xy�)�/ɚ0 ��/�%Q.�UB����Q@/4C��R�T/l�s/��$0n$����}0�h�{�z����/�N0���/��8/,�I�f� �W�/�����{%0+>0٤�.8��.�����M0��/��0��# �ܪ�/Y�
���z.� �0����ϊ�bS/����~M0�%0d��#�,�y�R�x����/66�/zv%0 u-�j���Ή0R�/��/������/܏/��+0'�0�C���02�)0~�0d���~R-��/t�/J$¯�!10W�"0��������u�Q��/��0�Z@^��t�0ތa�w���e�bA����-�&�x��[qP0H|��`W0�$ɯh�8�� a�Ќ
0P�2.���/z�4�VF����/�[�.��e���p/�e�����P�0��0=L0�s/�Z�$q�/��/���/;��p�t�|@�/ �,�F8/��:/�N��l��.�i�/��q.���/�ЯNYl�`K�-��V��D&��u0L��棯m�0���д{/@m��d�A/*��/�^01010���a�YQ0{:0H�?�L&�/�.
�0O4��\C��2G0�d%0�|"/(9F��i�/b���-�/���^�0#	�/6�/�W�� ��0���*�0�-1�/B�ԯ�c50��-'�0`o0�NO� .,���	Ze0��-�U����L�JS��a0,�R��츯`(m.�q/=�J���[/��Q��=d�F�	��T����.���/]U�0�E�/TP�8ꀰ��.X,���p0`>0�D���uw�*5��B��.��ӭ��_9�����,�����������/ P!.H�����_�� 0d��0IۯJ�-/������մ*0k00��@�l/�ȯN7����n��80X�a0(��/;H�/`���/���/���,�/���/��N0��*����.�2/L�
0�]/8y<�h0&��s$�-���>���yO�)#0�e0�ބ�Σ6�>|����E��ޏ/P�.`�$��Q���_L�̷"�@|��F,8�����b�.��l0]�/ x�OI�B�ϯ kׯz�`��^d0bj0���/ �^�G��i�%�A�H��0��/_)�ֈH0�f��߈ 0�*0��0ɯ�k�d�l/UK�/�
�������:���0�WX0�|0q�?�[�/y��?���_��B��c�#_i0<&:�Z�/�1�פ
0�-0��r0���/��/6��B�m.y�0�d�/��0w���x�]�������ђ�"����c������<���`�.�ǯ�0���h�/!��f��/�^@0���D`$05��/��[�5?p0He�/ �q�ࣚ.�﷯8��/s-0�.��}/�Wد��5���0;�į;f0�c50Ԩ��|��u=�]{����0�zz�3��/Cϒ6��@�fd��"=�`A�Ԅ��V��6�^@���?��A8w�6 @�E�G8�w��5�6o�B�f�>�f!��G�98�/Y��/���?8�|�6��D��/?��l�6�|k6I�C8��68�S�QL64�,�D�6�5�5ȃc6R;8�܂6�X6���7�fD�YVD�4BB8#�D8(�7�/t6k\08*MA�����aNR6�;�)u�6q�v��ED��*����f6Rb�6�m���(!�i,X6�C�.�t6�}?���D�q�V68A8� |�B}�Q�;�_�?8
B��'���A���6�cE��B���6ǭ>8,93�3A8^x6��B���B�Efr�	v�6xp����$6�ȷ��C��ED�0�n��T��S�1�k�6�-@8������=��򨇶�i�S�}�܈��kD8�0�o$?�qF6�LD��I��ـ@�d'��j�D�A8�?��S��gB�>s�6��R��jD8( t��</��I@��Pk6�r��lq6'@8ʶ?��hV��B8�rs6ʑE�v�:�r�+6�D87�;6��C�Īa6ȵV����K�>8n@8uD6�*C���A8�1{67A8�Wo6zC�Y��|
�O�?��%o6�,D�G�M�����B8fy{6�=8W�u6Z1B� oA8�D�:4J6��@8��@8M��'G��W6a�6g*8�G8��C6��6&�h6V�6-�P6!�18�@>�F>��C8<�I"���C�2;8Dh8˘l6�B�l�A���7��b�8�5A�\b_�Y�;8��B�J�<7>;s�(?8*4D8BD8f�e6�A�����cS��a�)6�T=��zC8�y67PF���>�H�?8��Y6�j�6̱B��F��営a- �h#<8+s=7h�;��i`6C�A89���k?8�46$)@8�r+���7��C�8�@��6t�ˎ�7$�h6�JD���6
@F�c�C� mC8C"�6|W6��D8=�G6�]N�[L6�C��v{���;�:����@8�*=8�n6]=|������r�>m7��x6�+C8Й��B�1�S���F6����Kfe6�q7���6��(���p��]A8��9���W�r�B�I�8�9���ً6���%hD8qY#���"���C���*6�FF8VSB�&\C��]�6q��7��C�?�@���(���6OF�6(�;8�Y6�
B��G6KQ?8��7͍:�w�y��*?8���6/w-�}.B��zC��)�7��5�}�7�ى���6~RC8S����}�6�{E��Y?8�f����7�D8�S6:`A6�D8s͎���<���D�C�6)7b�n88�&�6kK@�Y`����7�6B8�@�E8��Z����0Z����M6�5r��s;8��k��`���|m6]�E8�A�ң@�$�J65�:�k�F8���7z�!�����#��6_?�lЃ6�C�h-6�;E8��>5|�A���_���@���A8��@����7������� D�� P�sB����|6��E8u-E6��.8�G8�r�=86�B8��V��VB8x0�����q�7q�K��z@8��>��my6�ⅶZIN�6��]��6���6ӡ?��f���2\6^�@8 ��5��U��=� ��5{Uu��b���C��$��r���&�DQB8ߝ�/B�6�98]@?��D8$�S�V�	8ӓC8�F��MA�r�0��lT�[>8��8�D�|����(C8��s6��>�$�A�Y2@�jv-8��>��o�ʬ���PB��@V�WR\�� *���Y6)�B8M�?8ftQ��=<���`A8�>8hB8�6>?8�A�=�<�U�@wD8<�5�ɷ@�F8K�F���6�rG~�ٷY�t8\�@83jS6F�H8�q@���6��8@�D�q�U�9hG�"����?8��D�����r�?�^;&8,fA8fv6Q4���^�6�t��I�/�p6�6}6a6�;7�f58��?8.�)���C��@8�CD��B8:���u@�)e,��e%8yiA8�c�?�.��TA8��F8�_@�zY@���_6P���-P�5+0Jń��˯�������J�P/�� ��:�-�i�/P�E�Z�0r��/\��.0P��/	�e/���,��/�E�/��� �5--42��Wg��B0hHe.�	�a,����/���/��=/	7�Ο_0J�x05�0�8�,�(�/̆���Rįox���0��}/����S�z/(2�-u<}0*<y��G� p�&�0�k��(:�����0ն'�v��.:h�dy�V�o0�/W�W.Y5ɭXm80���/B�ׯ�_M/��i��\tO/+�������s�/���V��/ۂ�T��b�m��в.�1�0!��Q�\/(�8�ܗ��r�ǯ�q0R��Rw02k�/�IݮV���/<F�.U=��-8�>`�0���.I��/N=O025��,����M����0��0��/jb0��X��$�/��$���1/<���ߠ0��>/��n�8�'0��y/�T)/��&������0��X�l7-��$/s��/j/�b/���Trk�Z֯��p09H@/h�����&��,��p.��Q��������> 0X��/�>+�d$�.��D�1ف.���.R��/)���]o'0b��/z���/ގ�-*�(��j�- d���+E�:�70n����60�).~�^02���-�H��/ӡد��z��4/�v�4�l����e�M��� ���N0ߦ0�ć/uU7�&_����	p0)�N��ɴ���/~��ր	.�̨�<= �BR����ǳ�0����Br��W�-���/�?�/�Թ.�\0�j�.G���W˹.ljt/�kG0p��0�Q/���ޞ����c���B/�Έ��A/��/w��/�;�[ί�!����.&{ޯhԲ�ZM���T�����Q���
0ct�/I��.�0]���@U/zׯ�%�/���/$;��l./+\4�oH�"߅��a�IwZ�ѡ9��!0T�/S\v����'Sѯ�x/�f .{`G�S���U0�%V�/K��!0�W��/\;0���g����/��#/�똯�)�.���d�/��ѯ�����bx0wD��DÃ�#����P篙vA�8�|�L���t�.*S/6g/�F/(�7�į�U�/JZ.�P0����M�ͭ/&(0Fy5���7/��"0wJ��S�&�J0��.��
0u��0��o.����B��.��&0��W�uZ�|��-k;	�f�-�#����%/v���NŜ/X^/0���U���N/��+��g%0�L0��P���=/}� 0�ɾ��0z�m.��\���o-�;�>o� t���ّ/��/�07w���>0��4��/�X0�?0��j���40&�T��ڸ/�(/�8��0�
�/-�/�K\��O0F-~"���9*���zƯ�qB-"uR��uP0�E���a0�g�<$S/|u'0V��/Y=�/2�0ۋ^0[4$/=�x�	-w�8׵�Be�/gx�.�µ0,1��ڔ/�ĳ���@��A/���0�p�n6�����66���/(B�|�k�C?�\�,/��j�'��/_��/�F���?.��/C̰/�L0�SٯT�0�Ι���)/
1{��k��В��50�-Ϯ�C</,�M/ML/�$)0l�ͮ>��ү·.�H�0�6�/��/���/N�0Be8��.FT�/)�(\�/�(/,N�/�i*�n�>0�$�c<Y0�_����ܯ��S0?߉0�;ү��/w+o/�/l��Y]ܯ��-^L���J�l0��t��-�5)�V�p0��..g����-*��/ޠ;069�0�|o/^Id/`��/��
/३+ɮ;/9ܴ/�dz0���/@4e.r&!0	z�.W	0/��f�/nă�S0�Z�/���/�k'��=���j�4�:�<�.��/�G0i�]�\	�/��
��_S�o[��80�uq/��;�8��q���/ɯ,��r�0�6����=�.S�;01h�G�0G����y�/vK
/p�*��<*0PKQ���P� P� PK                     0 checkpoint/data/29FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZi��4�e�4���4qՆ4�0�4c��4q�4ZP�4K�4��4a�4^�F4��4�1�4e�p4)1g41>G4x�R4"�4�l^4��4�G�4�
{4��}4�O�4��v4v�4���4=\�4g�4)��4�O�4EZ�4��4�J4ț�4�K4��e4a�|4�l4���4�pr4	�4�_�40�N43�4�>�4U4I�<4�u4_m�4�3C4J7O44�4W\�4�w�4�o4@�\4��4�n�4ݍ|4~֊4nI4���4(�4�X4Ç4�_n4���4-Ą4o��4�Æ4�z4.[4�Uz4���4��~4K�n4KU�4=(h4_o4Vȉ4��t4*��4�'�4�W�47��4 nM4�%�4��[4F4$�~4�g�4�щ4���4xq4��v4H>�4B�d4�;4m�4㏆4��r4d�4ʊ4
{�4N�|4��d4�4��|4��~4j��4t�4v@4���4�-!4?{�4(�4˰�4!4��42WN4�44��]4I�4r4ߖ94쁄4V�4�}�4�q�4gh�4�DD4ק�4��e4�X�4XX�4�4�4Y>�4yh�4��C4�]�4��4���4��x4d+Q4�D4S!~45�4N�4A�4n"�4�(�4��4�&�4C��4��@4�{u4�@�4�~�4vis4cz4�5�4�4q��4>Y4�	�4�W4@�N4Q�4���4SP�4>H�4��4E��4���4�|4$m4��4�!�4��40�4y߄4l�4u��4�]G4��4��V4,�>4�܇4�j�4tBl4���4�7�4�z4��e4Ei�4�L>4���4�vL4K!^4O~4�o�4���44f�p4`B�4���4� �4j�4Q�4�gs4,\E4�q�4��4�'4S��4��4b44�)v4�}4��4M�4D�4 ��4-i�4��4���4%�4d��4��4'2�4��s4 �4���4��w4�$�4��4F�j4w��4I��4���4���4מ�4'�E4�_�4�X�4fst4zXF4(J�4�l�4KI�4e7�4Y�4�}4��Z4��B4��v4HZ4�Ph4^݁4\�s4{a4���4��p4r�D4~p4dV�4�bU4�c4@�4��4�4�D�4�4�y4���4�0�4#�4�)�4��4yŀ4��4��54 �}4��4�4�T�4�4z]}4Qx�4�c4���4k�4�4�U�4(?�4�R�4q�4�Y�4�}4<e�4/��3���4/"�4���4��|4�L4FLl4��4���4��49�4�Ǆ4�Nx4`��4�r�4�!J4�a�4/|�4ނ}4߳N4�
�4jy�4��I42J�4�4c�4xǀ4�ć4q��4�Kt4��j4�/�4[$�4��v4=�4}��4��O4wg4��4"Ǌ4�*�4�j@4]��4���4��4�A�4a��4�T�4R��4�OS4�&�4�3i4�t�4/Y4�s4│4�ނ41UW4k��4���4i�4X��4k��4t�4��[4�{4�zR4>��4��4*$�4P��4P�4��\4P.�4���4��3s�4�W�4�\4�&�4�Q�4�E4���4��4ƅ4�ȅ4�h�4�pA4���4���4��y4W{M4Q��4�~4;P�4]�Y4Ý�4"g4�@t4��4.L@4$=�4�l4�y�4��t4��4�$U4��4�Iy4�0S4�&�4�c{4=�4�4���4 �y4��4���4��|4��4�΃4۽�4��4t�o4�І4?Ӆ4w�4N�j4ui�4_�x4dE�4��t4���4rބ4�HK4��4}4?G�4eSu4��n4w�4�T4��D4%��4�V4�{4�n`4�4㋄4��)4b�N4Q��4P��4�m�4In4Ar�4���4ۆ4���4�Ղ4��d4�у4o)q4��4�ׁ4��4��4ކ4r�4U �4�/�4�V4G�4��4AIn4�+�4+9�4N�4�%�4ʇ�4�{�4��j4e�}44��4�s4(�4e�{4�ۀ4���4/h4+�;4�́4t��4Fك4vB�4W~�4]��4�n�4 6�5Z��5s�5l��5�3�5Ic�5���5�$�5���5N~�5���5f��5P��5�j�5���5��5��5��5���5��5��5��5a$�5'_�5�x�5g�50��5���5���5�W�5@�5R��5v�5=�5��5A��5�w�5��5;{�5y��5�x�5,�5��5o �5a=�5QT�5j��5���5��5]��5��5�a�5�,�5��5��5=V�5�k�5$��5�
�54��5 ��5���5�d�5��5Ľ5��5���5~v�5���5��5���5!�5��55#�5�?�5-�5��5¨�5.�5=k�5~�5��5p��5��5A��5+2�5}��5��5UO�5.c�5�W�5��5j��5X��5���5�Ϋ5;��5�@�5���5���5���5���5�`�5?O�54��5��5Sf�5>�5_�5 A�5��5�ʹ5B~�5�=�5u��5��5��5���5�k�51	�5�:�5���5$x�5h�5�&�5�:�58z�5#��5���5��5A��5�Ź5�٬5`��5`�5��5C��5�8�5��5,X�5l�5�V�5}�5�(�5���5��5�1�5U��5q��5A8�5<ݲ5��5T��5�K�5��5��5��5O��5�+�5e��5A��5���5-��5�+�5ˌ�5���5�`�5:"�5{��5B��5k��5^��5<��5�t�5�/�5�X�55Z�5�9�5p�5���5 �5���5�3�5��5���5}�5闯5C�5�,�5��5Q�5��5D��5���5}��5h�5�ܯ5���5[��5��5��5��5^��5��5��5|b�5�0�5jG�5�%�5���5��5�3�5�5�"�5d�5l��5���5��5+��5�'�5 :�5A)�5+��5J9�5bW�5w�5��5�^�5��5
��5���5ֶ5��5J��5Z�5D�5�y�5-�5�	�5x��5%��5཮5���5l0�5D�5LF�5�w�5���5"��5��50L�5�w�5,��5��5Jx�5w��5���5�d�5���5���50à5Ľ5f/�5��5���5|�5}�5H7�5X.�5���5~�5ȴ5���5(1�5VZ�51x�5Ra�5�߲5ψ�5v��5�>�5�Ю5�ٵ5騽5�5���5���5h�5/��5�H�5�~�51s�5�o�5�ƭ5�n�5_m�5�w�5Ğ�5s��5�Χ5F8�5�n�5C'�5��5�<�5��5��5%��5C�5h�5>Ĺ5�"�5��5�N�5h��5�b�5���5Eh�5�5ۻ5���5�-�5���5���5���5"F�5��5T��5|�5y:�5=��5���5�k�5�t�5 w�5Χ�5�d�5}Y�5N�5�/�5Y�5�Z�5;Y�5��5��54�5���5�2�5oP�5tI�5���5+V�5�~�5��5YG�5ؔ�5wF�54=�55�5���5uݽ5Ɗ�5�"�5�n�5��5�51v�5��5}�5�T�5�m�5O��5&��5���5r��5�5
3�5_E�5�5\S�5���5p��5�A�5���5~�5n�52��5�%�57q�53�5X�5���5wt�5���5�ٮ5Z��5�Q�5�ҿ5{��5�ھ5'��57�5���5�Ґ5yg�5h�5�̰5s��5A�5'��5���5e��5h)�5}�5�h�5uW�5��5�;�5l��5�+�5��5^�5���5��51�5ճ5�/�5;�5�~�5<��5c��5���5z��5���5D&�5�ټ5���5�ֿ5@K�5���5�5Y �5�۽5���5�;�5��5��5�Z�5�D�5y�5�o�5)4�5n�5���5]�5�޶5$K�5��58C�5���5���5^Ժ5� �5���57B�5���5aH�5��5�;�5	��5�۴5���5��5՛�5��5�0�5{��5b[�5�j�5�q�5�h�5�b�5��5!��5OL�5���5���5���5��5���5��5Y��5ļ5�,�5V2�5���5���5�,�58��5J4Z�4� 4��3��3���3=��3�v�34�:4�	4�2
4b�3�4�46L
4(�4�s42m�3	4��4��4�4|��3��
4k�4���3d�4p�4kr4[&4�r
4��3���3��4���3���3~\�3d*�3xk�3S4p��3���324mz�3+�4���3���3͖ 4#g�3�F�2ɻ4e� 4�G4��4�= 4-E
4'
4`�4.�3�p4k[4# 4q�3�04���3��4;�4'�4G�4E�3�3_,44o4���3�;4��4�o�3Q��3��3��4�r4�W�3���3��4,�4��4�~4+ֿ3�44�+	4[!4�
�3Y4�2�3��4�(�3U��3)�4`��3�m
4/4��e3\�34���3f�4�4�s4�4�/4$�3�Y4c��3�4��	4冟3�4�)4���3D�4��4��4zW
4�e4�^4��4�@
4V4�
4��4M�4 �4Ѯ
4e�3�i4��4L4��4\]�3=�4�j�3|n�3�4�$4C�4��3ͨ4J�4׳41{	4�G4'4�`�3.�4�4_�4]ڞ3_�	4�&�3��4܉4\4��3��3��3v�
4\��3c��3�4J�	4�i4�v4�4�q4w4� �3&�33�3�94�34X��3%p�3�X�3_�4�(�3Ϗ4��4q 4��4$��3�4�4�S4�Z4q�4�)4�� 4�q4��	4&�4�	4��4��3%4c64Cj4�Q�3�f
4s?454�%
4ہ4���3��
4��4$�4�A4N�4B4��
4IB4��
4�z4B��3�u�3R1�3T.�3n�4��3�/4<��3�?4�u4G��3�9
4�V�3O�3�4;-4E%
4��
4�;�3 4�^4?}�37w4��4#��3�M4!#4��3��3�4��	4F�4{�
4��
4���3�3���3O�4�C4c�
4ϥk3�4�
4�t4B� 4��4��
4 �3�~�3�' 4��4}}�3�M 4�4�[�3��4#�3�
4�j�3�
4g4hz�3��4|T4-�45��1�L 4N�3OS
4�h�3a�4|(�3�
4�g�3���3x�	4�:4�4��4��4�f4T4�]4v�4�4��4�^	4��4��3g4(�
4��4R9�3E4څ4��3��4WB4�{�3�z�3�G�3��3yl4&E4�C4�47p
4>
�374$A4�
4�4��4��4�(4�94G'4��4c)�3��4c��3�4ʹ4LS�3lc4{��3*74J��3#t4(��3td4�
4NG4&�
4�� 4� 4p4�ƶ3Z�4��4�I4��3�z4i4��4�	4�4��
4��3L� 4��	4?2�3��4�8�37� 4��4�}
49�4Lb4�4��4�g4�u4��	4���3}4�	4���34��4Z4]7�34h�3ʧ3ފ�3�7	4��4��
4���3U$4Ʀ4�g�36g4�d4F�4�
4��4U
4p�4��	4L�4܉4pZ4� 4.#�3~�4Ŕ	4��4��4V��3��
4T4�q4�74�?�3���3��4�U
4�3 �48�4%�4^z�3��4Qh�3��4��4H�4Y� 4�4ɵ�3!54ΰ�3�v 4�Z�3!A4:6�3���3�*�3��4�]�3��4�v4�)�3��4��
4\� 4X��3��4fm4��4�4�a4�4�4F��3�[4Dy�3�ʽ3�4vq4 �3��4���3���34w�3Y�4�3i�4'4�4�H�3n�4��3�+4�5�3�
4��3�_	4i:�3��3��4i�4�r4�|�4�4�+�4��4�\�4H�4P��4��4���4w8�4X��4 ��4Z�4
�4r��4ݢ4��4lϠ4ɖ�4�4�r�4�-�4�1�4�p�4�	�4�+�4��4^��4Ѧ�4Eә4a��4p��40��4ƽ4;��4W��4D�4V��4��4�4���44��4+��4&��4���4!q�4�T�4�X�4,��4��4j�4q�j4���4�.�4ŷ4���4J��4��4���4���4>��4 ��4�F�4}�4os�4_��4���4x��4yߵ4���4��4���4�ɴ4X�4�X�4�h�4��4��4v��4���4T��4�J�4;��4�/�4
q�4�ұ4c�4���4Q|�4Ѱ4D4�4�+�4�,�4���4˰4U��47��46y�4$3�4ﮘ4d�4��4��4qմ4��4	-�4�2�4џ�4���4Y��4�֥4�H�4�z�4�5�4+ڸ4Q��41��4�4+&�4@�4�p�4��4��48��4{c�4�Y�4��4ݹ�4��4�A�43��4��4�;�4_��4)��4�@�4���4�?�4��4`�4M��4k�4��48��4��4Ķ4�n�4��4Ϻ4���4#�4��4��4@��4W��4�W�4���4��4���4o��4�m�4�K�46�4ι4��4���4+�4���4� �4��4���4Bȷ4$m�4�8�4��4��4>��4s��4U��4wպ4��4!G�4��4\.�4�͵4���4}�4*��4�_�4���4�d�4,լ4^Ҿ4�˻4�]�4���4̊�4��42~�4\Y�4���4P0�4��4��4g��4�k�4Ѕ�4t_�4���4o|�4$ֹ4UV�49��4\�4���4��4E�4��4��4���4 j�4��4z��4���4��4.��4[�4���4���4~�47A�4�$�4�b�4?��4��4�j�4o8�4�Ѵ4A�4=ͩ4w�4���4i�4�S�4��4���4&w�4�ެ4�ݺ4֍�4��4���4���4��4��4m�4Б�4�@�4���4���4���4�ȳ4��4^��4��4?o�4� �4в4��4ٷ4j�4V��4�װ4�0�4�5�4R/�41F�4
��4L�4)#�4Ng�4&�4ݬ4礍4�4Y�4�Q�4h�4-v�4��4\�4���4RV�4�3�4ӽ4泺4i��4Ӆ�41�4��t4���4<�4���4��4�n�4��4���4ڐ4��4I��4X��4x�4���4\��4���4-��4�x�4��4<�4���4թ4O��4�7�4\f�4�m�4?W�4]>�4`ɷ4u'�4�p�4�˲4,1�4s��4ƈ�4���4�F�4캶4�7�4��4t�4Ea�4^0�4#a�4>P�4Nӻ4{��4���4��4$�4*��4A��4��4va�4���46��4��4�4���4�U�4��4ei�4��4�4iα4}:�4���4��4��4��4;�4G��4��4F+�4���4��4�?�4���4�@�4��4���4��4d�4ú4�4�k�4�5�4���4u��4_'�4x�4��4���4��4�і4��4��49-�4YE�4R�4y9�4���4�=�4�F�4xp�4<O4�G�4�Q�44ر4�i�4�ͺ44�4�o�4v2�46��4��4)�4�m�4��4}��4�۫4XǱ4cۤ4�W�4��4�9�49��4��4�;4s�4���4
�4nٱ4gM�4jz�4O�4t�44O�4�X�4ǵ4�T�4�ó40۝4bU�4tn�4���4_W�4���4�ٺ4j�4���4[��4��4���4h��4n��4���4�!�41��4 )�4��4"��4N��4�4���4]+�4:m�4��4ڽ4�J�4_��4"з4
�4÷4�
�4�$�4��4�4|��4�ϵ4Y�4|��4%�4c �4��4��4���4�Ǯ4&��4Rf�4�4:ɺ4+ʨ4��41!�4PϮ4K��4ǵ4[ж4C��4�w�4�5�5t)5�5M5�c 57!5(�5i�"5�5�5O�'5f�5~B5j�5"5�c5|5~5�C&5�%!5;�5��5g�5�]5tM$5��#5 5��5U�5V�5܄!5��54�5��5^�5r�,5r"5ޕ$5�5Q�5��5W�5�(5��5�I&5��5�C$5(�5�U55i�"5>�5J�5�%5��5SB5O5w�5�Z%5�5W�"5+�&5�52s$5��5�$&5g 5��5�5;�!5�5}�5�5B�5�B5�!+5�+%51Z5@�5o�5q5���4Ӡ$5)�5[�5(]5�5�5=}5k 5�_5�='5 �#5�<5/�5�5��!5�$5�5��5�U)5�5?_#5��'5�Q5��5�+'5�)5ˤ#5�5�h5b�5L�#5Sf(5��4) 5�$5��5��5�p55n"5B0&5�(5!# 5�#5U25�5��5�0%5*$%5'�5k�(5�5o�5O�535��5@�$5��%5�!5�	5[�!54R5]�5�5��5I#5�(5��5� 5�'5�M$5j(	5�<5�15��)5'�#5>�!5)M5�%5Z5E� 5'&5$!5t0"5M�
5�45��'5�&53I5.#$5Y�$5�5�[%5�N5�w*55�5�5ž5]L5�t 5��5�I5mB5:N�4�w$52�5W5�5��#5h)5}�5I5g�5�-5]5�,5�@5h 5]�5��#5!5�K"5%}(5�o�4h�'5Z�#5D0 5�%5�n%5a�%5[5�5��5�	5/�
5��53�5��51W5$�5�a%5��5n5�r#5��5�5!5&�"5��5~5�:5$�5��5�$5�O!5ea5l�!5}�5�H&5��&5�d5$!5�5��*575x�5>�5��4��&5�,5��5�65��#5eP5!�5��#58"51]'5b� 5�5�%5�q5�(&54!5�!5? 5�5`�5�d#5��5��%5��!5��	5��5��5.b5�5�H�4� 5�)52+5�
)5�<#5�{%5�j5�Z5��)5�t&5
Q5��(5G�5-� 5�$5��5�75�5tg5/��45lo%5 �!5
�#5�<5,9!5�p(5�= 5�V5��"5N%5L�"5��%5Gb5��5p�5�U5,&5$j5�c5� 5*�5cw5�M5�$5��
5<9$5V�5`&!5H�5��5y|5c�$5Za&5c 5p�"5�]$5�B5�0 5$*)5^5ҥ5 �"5N�5�5u�#5��5Qf,5�q5-�5�5<45��)5�=$5���4�
5/!5�5!{ 5I�$5!�5U�5��5�5��5�	5&5�5�5��5q�*5��5�C5=�!5"�$5�d5\5�H5��5�K5�"�4,�5�'5?�%5�x5,5E�5��"5�%535x5 �#5ˌ'5��5�!5S55�5���4dv5	5y�
5 �5M�#5�!5g�4�S$5B0!5�5�'5s#5}��48�!5h�	5��5��'5)(5l�"5�"5�5 �&5�$5� 5��$5��)5�� 5d�5�5�E5,'5#p 5�#5	�!5`S%5) $5c}5'v5�d!5z�&5�5%%5��5�)$5�B5j5�5�G5P5�"5A5S6*5H�5�A$5��5�5=
%5ۈ5��5ˡ5��5��	5tO&5�#5?�)5X> 5�15��5m�5=?"5�5'5"�!5�5�*5i^!5��5��5ܿ5/�5�5A�5Y�)5��5�+5B
 5o!5=�!5b5I5%5t�5s�5�85��(5��"5�p5W 5�`!5�t5~�5?/$5��3��3Ʉ�3���3R��3Y��3:��3��_3n��3X��3���3��3��3<V�3Z2�3�Ӳ3�p�30��3n��3S��3�3��3�a�3��3i�3�)�3���3{��3��3���3?]3���3��3���3���3���3 ��3	@x3�w�3z��3�f�3��3?��3B1�3&�3���3�k�3i�3�:�3��v3���3�
�3��3���3�"�3Y�3��30��3)��3�(�3��3[f�3��3�9�3i��3z��3��3EVU3���3X=�3���3 ��3��3��3 @�3���3e]�3���3l4�3�	�3s{�3���3�,37��29|3��3Q#�3�&�3��39�3���3d��3�
�3�*�3}�3a��3���3J��2g��3mY�3.��32S�3�'�3���3j��3~��3���3�E�3��3 ��3|Ս3�eg2�@�3�P�3���3N��3j��3���3�#�3��3�V�3J�3��3a��3���3�Z�3v&�3G�3�M�3��3&��3$Q�3�r@3|)R3]$�3��3r�r3��3���3U{P3y�3 �3��-3�3XH�3���3~�3[g�3�v�3���3�%�3�=�3�3�3�X�34��3�t�30�3��3餂3A��3n�3@%�3��3o��3B��3߼�3���3��3g��3E4�3�i�3X��3�b�3��3o��3���3=+�3���3�-�3�K�3s�3�3��3S��3i��3�/�3f�3<��3���3.��3�ه3�>�3�@�3O�3���3���3P�z3ƽ�3u��3��3
��37��3���3�l�3ǽm3U��3V9�3�OV3 B�3���3���3$��3s��3R�s3���3�}33=��3�#�3 ��3~��3���3)��3B+3B�3��3K�3�]�3�e�3���3_��3���3f��3wg�3�%�3���3o��3���3��3�
�3�5�3^k�3���3R��3���3�F�3��3�w�3A��3�ד3#�3�3\�i3b��3q1�3���3��3d�@3���3���3�%�3�`�2�E�3,b�3���3��3*��3���3�B24̇3���3
�3l��3I��3��3!�33�3J\�3|��36��3^�3��3���3-��3m$M3�6�3�x�3W��3A*�3���3��3��3]��3��/3���3I��3�Y�3 �3��3�K�3���3l��3K_i3���3���3פ�3Xc�3&z�3���3��32��3�.�3���3N��3���3T��3��T3e3��3��3L��3���3���3��3���3��3S"q3���3 ��3��3zQ�3٫39��3;��31��3�p�3|^k3���3���3�G�3�"�3�Q�3"��3=7�38X�3?��3��3l�3�|�3���3D��3��3�vA3���35�3���3�3�+L2�=3���3��3���3�3�3+�3�
�3S�3
�3���3�x�3
��3�#�3�,3���3Ӧ�3���3��3���3� �31�3��2i��34��3���3�:�3>��3l0�3u�3�(�3Ç�3���3���3M�3���33��3�0�3�H�3�Z�3$_�3�t�3���3I�3�_�3ʃ�3_�3�.�3�#3���3R��3�m�3�{�3� �3�wp3ki�3���3���3�p�3���3���32��3D3�3z�3���3֔�3P��3��3���3;o�3���3��3$ȝ3O��3z��3���3���3<�3y��3R��3��3�U�3mP�3H�3�'�3Ϯ�3���3\��3�%�3�ɥ3c�3�i�3��>3�H�3��3��3[z�3-��3N�3<!�3;�3T2/3��3}��3r3�3b�3
_�3^��3_�2S4�3hM�3�\�3��3K��3��3���3E
�3<k�3m�3���3M��3���3M�3��3+�3\��3���3Wa�3a��3�3o��3��3x��3���3���3^��3%Q�3�\�3@j�3$��3���3�r�3���3�3���4���4��4��4�/�4x��4X��4eĀ4J�4
l�46C�4E��4�k�4�`�4+�4&��4i�4�
�4��4���4g�4��4��n4q��465�4s�4�΋4��4�'�4S�4}A�4���4�5�4��4�ق4Ee�45�4_×4u�4�)�4 |�4�7�4�4�A�46<�4(�4�Ȱ4�X�4�-s42W�4I=�4ם4�0�4�v�4�Ǚ4��4��4\ӈ4�4n.�4%�4�'�4�H^4�a�4-\�4�A�4�A�49�4]�43&�4X��4��4jX�4��4�Δ4�Ô4p{�4��4���4��4㒟4��4���4��4�B�4�g�4�R�4���4ޮ4�y4}Fl45��4���4�v4/��4_��4��4�C|4x�4kZ�4���4�=�4�z�4�`�4Uˇ4�ˡ4d�4�Nf4�\�4��4P��4���4qb�4#}[4�_�4+��4�4��F4�4f}4��4!��48��4�(�4���4)�4��r4�ޝ4��4v˨4�|�4�t�4Q͚4�Ԡ4[4�>�4�^�4�'�4�u�4}��4bq�4 Ϝ4�I`4���4�g�4�O�4J԰4b̓4T	�4�m�4YN�4Os�4và4��4Wu�4��46��4E\�4t��4�ؠ4��4�$�4ۄ�459�4;=j4�O�4�ѥ4�4�4���4<O�4�W�4H��4v��4��4�ب4���4��4Q��4)!�4y�4[ǰ4/b�4��4�ޗ4��4{կ4N�4�	�4#C�4��4���4��4���4�y�4�ߌ4�=�4�w�4�X�4�Xn4���4�݂4�Ў4\�4�^�4��4�'�4���4�46!�4Μ�4�B�4�Nx41Ӎ4��4tM�4��4M�4�/842͜4���4�4G��4а�4���4���4���4�M�4\X�4a�4��4{�4�!�4L�4=��4vҖ4��4��4�]�4pm�4v�42(�4�4�4Iѥ4 ��4B*�4E��4AΠ4
�y4��4q�4��4�F�4r�4�g�4p�4Vw4�:�4r��4���4X��4�ɟ4�i�46Ή4~[�4�r42��4MX�4��4QE�4��4b�4Ig�4آ�4�Ģ4�+�4a��4]ӗ4�Mt4���4���4�[@4t�46`�4���4EQ�4��4Hs�4���4�z�4�C�4q�n4��a4��4�K�4�4F5�4��4u��4�׬4�f�4|�4�(�4��4�u�46��4��4	l�4�A�4�W�4ٝ4���4�"�4�י4(��4sh�4���4�B�4"7�4�/�4"�4e�4.��47��4��T4`��4��4���4D�4eu�4nP�4A�4��4�{�4��4˅�4׳�4���46��4]�4�Ԝ4ɩ�4
��4�Yx4':�4r�4趘4�˟4B��4���4�У4��4���4�K�4y�4O��47j�4��4���4��e49��4���4Ј�4\m�4�˙4J�4�G�4i�4Iے4�&�4� �4.w�4��4e��4��4�b~4Nқ4���4��4�4	�4��4��4ơ48��4q��4K�4�}�41.�4��4�>�4D�4͕4+�4�9�4�k�4���4I�4ǡ4��4���4�!�4gŋ4�?�4�%d4���4>�4�}�4���49 �4c?�4�Y�4�<g4J�4�:�4��4��4n��4�~�4�ŏ4Mt�4��4�+�4�)�4�4`��4F	�4*^�4zm�4�ѡ4�_�4��4�4�	�4H��4��4���4ބ�4Xb�4�	�4Zr�4�1�4�4�>�4�4���4V��4�4�4�V�4g|�4t^�43��4�4u��4�4f~�4p�}4�K�4�4*�4���41W�4�4�f�4���4)خ4�`�4BO�4^��4�l�4!�4�4�4Z�4�4̠4b)�4h�4r��435�4F#�4��4Ҙ�4S�49��4���4f��4�Q�4�!�4�N�4�`�4���4z�[4�T�4��s4F��4�̌4R�4���4q�4J/�3є�3���3�p3`��3O�3�O}3�/v3L��3���3jF�3D�3iV�3�x�3���3+�3��3��3���3�Q�3���3���3/��3D>�3f-�3�R�3J�3ܳ�3��3o��3�c�3���3�E�3Gl�3
4o3:�3��3 W�3��3���3���3���3F��3\x�3x��3Q0�3(��3�f�3q��3��3`L�3(��3)A�3��3���3(�3��3�~�3��3^#�3���3�o�3��J3j]�3l��3z�3�>�3�ڷ3��3_�3��3 ?�3�n3Z��3�@�3ce�3���3���3;R�3���3X@�3�<�3{��3V��3���3\��3�*�3k5�3���3r]m3��3͜�3��3}8�3K�3f��3`3�3:G�36��3��3��3a4�3�ka3P��3���3;�3o��3�N3���3+��3܇�3��3��3�Π3��3	�3�Q�3���2r��3��3N��3���3Ր�3��3L��3���3�u3���3���3���3�`�3��3`��3�g�3���3���3R��3�^�3�O�3'=�3x��3I)�3g��3�ԝ3m̺3�4�3��3&K�39y�3a��3�3L{�3H��3���3#��3r4�3ZH�3��1��3���3�+�3�d�3�Ε3�!�3��3X9�3��3�C�3�P�34[�3�3���3��|3"\�3%��3��3�{�3	�3.�3-%�3k��3���3K��3���3 �3zs�3���3�	�3@��3�Q�3f�3$K�3$K�3�E�3=X�3�`�3�Uw3�Y�3	g�3���3��3L��3c4�3��3 	�3�I�3��3��3�	�3��3���3�u�3?��3n�3���3Ddp3��p3�݈3.��3���3���3�>�3���3�3���3 k�3���3��3w9�3��3��:3���3�\�3S��3���3/�3���3^��3�gq3��3��3��3��3a[�3��3ID�3�3
��3*��3(��3���3�[3_c�3���3^��3w�3""�3��3���3!��37��3��3_��3��3�p�3s��3�f�3���3P��31u�3��3E�3���3���3Ii�3���3���3�<�3{�~3 0�3'��3qb�3�D�3���3V��3�^�3�a�3�n�3�ֻ3FZ�3֌�3���3�D�3B��3z��3���32W�3�_�3ߎ�3��3D�r3��3J��3���3�0�3Ȩ�3Ɛ�3�r�3��3�¶3�J�3� �3
B�3���3��k3b��3��3\�3���32�3M��3g5�3��3�H�3�E�3o��3�5�3���3D�3U��3�a�3C�3?�3��3�O�3��3�F�3���3��3wK�3̠�3q.�3-�3}t�3��3��33��36�3�0�3d�3�L�3��3?_�3��3��3��3�9�3���3k;�3��38q3��3h��3[��3��3��3���3��3��3�e�3���3�[�3ٙ�3�O�3 ~�3���37	�3̖�3qo�3p��3��3a��3Q�3��t3m��3��3ۉ�3���3�1�3���3]h�3C��3"c�3�B�3�^�3���3w��3�`�3x�3r��3_��3!��3���3�B�3���3�h�3��3Gx|3))�3N��3HM�3��3;m3�Yt3��3�3ҟ�3Ҵ�3�2�3(��3��3KB�3*��3ڑ�3H��3�F�3X��3`��3[�3��3|��39��3�b�3��3ۖ�34s�3ђ�3�;�3��3��3���3Xw3�]�3�{�3�$�3.�3(�3�m�3��3['�3
��3�S�3��3��3qj�3 "z3���2b��3�"�3���3l�3x]�3���3�d�3��3�]�3h��3(��3�g�3��3si�3W^�3EC�3_#�3���3�!�3i%�3�]�3L��3��3���3�;�3/��3Ye�3�3x^�3���3{Yx3R��3S�3R��3���3���3���3֓�3���3�<�3c��3t}�3L9�3�Y<4H�M40(K4�+4\�4*h94��4)�4�74�R@4s#>4�84��3qF94F;4�F4[�<4�l84)�4��74:p74�)#4T=4�Q=4��14 E64��4f�M4�<4 j>4�,44�>4�:54P�+4M<4�4J54�4n\L4�4��-4e�>4�=4�64��
4^E64�aE4��24N L4�..4C4�14��44�64��M4�N84�@4��:4=�)4"4��94�%>4SY14�T4~�54�/44V�N4��74	Y*4�u<4��!4&�.4޾4|=4��64�&4�|>4��/4a�4��4P�3�	/4�44F�4/�!4�/>464\"4R:4��"4<�84�94��M4K4A;4�:-4N4v?44��?4?4��04�E4�k?4�D-4�4�74v�14�54�4�3"574��?4d�B40��3��74<�94�4�n64��4N504�P�3*$;4�J45�J484wI4�pN4B =4�QJ4n�84��E4�*:4a�M4r�&4��M4��?4�?4�?4��64�.N4uIN4�<4�+84s#4�!4cM48i>4��M4��4V@4>4�a44��M4f4��:4:#4ǩ$4�d%4�@4Ê74� 84RM)4�84b4�G4�a64K4��4��:4
4�24�$4$V84�MF4o�M4��?4��94NM4�X�3ШM4�4˃;4�m?4�� 4e�=4
�4i�4Hh�3�'4a�34[>4�N4.*,4\N4�	L4|p74=�94,>@4#�K4-b@4�N4�n54�
;4�d@4�T4l:4��@4��4�/84�*4�84�y>4� G4p�84�J4u�3\�;4�=4��;4�M4��34(F4Z+4�a?4�PN4��94qH4�64�L<4u3(4�'I4��94�iM4�4<4�JN4:�@4,5�3�V@4��:4�04�>4c=4��L4$�>4�4�V=4�-4�>M47�?4�M4|B4��=4G�?4��4=�'4'�>4�A4-~?4J}?4I�?4$�?4�3+xK4i�>4�]94C�74�m4�;4�w94�F4�	74<�<4$b>47�B4�A?4��:4��)4� 4�N>4�gM4RP44�954!�84��?4A64�}?4-M@4S�.4��=4��54��64���3v�74�z+4��;4-�4)�L4i4�#4��	4�14�[#4��/4@;4-�N4�=4\�;4x[:4߈64��64F�M4r/4��64E<40�4 ]+4ˉ%4��M4��64�j4W�74�w4b4�*4[�54�64&�4�u4�l4�M4Q�4^ZI4�984�+74�T-4W4z�?4�2L4��74�*64�I4�Q&4��F4R�74�34��94!��3a�*4��84(�L4NM84
4�84�'<4vj?4Į<4fd84��74j@D4�w84��;4��M4�4��4�F4M;4�H14$b34��M4�<4d�/4�_L4��4�(4���3c34�;:4!�4A94ƝB4ڗ94�T84s;4A�N43HM4g�94�34_<4<9N4��;4ԅ4�4�Q;4o�54<w74�;4�@4f.4˯3�46*4��N4��;4@;4��(4c�3/k?4�j<4S�'401I4�94f>>4��-4�0.4�\74V~<4��*4��44�|?4�64X�4J4cn?4�?4	564��94�<4�TN4��!4h =4�EK4��?4�94�BM4=U4f?4t�(4ζ64�-4aH@4[4��M4H�'4M�4x] 45Q;4�zL4P]%4`G<4�@;4ß64�.N4��4�4��4k=4W�3 @4�X44l0*4�14�,84��F40,45�:4��3ɢ=4�>4�r;4D4�M4�I*4[N4�`�3"[4T��3�2N4��3M�?4�&14p�4P@M4Y�?4>�?4�m42"?4�/94��4NH�3��4�G4�]L4��'4Q4��34UN4�q64!n)4��@4�&-4φM4��5�545�|5!5}C5��4��5G5C��4v�5:�5��5;�50�53 5��58p5,�5��5PV5��5y�5۝5-�5��5�5`5��5י5�5a�5�45Y�5ؔ5,`5��	5�5�A595�H5�5S7�4��50�5EO5�r�4�w5��5�X5~�5�*5�`5�5d�5�A5�R5��5Y�5\t5ݻ	55 5�(�4?l5��5x(59M$5�n5��5�
50y5=]5�15?5�5�r5��5l5�5t�
5IG 5�L5ڤ5a�5��5t	5pz5A	5�5�Z5�v5I%55��5fA5�F5��	5/� 5z57k5�V5�5�/5��5R�5*5.5��5
�5�5h%�4�5q5�n 5
�5�5�,5.5�V5�i5��5��5:�5��5�5_�5Ы5K�5��5��
5k;5��56s5z65���4�)�4�_5��5�D54Z5 !5�5|��4q5R�5�V53�)5�
�4�H5��5�c5c�5��5J�5З�4�v5FJ�4�A5�5:�5�� 5��5�`
5�5��4�	 5�5^�5�Q5[P5VS5ˀ5cZ5�!5@G5�(5�m55�5R'5��5��42S
5Xg5p�5J
55��5z�5M5��"5�H	5�35��5��5M5��5��5��5��5�Y5��5��5��5ND5+�5��5\s5�5�5��5�5��5S5�45�5��	5�3 5���4���4��5�0	5�5-o5��5ڬ5�V5%�5��5��5_�5�5��5�h52�5�?5�	5 5�D5��5�5��5N85.:&5dY$5L�5�5�a5�05Pj�4��5h�5P�5�/5<5�r5�5��5�o5S5��5��5��5�5��505�{5ͳ5w5-�5;"!5�K"5¼5��5��5��5�V5�5�@	5'�5�5z�4�+5)�5�)5x�58�5�5�b5cv5���4�~5���4QM5�z 5El5J5�q5T�5�~�4�+5ј5��5�s5�5^�5W�5;�	5D�5�5�5�?5�_5�}5Ld5o
5UZ5�5�.5�X5�E	5�'5&z5�R5�5�
5n-�4b5��5@V5��
5�j5��5�k5�5IA5�}5#5Ǩ5X�5��5o�5�,5�#5a5u5ݐ5��57I5�Q5m�5�	5[�5ز%56�5��5��5��5;�5��53�5ԯ50�5{�5��5��5�H%5ڌ5�5�;5z�5��5�5r�5��5��4�Z5K�5�e51X5x5#C5@�5֪5�s5YJ5,05t5YM!5-5GI5�O5:5��5N5�U5�5O55�5�5yu5&�5��5f<5�۪4��5�5Ld5�5�5�4��5�}5��5�p5�E�4n"5�5c�5Ƭ5M�5�5��5G�
5�,
5a�5N� 5�5�5��5 �5yV5��5A5�95,�5"J5P�5��5H�5��5�
5�4#5~�5�5�5�.5y�5Nu5۶5El5�5�5O�5�5{m5,5�E5�5)��4f5,�5�5B(5A�5l5��5+7 5��5!j 5^�5�5H��4�85-6"5@75r�5�S5��5�5��5�?�4�u5 �5�5�5�B5�U5a�5v=5�w5;�5�
5�5s�50�5��5ID5	S5�95G=J4��>4�qC4�G@4�JW4k�X4p�V4YKX4�xH4��4~/A4�iM4TP4ϨW4�o4��F4�Y.4�?Q4eP4��"4��W4�W4�6O4��U4�YT4�R4�V4�T4�V46�T4�.@4@�=4�S4OUT4c�U4��H4�HT4�yT4�RL4�2R4{�44K�4X4Y�V4-PQ4)�T4�+W4߅;4��T4�yX4�m$4}�W4��S4��V44�X4�NX4-�D4�%X4��W4�ZX4j�N4˵$4�1�3��W4�5T4z�T4kX4�:F4g�R4��4�?T4Q4a�G4X�G4�W4��M4�3X4��T4}�H4W�W4�54�L4��:4ZO40V4��V4/�O4�cW4UkK4*�H4Q�<4�4��R4�3U46T4�E49oP4�34�2C4�_U4��K4��G4�W4� W4��B4��K4M�Q4��W4MK4߇T4�.46IX4qpG4�$T4-%T4��V4BOW4�H4�C4�W4F4��H4BcT4�4�@4�D4ƠR49uA4q�V4XR4�H4z@4�4W�*4w�04J�)4D�T4�U4�]X4ĔU4�O4.AU4k24ѽF4��D4��W4Ҧ4�)V44�T4܌E4GT4uX4s�T4T�V4L@V4l�S4�pG4�OT4�uU4��U4'-L4��R4R�T4)"O4K{W4U|X4�64;�K4ё24�NX4Z�!4 �A4 4X4EF04��U4X�T4�TX4)W4�WH42�T4[�4��W4~�N4�W4 fC4<�H4+�>4��H4RxG4�FW4X4��U4WDH4g�?4}�S4�G4+*X4��C4�ZV4�X4�Q4m14r}H4�<4*WH4m�H4��H4��V4�sP4��I4�G4zW4i0C4|�4��H4_"W4��T4��?4!�R4�?X4�	W4��G4��X4�V4�5W4O�S4��S4�=4�F4��4��3�:4-�X4�	<4�LW4��V4��B4�W4yP#4�%R4h�K4u*74dX49$4DQ4��U4+�T4ԦD4�X4tMW4�&4��4;V4U4�44��H42N46�:4��S4/hX4 ;S4�,)42e+4;X4%�U4�@<4vS4}oX4
wX4[�P4��4gW4��U4N\D4�pT4k�G4�P4|I4��H4�?4 �B4n�H4�Q4�PF4UW4�T4��G4��R4�vD4�8.4G�"4��V4�B'4T�R4+4XS4�F4�LW4i�R4�SU4�34�$V4YnX4s�4�Q4 /4kgU4:�14��P4{�%4�XH4w�V4�K4O,H4��T4�zX4�TK4�P4�YX4�_R4��H4TU4
mX4��F4��/4#tQ4�jX4�H4IX4��&4<�A4@4��/4�X4�S4"Z'4�X4�W46�E4`F4Ȁ4��X4�3S4�W4��?4y�L4��!4�U4�@S4�Q4ǸT4~G4��V4��F4�i>4�4gH4�lO4h2�3�%O4}2W4L94:�S4��H4e5F4J�H4��Q4n�W4�%W4w�V4	�P4_W4O�U4r�Q4ڵF4�164#�H44�4��H4m44:2X4�64��G4i�E4�G4%�N4p�N4aI43>U4��W4��Q4RGX4��B4�HT4ĐH4�%V4v�V4,*"4OM4�T4��O42<G4CS4ٓR4��V4��U4*�V4�H4�T4АV4B�,4�5K4ˮQ4
,F4
�P40�W4W1X4R&W4Y�U4��V4>�H4��64�~R4�8T4
�T4�S4�rX4�L4�4�J!4�?W49.U4e04��V4��W4֌W4��R4��U4��N4�Q4'pS48�H4?�Q4�@4�D4�V4*�Q4��"4��O4GcX4�7416X4�nQ4c�A4ޅL4.T4�x'4]xT4�U4Y�H4^�T4� 44�>X4�gW4�UX4�lF4��T4,T4A{B4M�C4% ?4H|M4PRH4�`;414�c#4��E4��S4�S4^�B4~~V4�R4�OD4��34��V4�7R4B�V49R4a&4R4�ME4� 4�f"4�!X4�DX4��G4Y�G4�H>4%V4}��3~�3o�3�o�3� �3��3�|�3���3��31e�3 g�3���3��3tf�3s�3�b�3#�3���3��3g��3�7�3�3�3���3���3�W�3A��3&�3��3���3Y�3���3%J�3���3���3���3ı�3���3���3��3���3��3��3���3���3�3��3"��3+�3���3-��3�k�3S��3b��3���39�3�"�3���3c�3 �3���3�
�3/7�3*�3:�3@��3���3���35�3�3�3F��3���3i��3$h�3k��3���3t�3 �3���3'��3��3�˿33��3���32,�3��3�r�3��3x�3��3��3���3}��3��3Z-�3��3��3&��33��3��3�^�3<��3�!�3��3G �3cj�3=��3���35U�3� �3��3��34�3�c�3��3<�3-��3V��3�o�3_��3�"�3a�3��3a��3��3X��3d�3i��3
��34��3�	�3�.�3E��3���3�r�3��3� �3��3Nq�3���3"��3�9�3F��3�3���3�`�3L�3 �3M��3J�3��3���32��3�g�3���3�K�3g��3U��3��3��3{t�3�3^W�3xy�3�{�3���3���3���3Y��3���3;�3��3H;�3���3���3���3��3�A�3��3E�3��3F��3���3ؽ�3��3w�3Zh�3H �3��3f��3[C�3���3-��3&��3	i�3g��3]��3���3<��3|��3�0�3��3]��3v��3���3���3V��3�3���3g��3V��3-��3�3NZ�3c��3���32�3�6�3���3��3��3��3��3�Y�3&
�3� �3g��3V �3I�3���3���3G��3G�3e��3̊�3�x�3wz�3Q��3$��3~
�3���3�=�3��3��3V��3���3f��3<'�3�3���3�3[k�3'D�3�F�3���3��3��3��3
��3~y�3c��3���3�C�3�3ʔ�3ZQ�3���3���3/��3���3H��3�G�3�3/n�3�j�3�!�3d��3G��3���3���3���3���32d�3r��3U��3	�38��3@�3���3��3���35��3���3zj�3��3j��3���3��35��3���3���3�~�3G��3��3��3���3��3���3��3qE�3W��3���3���3��3��3��3��3��3qt�3j>�3��3��34y�30	�3l��3���3;�3F�3G��3Mh�3��3��3'��3�3f��3*�3w��3���3��3���3^�3���3a]�3/��3���3H��3��3��3�!�3F��36�3uC�3q��3p��3y��3ZN�3���3,�3�	�3�r�3�3��3���3'��3��3(��3��30�33�3���3���3��3�n�3���3��3b��3$��3e��3zz�3��3���3��3��3�(�3��3�}�3x��3��3,��3��3���3͇�3ȉ�3�<�3��3d��3��3��3Q��3�2�3�]�3���3�P�3���3M��3��3� �3��3x��3x�3j��3��3���3���3&�3�M�3>�3/��3j��3%��3E��3�)�39��3�k�3���3)q�3���3��3��3`��3>1�3]�3�w�3+�3R��3޼�3`��35�3�$�3�U�3���3��3���3~��3P��3��3A
�3���3C�3B��3���3���3���3�3���3�3E��3yP�3��3���3g��3z��3B��3)��3�_�3���3���3���3+��3c��3�3�c�3H��3S��3���37:�3���3%�3���3.��3��3���3��3br�3���3�(�3���3Q��3��3���37$�3N�3��3r�3�3�	�3��3�3���3��3�|4o?w4tn}4�c�4��}4)�|42�46�w4��4]�w4x�4���4�!�4?�4m|4��|4���4}�w4:<z4��}4��}4�2�4Cŀ4%~4�m}4��w4s@}4���4��}4 }4��4a&}4t�45�}4J�r4��}4Vn4��^4E)�4��}4=B|4(�|4���4�Z{4N�|4u�z4��}4X�4�_}4�Q~4���4���4c��4E�}4ޞ�4ԛ}4I�4���4�ɀ4��{4U�u4�^}4�a�4�u�4��}4�|4��}4��}4�g{4Ct{4�i�4>р4�|4<�|4y�}4v�4�w}4��|4hK}44��4߉}4�k4M~4kc|4!(|4 o|4|�4�Q�4�%z4�-{4�΀4�y4��}4
O�4�*}4��}4���4<��4�Ȁ4�4�{4K��4ĭ�4��Q4||4[F}4vOh4a�{4�O4�}4z�}4��h4;�4��|413h4:��4!��49O4�o4�<�4�+~4��}4*��4��}4��}4a~4��|4:�|4!�}4�ʀ4\̀4d�}4���4���4I�4_�}4Q�{4��{4�y�4͎�4�}4_|4,at45�}4G3p4|s4g�4�X|4ᢀ47�w44d�l4�Xj4"8�4w�4_�4)	}42lx4n�{4"��4f>4�}44V4�iz4��4�N�4���4��|4�z�4ޱ}4�m}4FE�4�J�4I�U4�\y4�*�4�4ąy4�4�؀4�z4�E�4!�l4�	�4�
4\~4�H\4g�|4�}4�i[4�|4|��4/��4i?J4c�~4l�}4:��4Ծ4�d}4�X4�4cN|4h�}4�ŀ4!�}4��4�}4rw}4zc�4g�u4��|41Ā4�|4>�w4+�}4��{4�Tz4��{4T|4�(X4.W}4�{4�̀4/Q}4���4"z4���4��}4�k4mQ�4���4��4xm}4��4��z4��|4D�~48�{4��4��x4^��4�f�4#ŀ4�u}4�o4�h4hY}4fg�4�N{48@�4�r|4�3O4:|4�a}4l�|4D�x4��y4�6x4 ��4y��4�;}4�{4�k4��}4�4P}4֙�4R|}41 4$|4}4H}4�<|4��}4�p�4���4~x4�4�}4$4���4��4�}4�)�4�}~4�R}4{N{4�~4ۘ}4�׀4$Z4�v�4�h}4�u4���4��}4F�4��~40��4�74F��4\x4�{4�t}4Z|4��}4M~4��T4; }41g4�v4��4�l4�7}4Ҁ4<�~4�c}4�}4��|4�h�4K�}4�K�4�|�4ӻ�4�:�4�:]4AQ�4ԗS4uR4b=�4��}4n�n4]�}4{�}44z46]�43||4Ն|4�}4	�w4ϣu4Zh}4�v4-�}4���4�}4W�r4s�u4��4�d4b`{4"�~4��y4e$}4\}4b�|4�[�4ZT}4��z4	}4�9|4`n4�}4Ǖ}4m�}4��}4-�4��4���4S<z4E>x4�4X|4xx4�{4y��4Y4ax{4@p�4P3L4?}4C�4׍�4.�{4_��4m{�4��4w4��4Aр4�ML4ߩF4�b}4rGu4>�|4�n�4��4H�}4EK}4��z4~�o4a��4�y4��y4�H}4;�41}4q�}4��}4��|4��_4�ɀ4�w}4[~4�Wx4��z4�z4��4'�X4]ـ4~4���4��}4A�|4o�}4�A{4�~{4<��4�M}4*d�4&|w4��4A�y4&L4�%�4��{4ڮ|4��4!kJ4�1}4��~4���4�aZ4&�4�4y�{4��4�[�4�4��}4��z4�|4���4\ɀ4(��4`Ez4�2�4KZw4[�}4}4�~|46\w4cr}4��|4#/�4�<|4�}4 �}4)]�4��y4L~4j�z4ʞ�4���4�|4�JR4z�w4H�4Ѡ�4�j�4u~4ԃ{4�ڀ4 w4��|4��}4��}4bȀ4�Ȁ4���4޵u4[<y4ć�4pŀ4��{4�f�4�~4�Ā4%e4�U4�P&i��&��-&�S,&ė:&�<&�*&/�/&+??&�*�&���%�[&�o�&O�& �&�Í%@n,&̒4&�V&�Ɠ&��?&�o&'#Y&5�&�E]&ٔS&��1&��&�.�%;j&)�@&&�&�ܪ&��&��W&L_&��<&�0k&�.�&��&��[&�o&(�7&�+U&���%��P&���%���&s
P&#Ʉ&}��&Φ�%��&'&��
&_8�%�q&��&踍&��=&�bF&Q�%t<&��&�nf&��<&��&�[9&�'�&V?&�%B&'�$&b�V&��&���%#&}&%�*&��Y&��&c�2&���%��H&�~&�G�&��{&7[&�'&�FB&Dw@&=SX&��&\N�%AD&i�!&��8&F&8�N&��%%{@&��&�� &'�_&��P&ӈO&��O&X&�7/&�0&��*&o�,&y�%2�|&6	&&�&>�:&��+&)/&���&�'&C�&��i&׵7&��}&HO&��&��:&d�#&�T&��%�\&�)&b&!�z&5�<&� 6&O�&�C&R�&@�{&��&�-&oO_&��r&��%��$&�^i&:*&�,&8+&jk&�a&��&� &�q"&���%i�&�R6&j�d&�c&q%&�dV&�O3&U?&�#/&��;&��%�z&��&	{'&�+&{�&X��%�/&�TY&x�&s�W&v��&8"!&���&��;&��A&���%�&ȷ�&�}&��8&-}&�-&�&��&a}&�I`&�;�&�-&J�&��&��(&�P&�5&)�&
�3&1�h&��&�:&E�S&�bo&�R�&�]�&6�&V��%��>&���%B�:&D�&Hs&�8�%�:�%=i�&x�-&�T1&��`&Y&��(&�C;&��F&�zR&���%�8�&��}&A�&���&�:�&q9�&3�_&�@&��P&��&aD&��	&��&��&*cO&�&f4�%�L8&W<(&,%&��g&f��&a&Y	&��>&���&��&
�(&O�e&��P&�|F&�2`&���&��?&0�P&��&g �&��&&|�D&1��&�DC&���&Ӏ�&�&�
�%��&`&�!&�{W&�8&	&�&�_&��=&o&��9&��.&�L&`�p&�&T�2&�Z&�đ&�&��&��S&L�6&���&��@&�Yq&U�&9�&$�1&���%��%�!�&��%��;&�2�&ؗ�&$�&�&�*�%�&��<&y &�s&��S& �T&/�&2*&�7�%�A&��&a$&-�T&3+8&g�&�V&JE6&z�%��Q&9�)&k(P&�7H&7a/&�k)&8V0&w&�b&&)Jt&߉�&B\&�&bq&�nS&�s&��V&S7&?&$??&=2P&C]M&�B&||I&���&�*&��>&��%à�%�I&/ۙ&ٿ]&g>&;3&X�L&�b&�� &j��%�:&01w&�7&�&��%��&��h&[
q&8)/&�2U&4�*&�qU&EjS&�'r&څ3&{#+&:�&�]&�X&��S&&jSd&��&�bD&��&M�_&�tJ&�˦&q1&/1&��&��&�+.&�&�O&�[�&&P
&7o&#B&P8&q&�%&�j&fճ&.O&S�&@�&2�&�h&�gu&�6)&�T?&k7,&^�9&�/�% �#&��&4Æ&=D#&F��&���&��[&��&��:&�h&|ވ&�}&�$&�0&��|&\[&�;&�Y+&��:&��6&,U&��&��9&��;&�lZ&��Q&�*&53&+�E&(~�&�&9��&:�i&&N&�|K&^�&
H&�n�&{�,&�!&uU-&�O&�Ο&a��%z?&~�N&_#K&z�&{�F&j�C&z��&}��%��K&k�$&<Ԉ&[�'&��&|��%ӣ2&��,&�>!&n�[&x�%& F3&��'&�2&�Z�&�I&�?X&GG�%5-&�aS&�&��&��*&�V]&�)F&;��3t=�3�L�36g�3�H�3���3n��30��3�9�3=,�3���3K�3�Y�31$�3��3�,�3�3^��3�9�3>��3�(�3d#�3�/�3+@�3?��3�<�3���3�j�3]��3���3S�3�m�3�G�3�4�3x�3��3i��3�.�3B��3KZ�3�}�3��3W�3�,�3
�3�2�3a1�3_��3:�3��3
3�3k"�3J(�3X��3��3k*�3i��3�P�3�3�z�3�m�3C�3��3pA�3Fe�3��3�5�3r��3��3� �3?��3 E�3�k�3I��3y��3��3*��3�Q�3]��3�(�3);�3-��31��3��3!�3/��3R��3I9�3���3��3��3���3��3�8�3���3�C�38�3���3�?�31 �3�	�3MB�3���3�(�3[a�3��3�)�32�39��3��3�0�3���3
�3��3�	�3�C�3�#�3���3���3oE�3�:�3y��3$F�3J�3W�3���3u;�3��3x]�3$�3��3��3|�31�3�3�3)��3P��3r�3XN�3?��3�i�3��3lY�3˧�3���3x��3.W�3���3��3*=�3��3�K�3�H�3f�32[�3n"�3�1�3#�3��3'�3R�3���3L �3�:�3��3��3�6�3�N�3��3��3��3l@�346�3���3���3��3�:�3�a�3�G�3�o�3A8�3��3�^�3��3�L�3-[�3L�3/�3�'�3f��3ޏ�3��3�i�3���3��3n��3��3��3n+�3�g�3���3�L�3O��3��3J�3�y�3���3i��3��3�9�3+#�3��3x'�3��3C�3���3|[�3M��3�Q�3V�3���3w4�3�7�3  �3C�3Ch�3�C�3���3���3g��31�30��3/�3�e�3�)�3A�3R'�3$�3�$�3���3d+�3�6�3.?�3�Z�3���3���3\$�3���3Y��3�K�3� �3�o�3���3���3&�3�u�3��3�X�3��3 ��3�I�3�3XV�3@��3"��3bN�3
��3�f�3`��3���3l��31�3���3�'�3�-�33�3^S�3�+�3�3&��3��3R-�3���3���3���3ӳ�3�3��31�32�3��3L7�3	��3���3���3���35,�3@��3��3l=�3���3CJ�3�3���1Q7�3�P�3��3*7�3�3�3t�3E,�3$J�3�p�3ٛ�36�3�v�3B��3���3�D�3��3�3,�3��3�3���3("�3�@�3n#�3g��3�J�3uK�3�/�3e�3��36I�3.�3���35�3���30�38�3��3���33A�3���3���3)�3�y�3��3�Q�3c�3�#�3i��3\�3%�3���3-��35��3�;�3�2�3�9�3��3���3���3�Q�3?��3�2�3�)�3�6�3���3��3;�3!�3���3���3[�3���3k��3���3��3f��3�"�3jL�3�<�3@=�3c��3�3�+�3��3fW�37	�3+�3;�3�0�3�]�3i+�3%��3���3v2�3���3��3Ti�3�2�3�(�3D+�3=��3��3�"�3�Y�3$@�3���3@��3��3Gr�3���3�2�3� �3���3��3Uk�3c�3��3��3�|�3u5�3l6�3h�3@�3l�3�'�3�2�3���3�3�1�3��3�B�3J�3��3>��3���3��3���3r��3� �3x��3j��3�D�3t��3���3��3��3��3�0�3OW�3/��3-��32�3d��3P�3��3!�3��3���3�b�3BL�3���37�3D�3�
�3�d�3���38�3�Y�35��3�J�3���3�U�3)J�3ɍ�3v�3.��3���3���3|��3�3[�3#�3H��3���3�t�3E%�3�5�37�3�h�3�2�3���3���3ރ�3��4�t�4+��4���4��4��4���4k�4���4Rj�4���44��4��4۶�4���4=��4��4w��4���4�>�4l�4���4�S�4���4җ�4��4���4���4I��4���4m��4���4��4F{�4���4��4���4��4D��4g��42�4�/�4,��4�4C��4��4���4<$�4R��4�G�4R��4 _�4�_�40 �4��4�
�4Z$�4�<�4�^�4���4f�4l_�4�˽4���43��4�~�4�4���4M�4�u�4`��4�k�4�G�4���4mq�4E�4a�4��4a��4W�4���4�z�4��4�3�4�\�4Uh�4/�4�@�4��42>�4�o�4���4I6�4��4P��4i�4.ر4���4$0�4Q'�4���4�u�4�=�4_;�4@��4�W�4&�4)��48"�4q|�4��4?�4T_�4vA�4�4���4F��4���4A��4��42��4x��4���4#L�4���4���4��4���4(��43)�4���4���4�ݲ4K3�4�#�4r2�4���4��4XI�4�>�4���4
��4]O�4�i�4�d�4���40޴4I��4�*�4���4ٹ�4��4���4�W�49�4#��4;�4X�4KV�4�R�4��4m��4�4��4���4S*�4���4n�4+��4��4Ԛ4�J�4}*�4J��4>��4/�4r^�4�%�4��4Mq�4�/�4�/�4}�4E��4�%�4ͨ�4H��4���4]��4<��4��4�|�4C2�4J��4���4�!�4�3�4�4E�4Sl�4H��4���4S��45�4��4���4e
�4���4�ի4с�4�&�4���4���4�$�4I��4mz�4�B�4���4l��43�4�_�4Rs�4�a�4a��4e5�4�4Z��4���4���4D��4�4�п4\ʫ4,X�4o��4���4�4���4�7�4���4�n�4��4���4?��4QR�4�k�4�,�4Ϫ�4���4���4�߹44�4(��4�-�4��4�=�4w��4��4��4�(�4�4��4��4)g�4r;�4/��4?p�4d��4v��4�]�4��4��4?v�4���4��4A��4%��4��4K��4cY�4�v�4��4�L�4�k�4Y��4I��4z��4�`�4���4�>�4�h�4��4{�4���4<�4��4���4���4���4���44��4�`�4s�4�8�4�3���4���4��4 ��4 �4���4�v�4y��4Rd�4���4���4I��4S=�4��4d�48��4�	�4���4HC�4%�4��4NR�4�r�4\`�4 ��4�`�4���4z��4�Y�4���4#�4'��4pñ4��4��4+׉4���4�>�4�e�4k}�4��4k��4	�41�4���4���4���4��4Q�4O��4�ѻ4	/�4��4�z�4��4E��4'D�4��4��4j��4�V�4�S�4���4�4��4!��4���4���4M��4�4��4}5�4��4���4Y4�4d	�4m��4���4>��4	]�4�U�4U�4�O�4��4z��4��4��4���4z�4���4V�4e��4���4U��4��4\��4*V�4�N�4?�4j�4�j�4�s�4�k�4�U�4���4��4�[�4S��4�^�4PK�4��4F��4!�4˥�4��4K�4SA�4k]�4���4`��4���4�+�4�4	'�4LW�4���4�B�4�}�4�,�4�d�4��4���4{�4�P�4v�4c�4���4�"�4��4��4���4a��4|}�44��47��4	2�4���4�,�4���4���46[�4�L�4�-�45��4;��4�&�4�t�4���4���4g��4�4B��4aU�4d��4��4���4��45K�4�?�4H��4=�4��4!��4�d�4/O�4.4�4��4��4���4\��4��4^[�4���4��46��4R�4��4B �4=~�4�C�4GB�4CE�4��4�P�43��4@��3�3q4�/q4��q4�xn4i�e4E3f4\54�Ag4h�3��f4nq4�g4��f4�
f4��p4�q49r4�cp4�q4޾q4Q�p4lr4��q4�og4��e4��q4�Lr4��A4��j4D�e4E�p4�q4�<n4	�-4�c4��c4'��33f4C r4"r4{>e4��f4_�p4EMq4��n4��f4��f42r4�r4
q4�r4:n�3\cq4�Y4��g4�ar4�q4��k4jdr4PLp4�r4v�m4g4��q4C�f4g4!_g4C}p4lq4�g4}�q4Ώ4��d4�f4rr49�q4(�n4��q4�Bq4�fg4��c4"+r4�$p4�+q4��f4ʑA4�q4���3��q4*e4�q4-}g40g4��p4�r4 S	4�b4�p4Iq4V�p4�bg4O��3��l4�o4�q4�lr4�rg4�e4]�q4!Wg4��q4�`f4�q4�e4lg4&�p4��d4��e4��q4U&p4z�`4Gr4-[p4+�q4��f4:��3��f4�f4��q4�g4Q�34̢`4�r4z`q4��f4Y�q4
sF4��q4�G4og4�sq4~jm457p4ԟq4�Lf4��e4W�o4�r4��d4J\4|�m47r4��l4��l4�T4Uyi4z:e4��m4�sr4Hg4��q4��d4��e4�e4�-r4�f4ǋn4��q4�wg4��4�q4�r4ǰq4&f4��p4G&g4�Mp4��q4�(�3�6g4�\q4��i4%�p4F�f4�f4d�p4�7o4��f4hEc4$R4��_4 �q4�sg4��p4W[e4��q4��P4O1o4ur4�Bq4��g4�5f4r4NIo4Qr4�An4��q4�34�Yo4e�q4��d4,Xg4�a4Gg45wp4��m4��n4��q48r4�np4O�p4��q4/eq4��d4�i49RZ4��p4�Vp4�r4r4Uj4`��3��q4ôe4^Id4%Tp4��p4mZg4,e4��q4�gq4]@r42lf4��g4ul4��f4v�o4u>^4�\g4V�e4ZXp4��p4MCe4�r4��3�k4��l4�-g42�q4�,n4u5q4.�f4��q4�c�3ѐ�3��q4�g4 Yf4�m4�b4�wf4[�f4�(q4Xq4�ar4�/q48|o4�-g4�~q41?g4u�q4i�o4�pd4�q4ٯq4��p4�`4�.�3"r4>�e4Pr4��p4k�`4D�q4W�q4�o4qer47�q4�q4��q4 �q4<�q4N�e4���3��q4�)r4�l4:14Ye4-�q4׽m4� i45�G4��q4qqp4Oe4�>r4,g4|�f4~��3
�p4"Ip4C�q4;�74�Ho4��r4rsq48�q4o�q4Up4��h4er46r4�#p4)�f4\�p4�-	4��g4A�c4}c�3�jj4l#r4��p4,/p41r4��q4�Za4��q4�`o4��p4��p4{7p4K�o4Zn44Kg4��l4q�q4�M4��q4/�q4�^4B�f4�q4n�q44�q4�o4��f4hJg4,6p46�o4Xc4�sd4�s�3�B�3;m`4��q4Oq4�r4�r4��f4c�i4��q4�=q4?�q4�q4�Zg4��d4&q4wWr4��i4�G^42q4Q;k4�Vb4͎q4c&r4��m4�(r4N~p4n�p43q4Cfo4�n4��f4��?4;r4�0g4��n4R3f4|\g4��o4��q4b�f4�`r4�Yp4�Nf4��q4�\4x-g4��e4�r4TSr4�~f4��q4r�q4��p4]�q4|ve4�&�3Te4)�q4C9o4]1d4s�p4�Wp4��q4��g4�Wo4�q4��p4�+r4� r4�q4E�q4�d4.g4	0r4�q4�0c4If4?kq4Ag4l�l4Tr4�q4��3��n4��q4�7d4�q4�a4Wg4�q4�Sf4��n4�9g4��o4�Vq4&p4�!q44�p4��d4R�q4��q4:_4�Up4�Nr4sf4��q4Y�q4�g4g�q4PeQ45r46k4�6r4@�f4�6r4�Dp4:�n47fp4FFf4 �q4��f4�q4Uf4{�k4��p4��q4{�5ڈ5Ơ'5�(-5��,5�#5|�5RT-5�!5�f5�� 5�G"5NE!5�'5�y5?�5.�%5i�5 r,5y#5�-5� 5�:5��,5�5��$5:} 5�"5�-5yR&5�M 5��%5�A&5�$5u�,5�5��*5�$5f�&5��5=0!5��5��#5��$5e�5�$5�+5n�5�$5�C-5�s5~m&5��&5K�'5�'5�n 5 "5B''5��%5��,5�#5�M5C�5�" 53L$5��5�h-5�5O�!5.E5#5��,5��5�"5�g 5�#5�3'5"5�1!5��-5�c5�25V 5��5W�,5�f%5P'5�'5��50"5��%5��5�5�� 5i�+5�E!5I�,5��5(!5��5�*5_�5�59Q-5l�5�^#5#�5��#5��*5J$53'$5�$55g#5��#5Q8%5�V'5�M-5Y�5�r5E�$5p�!5�05��#5ˬ5.Y-5��5�b#5 '5�� 5�X+5o�5�8 5og!5�"5v�5�>5#5T�&5VF)5U�,5�$!5�[5�Q5��5�m!5*6&5>l5#i5?H,5n5˝-5a-5q'5U�"5��&5	�5��#5�;+5�5C'5��5: !5a�,5� 5�,5��#5b�,5 5(Z"5m� 57D'5�&5�&5�-5O-5*�&5��"56�"5�!5��#5��"5�q&5�25-5�R5�5�65	b$5��5�� 5.x5C�,5��"5��5]q5�w"52v-5Tn"5��$5r�-5�s5Q5О5�h%5T�#5i�5#�5�T-5�O!55�!5b�!5�-5�5/5J5�)5.�)57�5G!5ޔ-5��&5��"5�5+5M 5cM$5>&*5-�5�
5O' 5}�!5w�5�e&5ci 5��5C5�\-5��5X�&5�}5Ԛ5t�+5V9(5�:'5�@'5l &5,5 M#5i� 55��&5yg$5 � 5�o"5\�5�-5w� 5Y�5�5��5��&5(�!5��+5g$5�v-5H�#5�V5�� 5
$$5��,5��*5/� 5K5o;5�p!5W!5�a!5��"5�j5\	5{55�E$5�C"5��5xi,5�5K� 5�"5 e5@�,5"�5�l&5��,5��5�J5 $5z 5�$'5r<$5h�%5��!5��!5{d-5.5���4�$5��,55K�565!M5m�&5��5.�"5;('5��&5>�$5$�5g�#5��&5�=5-B5E.-5d�5J#$5e5�'5}�#5�|-5�#5�75�.5��5��%5cI5J�5x�#5�h-5�#5�I!5Fz5��$5P$5��5�5y�#5�d5��#5ɦ)5�)5�n&5�� 5	k-5�C 5H�5�#5]�5=-5�P5�k)5� 5�5��#5��5!�!5� 5V5�p5~'5A�#5i!5Y
&5�X)5+~!5�!$5�r5]=#5�Y5��5/K5�#5X&5c%5"Y5֡"5Ȩ5"5��5V?#5��&5��5]5!5ޙ#5�'5��#5��!5�*#5l�&5��5X� 5b9+5;�5�5P)5��&5��&5�9-5Z�5��5+�#5[�,5j!5��5�q!5�'5�k$5�-58'5�05{}-5�9 5�L$5,$5�5�%5��5Y�5/,'5��(5��5��5�-5Z5;v5<k,5�<%5}�5&5Vm#5�z5?#5��"5G�#5��!5jN+5�#5zu5� $5u�5Z�5�#5`�5`'5�45m�+5i�$5w�"5�5k!5U�"5��5a~)5A85�q 5��!5�<-5�$5��*5}!5�x5 35zV5C)50�!5g5 5�"5� 5�5��&50-5�5p�&5�!5�4(5 $5S'5��!5�,5�~#5��5�(5f"5��5�,(5�"5A�-5�"5�� 5�%5[�%5S�:'޲W'��
'ݢ�&�N'MuW'�ID'*�E'bT&�O�&m'G�%'��&�Y'H3'�A'#�J'��H'WH'P�0'8s^'��-'�E-'�)^'$�`'3PC'!�8'�=�&?�O'R�q&'�b'PD?'�T6'��$'ƈ;'Z�G'��'9'�#''�M'^PM'uLD'-�T'�<'�O'˨�&,�I'�P'^V'P�P'K@a'��@'��X&[ZP'Q^>'18J'�2Q'==U'Md^'! X'vVC'��L'�K'�@'.VC'��@'8''�Q'��1'�QL's^W'��E'�S'h�F'�pK'J�M'��'���&�UR'B"e'��S'�8'^XP'/�'��`'�aF'�kG'�'ڌ�&6�L'�yJ'�C'�8H'��M'�P'j�N'T:'�Ɍ&�7'��D'd'�DF'#Q'N_b&M�F'���&љ''�#'R�7'�AD'�;u&��@'^�&=�^'�3+'E�S'�<G'�L('�a'.LH'~<M'��Y'�	R'��'H�5'�H'<+'].E'��!'`)5'��Q'�B'�e1'�`'6K'8'`;2'�4H&En�&�NZ'
�U'��&I�'�]9'���&��A'_>\'�'&֙M'�j�&��W'i�>'(q'��&5�I'b:'��R'�&@'x�c'��/'�_&	J'&�E'$\P'��.'0�"'^�<'Q�Z&�wl'�T'}	L'4BV'�8Z'g�J']~N'��6'?'���&�t�&1Q'TV>'��6'��['�e;']�&��W'dF'��U'�8F'2��&�S�&�Q'2E'��d' @'�~`'��-'�C'�$-'u+'6�&��&��'�{?'pSG'|C'��`'��G'��('L��&�I'4�F'��F'��\'~gS'�X'��R'[��&��D'�SS'���&''<'hz('ќK'n'O'�Y?&�u)'��8'��'�-\'�)�&�@N'�D&kǾ&��&�d&cI'�#c'��M'��:''~''@B'F�H'saD'V�.'�~9&��'mI1'$�I'��T'��J'~�M'���&aj'��1'hJ�&�JI'tJ'PH'��M'��N'=�X'�\'�3'�L'��H'�_M'҆�&�"k'��&�JA' �o'��0'	�0'�R�&�bY&� M'�LY'}�B&��5'#�2'��J'W[{%�'y��&��!'�X'��M'�M'7S'V�H'��&��W'~�7'�G'�S'ԥ#'~8='%.'b'u,�&1�'�" '�\\'��c'��&�%'ZZ'G�"'�w�&��$'�[�&�-'A�)'X9'?;�&(!2'�)B'�FG'�I'y&�h;'4�H'aD'7(['�t3'��'
Q'�cK'rHJ'`;E'G�M'/�'�ƛ&�Y'N�('�@'Z�&�G'�z]'�lW'�H'�"@'j�G'l#g&�(�&��&V'8'�MQ'�'*�0'T9'�C'B"h'�-'��'��?'���&�(7'�f'-c'���&���&��='!V'A.�&LrC'�'�T'\=P'�kO'�IE'ղd'>HY'JL'&
0'p�Y'GJM'�6'�)M'QZ^'��W'�0'Q�`'~�&��E'��&� T'uY@'H'�PI'��&��O'=RP't\'�$'8�/'��A'-�n&�L�&w8G'h�"'��c' �L'|�H':�N'F�G'+``&υ�%��K'�^1'oN'��T'W^'Q�?'�W'5'-�:'�3"'�<�&�N�&	J'߿�&�L1'�qZ'�>B'�3i&�X�&G��&��'q�E'�!1'�5'$I'�1('��0'��A',�s&5�O'F8R'G�%��B'�(�&`+L'KL�&�!Y'W X&z�I'�L8'��H'��5'T�0''�T'+@V'��&��R'�
T'��&�)J'\�F'�H'*�R'� �& 5M'��8'�:'�)F'�SD'��E&K9B'U�G'fZ&��^'2�I'�I'�3.'m�'H�>&1[�&��z&&n:'�'4''8fQ'�2'e߆&�U'�HB'�'P'j\9'��Y&0�<'�E'��&��V'�=W'��C'x�f'�Y'��3��3,{�3���3���3M��3�3s�3H��36��3���3=s�3V��3���3���3���3���3�j�3���3׏�3a��3/��3���3��3p�3���3� �3���3)��3M�3D��3X{�3���3�~�3�?�3���3//�3W)�3�T�3��3[�3��3���3dB�3�g�3)��3؝�3�3���39�3VU�3���3���3��3�m�3��3M��3�`�3��3��3�c�3���3ֲ�3���3;��3�Z�3�F�3�p�3 ��3��3��3���3Us�3���3G��3p��3p��3���3�y�3x�39��3�`�3���3�`�3��3�r�3���3P��3F��39��3���3�g�3�0�3�j�3��3���3lv�3aH�3�w�3?3�3R��3�:�3!��3jG�3M��3��3�n�3w6�3��3_��3`��3J�3���3��3��3֔�3H��3`1�3���3�i�3���3܆�3�K�3 z�3.`�3?Q�3Z��3~M�3�S�3�$�3Ή�3\��3փ�3�l�3} �3�}�3?��3�=�32�3�!�3�z�3��3O��3��3�L�3d��3z��3���3.n�3��3$<�3�o�3�9�3.��3��3���3�e�3nv�3���3��3��3A��3��3	��3q�3�H�3,q�3�{�3|p�3ك�3���3<$�3���3rP�3�{�3�[�3�>�3:��3N$�3���3���3�E�3�3ZI�34��3b��3U��3Ʉ�3ǌ�3��3���3�K�3�i�3�k�3���3��3���3�l�3�`�3���3���3{��3�:�3��3k�3�d�3���3$��3�J�3�|�3-|�3���3��3��3�{�3�=�3P��3���3�V�3-��37�3�D�3���3��3P��3���3���36��3��3��3���3�m�3���3cm�3%	�3S�3'�3lf�3�}�3x�3FF�3���3�3w��3��3�3�3|}�3e��32��3EY�3��3��3E��3���32w�3�3�3���3(��3�Z�3D�3JK�3^!�3\��3���3<�3��3�p�3%}�3�|�3Y�3�p�3���3���3l�3���3��3��3}d�3�8�3a��3W��38��3\��3[K�3]W�3�|�3	!�3q��3~s�3�g�3�<�3�C�3Ǐ�3)��3�&�3�v�35h�3���3Pj�3g�3~�3��3�|�3���3��3�:�3w��3J�3K��3\��3�_�32M�3Y��3d>�3���3^�3��3��3���3>��3��3(��38��3���3b�3��3X��3Ø�3zh�3��3"��3!�3_�3ɒ�3��3<��3��3Y�3�3�B�3���3�z�3\��3�L�35\�3��3�]�3d�3��3��3���3E��3T}�3X��3��3���3^L�3��3`��3n��3.��3��36�3���3���3ku�3f�3���3L��3K�3�H�3s:�3y�3��3���3mx�3U�3�}�3�3ߜ�3���3�4�3�3���3���3���3h��3f�3�X�3#��3�Y�3]�3��3A��3���3`G�3>��3���3�d�3,��3���3}�3���3\��3T�3��3���3��3�W�3�3$B�3�9�3���3nN�33��3���3��3�h�3�K�3�f�3?v�3a��3�Y�3���3O`�3���3�3�3j��3NT�3GC�30��3��3Y �3^o�3V�3�R�3�h�3R��3���3\��3�"�3���3g��3{o�3�6�3�e�3���3|q�3���3��3l*�31y�3�r�3P��3�w�3&}�3��3���3�0�3j��3"J�3�J�3���3*.�3G��3���3�$�3->�3�H�3
x�3Μ�3���3�F�3M�3`�3D��3�_�3��3�p�3�>�3q��3݁�3!��3O��3[�3@��3�T�3lv�3A��3@H�3���3h��3G��3���3O��3.��3��3��3)_�3\�3 !i/��9.>�G/.g/�}�.5H/��b/��/��0/�[/=%i/�=/���.�I/rT/W�-/t,/5c/X /QQ/�m/�za/�Q/�E/��U/�X/:MH/+�m/_?/��5/i�G/�7�.-:/��j.��N/��V.G>/%_/Sl/s�B/'�\/T~�-tm\/݉.�A/c�`/X/xYX/�Un/���.k�M/��>/޳N/��[/��k/@=[/Ai/�X/8CX/�s/{<k/g`n/f6d/Q,7/UWq/�5/� X/�qY/��l/Z]&.��d/"�W/q�U/�ab/i�a/���.�F/ᆱ.Jj/~�U/A�m/{3�.��.Wmb/{�b/(ݵ.��.��[/��a/�?P/Z7X/7�\/q�s/�\&/�P`/��f/A�/z>E/��V/�i/o��.��(.�m/t�P/,4^/��i/�`U/�U%.�{_/[O/0�"/9i/��R/q�-?�.��.��n/�W/�m/a�5/��_/�;Y/}��.��8/ٌ%/�N/�zo/�b/f�Z/��A/cq/��f/�.���.��]/�=*.�E/B�U/�X/y�`/gi/g�.�EJ/Ts/l[U/�gk/[�X/U^/$�/K��.PX/l�D.��]/�9^/ӱF/\�R/�xe/b�f/��U/��.Ηd/��M/�b.�/H/x�!/߸/��]/|�(/8k3/B�`/ֹ[/H�2/�G�.ҘW/��e/���-�v]/dg/Ph_/TQk/�o"/��6/p�i/�T/�Q/}b;/J�d/��[/�7W.�
a/ҝ</�	`/��U/Q,/�ut.}t;.�lv.y�l/�al/��d/�`/���.�<9/l��.�"�.��B/��T.XD/�YS/C�S/�$</�]/�B/h�g/g{l/7PO/nm/�ӡ-�Q/��M/��i-�v.��^/ʽg/w�T/�gZ/-k/��C/U�.�HV/'�.��`/4yT/�Ua/�Jc/�~3.��`/9�P/>OU/�+H/U!/�Q/�C/gq/�c/��T/�d/�b/,�I/֕4/�d/�^/Ka/k�q/]�D/[_?/9�b/�M/څ6/��/S�H/��q/��d/��j/cV\/��X/Nb]/ǺR/�&`/�3^/��_/��L/
#i/�m/@�:/��M/��/Q8�.=I�.�?q/��.��_/��X/�<G/��n/JJi/}(/�W/oZ/f�l/���.C�a/�s/�X/-Vj/�FH/LOU/��\/�X]/�aW/ֈ`/�(]/#X/u�;/Ơ_/��j/�gW/§L/��h/��b/�v@/��Y/.8Y/.`/�S�.�tS/��.�Ԓ.A�M/R�5.��l/��/ 3l/�ݒ.�aE/d�e/�i/X:`/�%e.Q�f/H�/��f/W�[/ܔU/���.��Q/'�l/�pY/8�a/B~�.�EW/�`.]�]/��U/�p�.��8/d�'/��R/�Z/��f/��K//�L/��Y/��./�Y/q�#/;3W/��h/}��.J�N/Խg/��[/�0[/*U/�~h/4�e/��Z/B�_/h�d/��d/-<.>�R/c1U/ڄ6/��Y/~��.�bf/G(9/�L\/�x/Q9M/�
%/�a,/ʶp/ư\/��^/fj�.�� /e.IWa/2�\/a�S/�a/�6c/v�^/�a/��t.��a/ΙI/�.j4Y/m�n/\�f/I#."�]/��.n� /���.��@/�?^/a�P/��a/�[.��I/k�Q/J#k/��Z/u�^/�*.ηf/�]/ �n/I�/��A/P��.�bj/&�b/�E</�X.|��.��L.[�E/UjT/dMJ/J�l/*�k/��:/�(V/���.��^/�T/��N/��X/Sh/$�N/�=^/�7E/R|>/�mf/�+/�?U/��.�'B.bF/^H/�Q_/��c/]V/6[/�7/Rjc/��U/d�5/��I/#�D/�Δ.�?T/�,]/��d. /9Cb/I�@/R /�_/Hue/&W3/�r5/vq/g�h/&x/�+S/'c/S� /'N/�[/�=/nV/Th#/�O/�J/ߊ^/R�O/��m/z�U/G?/��^/�q/��k/�#(/��4}��4ef�4^Ȋ4ia�4�j�4��4��4ӻ�4�A�40�4�4#8�4�Њ4و4̵�4ڊ4��4 Њ4a�4s��4�4,b�4h�4���4��49��4W�4���4�P�4g��4K��49��4V��4�j�4��4�f�4د�4�d�4�э4���46��49��4J/�4Բ�4�l�4[��49��4���4���4��4܉4���4���4���4H�4��4�4�֊4,�4��4�׊4y=�4���4��4@K�4�׊4���4.�4���4��4��4+I�4�l�4d��4K̅4_Պ4��4YA�4��4��4V}�4�1�4��4cx�4�)�4Ge�40o�4�Ћ4)�4W��4���4�Ս4r�4�[�4��4��4z��40�4�4�4.č4���4��4*ԉ4��4��4Ս4��4E��4m�4섊4:k�4{F�4�8�4��4�4K�4��4��4��4]ԍ4c��4�4d��4�4ۖ�4�E�4܍4QƊ4"��4b��4Uӊ4���4�ۊ4U�4��4�Պ4}��4ӊ4̑�4ԍ�4�҇4��4R}�4V�4F�4Z��4͊4U�4���4��4��4�2�4Ux�4�&�4l�4=��4ő�4��4K��4X�4�`�4���4���4ȍ4�Ȋ4��4���4�ލ4-�4r�4���4���49̊4֣�4��4l9�4�|�4��4�z�4���4�x�4b��4(��49�4ah�4/��4쪍4�ԍ4 �4?��4���4��4���4uǉ4̊4]c�4�4� �4i}�47��4$�4о�4�T�4Q��4
�4nʊ4���4���4��4~��4���4���4���4��4� �4j��4�]�4��4�Ί4X7�4�4f��45΍4�/�4[U�4�5�4 U�4���4娊4��4Ԩ�4��4��4�ߊ4�R�4LĊ4��4fό4��4ۼ�4��4��4�4Zz�4�K�4HT�4�׍4���4um�4>�4U�4�)�4Qۊ4�[�4͂�4�V�4���4͊4��4)L�4��4��4��4��4	��4�}�4���4"Ĉ4�ۍ4u�4e��4��4�ݍ4g�4C͈4c��4��4Ҥ�4 ��4���4�ˉ4�4�r�4�9�4FC�42Ή4���4���45ɍ4�b�4��4�{�4Q��4.��4�4�4Ɗ4 ��4�=�4�Ҋ4�͉4�Ê4�4Զ�3 ��4�Ŋ4���4N��4��4:��4�r�4���4痈4	ފ4ଊ4pډ42*�4�y�4�a�4�4 ��4�Ԋ4S֊4"Ċ4l[�4�ˊ4��4��4q��4$��4<��4���4^Њ4튈4zߌ4��4�̊4ӷ�4���4%�4���4���4�q�4RÉ4X�4��4�ވ4#��4��4���4~V�4��4!�4�4�4���4�I�4�_�4�4,��4o�4�È4�C�4Ժ�4���4/�4���4��4��4�ƍ4���4�.�4�Ɔ4FU�4���4�Պ4jԈ4���4b��4��4�e�4�.�4��4¾�4��4'Ԋ4L��4l&�4���4��4Ύ�4�h�4���4r�g4*�4���4��4d�4�Ɗ4��4�l�4@��4�=�4љ�4Z��4bۊ4+��4�3�4�c�4跊4��4��4�Ȋ4}��4��4��4㱊4Nӊ4��4>��4�K�4�4�ۊ4ݨ�4���4�e�44`�4Fۊ4)��4�ډ4|��4��4զ�4[��4��4s�4z��4l�4]Ӎ4��4��4�ǈ4��4�u�4	Ɋ4h��4�}�4���4��4:ˌ4�8�4;s�4�׊4HЌ4`4p�4�È4��4��4 �4dl�4dZ�4rތ4��4�y�4Ef�4�ƍ4�2�4Ά�4>X�4�Q�4͉4bC�4+��4�Ȋ4���4� �4 ފ4�42ߊ4�H�4s֊45��40�4b��4�Ê4�Պ4���4*Պ4n.�4���4��4C��4*�4�
�4�4Uڍ4ڶ�4�D�4�5�4��E4$ME4a/G4�F4�4G4,:G4{�F4CG4|2G46A4��F4�G4�@F4ӟF4:AG4��F4GG4G4�+G4aIG48mF4�FG4(+G4z�F4�G4�}D4ĺF44G4s:G42�F4�zE4�G4�uE4o"G4�F4�G4,B4��F42�E4�*G4x�F4�\F4��F4��F4_G4�?G46G4e�F4�>G4"�F4��F4�F4�#G4�;G4zG4�CG4�BG4��F4^3G4@G4R�F4�8G4�aF4w(F4<+G4W�F4'�F4G4DJE4nfF4a�F44G4�+D4ǓF4�AG4�&G4<G4�IG4�'G4�G4�3G4�@4N
G4�
F4�iE4$F4ÃE4JG4He?4
<G4�bG4G4��F4[G4�qF4�G4�G4n�F4�$G4�D4=�D4��F4�CG4�F4FSB4��F4�G4��F4�rD4�-G4K3G4.�F4�vE4��F4`�F4�IG4�5G4��E4[�D4�F4�:G4!G4��F4�'G4!�F4 G4T7G4��E4 �F4��F4� G4RXG44G4G�F4:�F4�
G4AF4��F4ȦF4U�F4IG4-xE4,�>4 MC4��F4|E4�6F4	zB4G�F4�]A4��F4uG4K�F4͢E4�JG44iE4OG4T<B4��A4�=G4�F4?AG4�{E4~�C4��E4��F4ZG4;F4��F4�4G4�6G4N�E4>pF4 �F4�G4��F4e�F4T�D4��E4�7G4�>G4]�E4|�74��E4�^F4�:G4�E4G4�"F46+G4axE4�G4�G4BG4��D4/OC4�&G4OE4IC4J(G4�TE4.G4a�F44�F4��F4��F4G4�,G4��F4�BB4�)F4+7G4�.G4��>4OG4��C4 �?4�pA4tF4lFG4��F4��D4�9G4{�F4�1G4�K@4BF4,@D4�C4qG4�(G4"G4Z'G4MG4��D4k�F4��D4�G4G4WB4��F45~F4y<G4s:G4�*G4��F4�!G4�GF4%OG4�F4s<F4��C4�cE4jhD4T%G4R�F4VF4xpA4��F4��F4��F4e�D4�tF4E6G4��F4KtF4G4�G4�G4	F4 G4�gF4=+F4��F4�F4KEG4~-F4J�F4��F4�F4�(G4�#G4��B4��E4�E4��F4�D4}SC4vG4�G4��F4� G46G4��?4#�F4>!G4�#E4�<G4\�F4E4Z�F4��E4.%G4t%G4G?F4�F46'G4��A4o6G4v�/4�F4s�F4D�64��F4�<G4<�F4<�B4�'G4��F4�lF4�?G4�3F4�F4�&G4�$G4,4E41'G4�G4J�F4#�F4)G4�54��F4MCG4��C4�SF4��E4� G4��F4B4�q>4C"G4�}F4H�F48G4�(G4��F4eH@4�HG4��B4�6G44�D4�G4�<C4ȲF4�^F4��F4�6G4H#D4ђF4^WG4��34�F4-G4�G4�G4.�E4˄F4�PG4<�F4n�A4��D4��A4>4�KG4�G4k�F4#!E4��F4�0G4(G4��F4��F4�PE4�G4��F4:)G4��@4)�F4�:G4RF4_A4�F4ݍ:4�=G4��F4�>G4�CG4jG4�ID4�D4n&G4��C4��>4��F4�-G4�!G43G4iG4��F4�F4@�F4+G4��F4-@G4�D4f@F4�G4bG4�G4^G4�DG4h�F4�F4EG4��F4{�D4�&G4XC45�F4�FB4f5G4M�C4]G4�F4F4:F4'G4�>G4�F4��D4YG4�#G4�F4e�F4�F4W<G4EG4�.F4�G4�F4mF4qG4�-G4AG4@.F4�F4Y�C4��F4s)G4��E4�A4zGG4��F4=�E4�G4��F4�C4��E4|:C47G4ܙE4��F4��F4��F4.g@4�D4G4NG4��F4�MG4�	G4f/G4*�<4�F483G4��F4v/G4"G4��F4�v@4��C4
TF4Q7G4�9G4�9G4�G4v-G41G4Z�F4_�
&�\J&���%�[�%�)
&��%�I�%J\&�%	�h&���%��%�ݘ&
�A&
@&ą�%n��%�u&�/�%���&��%I�%D
&OdN&>&{�&�m�%޻2%jF�%�[�%H�E&���%U��&^Z�%ٛ&/��%���%_�%&ƞw&��% �&�&�%�%�Z&�d�%h�%���%�&&�r�%g<& ��&��E%�c�%ˠ%x��%�Ɓ%ճC&F&��>&E��%}l�%t?�%��%�1d&�/�%���%�%�Q�%GZ&���%@�%�?|%��%)��%ta�%tS�%,�%r��%�M&ju&�ly%���%Ҋ�%��%�2m&��*&"f&Ǎ�%�z�%���%v�&DL�%��%���%�K�%���%^&-lf%��9%d&Yx�&��%�/�%���%S�%-��%ɒ%���%��%=��%���%�7�%K,&u��%��%PS�%��%Y�%G�W&�V�%��%��&ɡ�%�&_�&�		&�&0&��%<��%T	�%���%A!�%���%P&�k%:G&H�&��%�(&�X�%�U�%�4&�&�Z�%�x�%xN5&'�%	�%���%�8A&���%�5�%��%=�%��m%�#&���%?1&Ϋ�%��%,	&?��%���%'�%�r�%1��%K<%Xd&Ux&��%�2&)�%���%��$&7�%t]�%���&���%��&!�%}v�%�]�%Y��%u&u+&�׶%2&*	�%(7�%�x�%+��%��B&5ņ&�x�%�~>&���%쨡%�<�%���%���%���%�T&c�%�P�%��%?<&&(�&��#&|r�%O�%#�%�w�%�[�%��&�=&���%ʔ%��0&��%8�&+#&V��%�<&���%��%��&t��%���%W1&�ND&��&5r&��V&�?4&�5�%��%��.&f��%�jm%�_&g��%���%H�%�Y�%%A�%�]
&��^%W�.&��'&�Q�%H)�%�\&��&��%��&�!�%Ů&9&�%��%v)&�5�%�h&P,�%77&b��%���%�ң% 6�&S�%�ɂ&ϛ&�z�%��%VQ&�-�%"��%��&�y%��%E��%�"&��%��%je"&Px�%�(&�R�%�&�%6�%ro�%R�H&��&���%�t&�%+�n&���%�h&j�W&v��%#-�%߾%=a�% �*&QZ�%D�m%9&�0&��%UX�&�	�%h��%5�%O�%;�%S�%���%��%�$&�ٚ%�[�%�¶%g��%�)�%���%vey%��%cՈ%5R�%��&���%�-	&C�&] &;��%-��%Uu&y�&\�&(�h&�ӭ%6N�%R��%��&�֗%��E&�� &{�&@E�%���%��&�Լ%���%>kX&� �%�?/&��%1Ү%5Ԣ%y�.&Q�&�D&z�%&l.&�Q�%�w�%�� &ֳ&&&���%B�%�T�&NQ&R?&�d�%�˥%&&�%.p&[�%�&m&�%�H�%�N�%���%��(&��&��%���%i��%��%�W�%���%t�&���%0׍%��%~y�%3��%��%���%�j�&�%�x%:Z�%�e�%�z�%���%$��%��&%��%��F&!�&qOB&'9�%��&��%t&�?�%<y�%r��%�Zh%j[&f�b&@.�%�Wa&R3&�w�%M��%4&`�%~�P&�e&�h�%��$&y(�%j�%���%¡�%�z�%�%`-�%$E?&@%b
�%���%̱�%�vP%w>�%�*�%Rc &�k�%�-3&.9&��%�*&a)�%~�{%8�#&�{�%�@&g<�%q/&'D&���%߯%�`%&��%&��%s*�%�Ӹ%�p&j� &�w &s��%}�&��%�T�%a6�%	�%)�&���%v�&p��%ֹ�%�X�%�B�%��^&�T�%�_�%^a�%!a�%�&ry�%n�&��%՟&�<�%�4�3s�3>W�3d��3�m�32��3)�3�3�ˬ3�b�3fy�3Xa�3�3 y�3dv�3��3��3Rj�35=�3O��3I9�3!��3Ҟ�38�3�q�3n��3��3��3�
�3�=�3�A�3h�3C�3(d�3Ղ�3f.�38�3��3�?�3Mb�3�%�3o��3n�3tc�3�y�3�d�3ҁ�36p�3Ur�3`�3y{�3.�3̊�3/b�3��3qn�3hw�3lf�3oh�3��32�3�U�35��3O�3'��3Wݨ3aj�3yƬ3`�3hZ�3�g�3�^�3AR�3�@�3Kl�3�
�3��3�p�3J�3�h�3M[�3���33�3�3��3�7�3h�3�B�3K]�39��3��3�n�3x]�3�A�3ݙ�3e��3��3�j�3�q�3~x�3U��3�&�3Y�3R=�3l��38y�3�Ȭ3�3k<�32F�3�5�3��38��3iQ�3���3�/�3�w�3���3E�3���3���3Nd�3�ߠ3�լ3@�3�j�3
J�3d�3�c�3���3�*�3�P�3@�3e�3ӫ�3
�3�R�3Wl�3j¥3�j�3t�3f>�3t_�34�3�۩3�Щ3�[�3�{�3i�3�ì3M��3�8�3�B�3�b�30�3��3�-�30�3�C�3�ߤ3yH�3�w�3�I�39�3z�3 u�3�?�30}�3]�3zU�3�a�3��S3`m�3��3���3�ͫ3�{�3m��3���3���3�g�3�n�3c9�3A	�3���3�Ŭ3���3[��3U�3ϰ�3S3�3.��3�(�35�3�t�3 �3a��3ZE�3�,�3@��3l$�3݋�3���3�L�3�ɬ3��3�F�3�ɨ3v��3��3�G�3qv�3�g�3��3Mi�37|�30C�3�p�3:��3\�3�ݫ3�F�34T�3]�3���3�|�3�f�3��3a��3�T�3���33q�3��3P`�3�s�3qT�3k�3��3�j�3�b�388�31�3��3�T�3Ia�3LW�3;̩3�Q�3-{�3�i�3�}�3��3M%�32�3�f�3�W�3��3��3�G�31�3�Z�3˩�3:̧3=j�3u��3y�3W�3��3?X�3n@�3\�3*j�3i��3==�3��3�3�ī3�b�3�B�3�v�3b��3<&�3�y�3&�3s.�3�n�3�"�3�X�3�n�3)��3�׫3R��3�R�3H��3�E�3v)�3SI�36s�3�\�3
K�3j�3���3i;�3�E�3���3M�3��3���3�_�3�y�3�=�3�g�3�^�3&k�3Y4�3ќ�3^R�3���3N��3�9�3ˌ�3Ղ�3x3�3H�3�@�3D�3�p�3C�3�ͣ3a�3|��3���3(d�3��3b�3`*�3[�3�D�3�)�3�Z�3q��3�w�3*a�3b�3�$�3|{�3p��3H�3�q�3OR�3g�3�Q�3�#�3�J�3q��3��3O�3=y�3�:�3(��3N�3�@�3>�3+s�3�b�3�W�3�d�3�7�3/�3w�3ȡ3�#�38��3>^�3#�3��31�3[��3���3�d�3�
�3C��3���3�7�3��3�̬3�a�3��3qM�3rM�3�e�3'$�3 `�3�b�3*A�3�׬3��3-�3S^�3�v�3n/�3z��3�M�3�i�3�:�3���3u�3��3�B�37�3^0�3�]�3x+�3+�3�ˬ3N{�3��3��3�&�3�r�3Z�3���3'��3���3�j�3&f�3���3Gp�3���3�4�3�l�3��3���3�+�3� �3�`�3���3�Ԭ3�&�3 Q�3돭3>լ3�Q�3.�3�o�3|Z�3q�3�b�3��3Qx�3��3©�3�v�3J֬3���33��3�N�3d�3�3r�3,�3rF�3�.�3V�3���3Qެ3��3퍭35B�3�~�3��3���3W\�3!j�3�[�3���3�K�3f��3ق�37Y�3P��3�o�3�j�3WO�3Z��3,��3#X�3�J�3į�3�g�3�w�3�\�3[�3q�3�k�3咥3횭3�-�3�ܩ3r�3$Ӊ4���4=�4.5�4G0�4��4��4T9�4`S�4BF�4ܨ�4y?�4(��4,$�4�H�4�]�4!M�4+��4�f�4��4��4;��4.��4�6�4C��4�ю4���4Tr�4�P�4!��4���4�4�4���4�1�4�4���4�4�%�4�Ɛ4齊4V��4�P�4��47��4ѭ�4އ�4�<�4���4Fj�4� �4!��4���4�I�4D:�4�E�4���4�d�4�T�4	R�4���4�ܐ4Wr�4L&�4�K�4�m�4�ى4�M�4���4�M�4dL�4��4Dk�4��4�4���4gy�4�X�4rm�4��4�Z�4�͊47=�4{Ǐ40�4'��4_��4�ڈ4�6�4;��4Ip�4�B�4���4���4�M�4���4�x�4���4�4�U�4���4�֏4���4���4I;�4��4��4k��4Ϥ�4=ޏ4O�4�Ɋ4 )�4W��4�א4=,�4�k�45[�4]�4�]�4�Ӑ4�k�4���4\B�4f��4�R�4���4B��4P��4���4�0�4ѧ�4Oc�4�U�4�I�4�-�4仉4�F�4�0�4Q!�4"3�4��4;��4L��4���4��4+|�41��4�|�4�P�4̇4FK�4�G�4"I�4�v�4(�4̉4�Ȑ4?�45=�4�f�4Lv�4�\�4�s�4H}�4���4?��48G�4Q:�4:R�4W��4a�4�m�4:�4�=�4�L�4Z1�4�̈4r��4߾�4T�4&�4�ϐ4�.�4$ؐ42C�4�ϊ4��4�m�43E�4>��40<�47�4"E�4�F�4}��4	^�4�K�4 H�4b�4hh�4���4涊4z��4*$�4ߐ4U2�4�\�4�P�4�%�4!�4��4b�4�6�4�/�4[��4�ˏ4��4��4-��4�i�4�-�4�8�4�u�4�}�4���4��4��4 ��4�/�41�4�Q�4�Z�4"��4 K�4[h�4W�4���4I>�4�\�4C��4D$�4��4�j�4Bu�4�.�4<v�4a�4���4Ί4.�4ж�4���4��4��4Q�4ň�4$ԏ4%�4^��4x&�4�4�@�4��4�p�4�{�4,n�4���4%��4s?�4��4]��4:��4��4_��4kq�4�t�4�֏4n;�4 ��42�4Ʃ�4YI�49+�4�6�4],�4�k�4���4+t�4lN�4<X�4��4�z�4�\�4��4 �4.M�4Y��4�X�4��4Q]�4%-�4�4�^�4�Ǌ4�D4&*�4�m�4�<�44��4n�4�E�4��4Y�4���4�a�4�,�4<F�4�c�4�k�4�Ő4�Њ4��45�4�V�4T>�4�։4�a�4��4�N�4u�4_��4B�4�X�4�N�4�І4��4��4�@�4��4vV�4
�4��4w��4���4
��4�\�4ܗ�4���4%�4:��4uY�4H�42d�4>u�4KÈ4��4���4<�4,ُ4떐4Jي4��4��4ʣ�4�ܐ4�X�4b��4�A�4w�4���4+��4?�4k.�44@`�4�R�48�4�Y�4�g�4��4��4	\�4ʐ4���4(j�4�2�4E��4��4�H�4�}�4�3�4��4��4��4&e�4�J�4?��4�`�4�R�4��4���4Cň4��4_?�4C��4�Z�4�k�4X��4b�4K+�4�Ð4�F�4Z[�4T�4؉4?=�4�4IP�4c��4>#�4�V�4}��4H�4�m�4T��4-B�4�D�48Z�4`y�4���4:�48k�4Rj�4�8�4VŐ4B�4�;�4�I�4cƊ4~i�4%�4�A�4�a�4#��4gD�4Ԑ4p��4f/�4���4�&�4�X�4�8�4YW�4F>�4�`�4�:�4��4��4Ŏ�4�/�4�4D^�4�+�4���4�	�4�;�4-��48�49Ð4�+�4���4v?�4�W�4�2�4�G�4,�4��4m2�4�\�4�4�4��4�Z�4"J�4R�4�7�4�`�4H�4�C�4 I�4�P�4���4/��4�]�4Cq�4$�4�y�4cÊ4o<�4�M�4�4�ڏ4���4�%�4yx�4���4���45��4���4��4�$�4��4vw�4n��4���4�,�4�!�4r{�4��4#��4,}�4{��4���4T�49|�4Ӯ�45��4(�4g��4�º4z&�4R��4���4�M�4���4@��49"�4L��4W9�4���4Ea�4Zu�4=�4,��4~��4���4p��4���4�v�4+��4&��4b�4��4���4o�4v��4�c�4>��4���4l��4��4�b�4'��4�+�4���40��4�u�4G��4y��46��4�4�E�4���4�4�0�4_�4��4��4#4�4�>�4_l�4S��4s��4�E�4�}�4�>�4��4cE�4P��4g�4���4"F�4e�4I�4R��4���4m��4$ �4���4��4�s�4?��4�4��48��4��4H�4}��4`��4���4�4���4�{�4�:�4X,�4�?�4��4U,�4=[�4���4!e�4��4�w�4ţ�4E��4Ź�4��4��4C0�4\�4T��4w�4з�4b��4���4�P�4��4�\�4��4W��4HJ�41��4�+�4��4�4��4�"�4C��4oM�4(r�4l:�4=�4e��4ԡ�4w��4��4vƿ4���4|�4/��4Y��4��4
��4`;�4���4��4=��4���4��4
w�4x�4<�4��4q��4-��4/�4�&�4M��4?��4BB�4%4�4�Q�4tp�4X��4p��4-��4A��4r�4���4G��4w)�4�@�4k��4��4�Z�4	}�4��4=��4d��4+~�4���4���4���4�r�4�d�4���4pL�4C��4&u�4B�4�f�4ޝ�4)z�4~B�4@��4&��4	��4���4��4N�4a��4��4���4#��4�7�4��4.�4��4V�4_�4hV�40��4�0�4�~�42��4�X�4k��4c��4I �4��4���4Բ�4Ɠ�4���4��4d��4|��4���4OY�4PT�4W��4G��4ע�4w��4�6�4���4x��4_��4��4r�4n`�4{�4�6�4��4s��4#��4�0�4o�4���4���4�8�4?��4���4�N�4Ɋ�4�4���4��4G��4q$�4U~�4
��4�{�4[��4���4�]�45��4S�4�5�4A/�4?��4�B�4��4�H�4f�4v��4J_�4�z�4Y��46e�4���4#��4��4�y�4���4���3?|�4���4���4x��4�x�4<��4�l�4j��4�4��4���4{��4ؿ�4R�4���4uˊ4�]�4���4���4�ѵ4�>�4���4���4a��4���4���4���4���4ϱ�4\E�4�:�4���4�4��4<i�41Ʌ4 r�4�|�4���4��4Y��4�:�4�)�4�v�4_��4=��44��4���4a��4��4g��4��4�4�K�48��4�O�4�h�4]�4��4q��4[��4���4-��4�.�4.��4W{�4���4���41w�4�;�4���4���4Sp�4��4 n�4�4=e�4��4ʖ�4���4���4.��4	y�4|E�4��4��4̄�4d5�4UԲ4�Z�4�h�4)4�4���4�u�4��4�.�4_�4d��42^�41��4ӱ�44��4�y�4��4���4f��4B��4�w�4J}�4���4`�4�k�43\�4
��4���4���4Oy�41��4c��4�6�4(�4���4i9�4���4{w�4!��4���4l��4�Q�4s8�4�5�4+!�4�E�4b8�4[/�4E��4s��4��4�!�4u��4�L�4��4���4���4�J�4\[�4�+�4��4t�4y��4w/�4�R�4���4v�4-��4��4���4�d�4�#�4���4i��4b�4��4�J�4�A�4���4���4f�4ܩ�4,��4�f�4���4��4u�44��4��4o��4�e�4�6�4h��4XR�4���4Oo�45s�4�4|��44z�4���4��4=�4��4U��4���4�b�4�E�4n�O(~XI)Au/),=)�Y))�|(br�(�')��F)�Q>)*�~(�E)Gܱ(��<)���(��)��@)F�-) ��(�))�1)f��(�S@)��W("c@)H�B)�p)".)��))�#?)�+)�ub(��)�!p(�uD)Sw:)�HB)k>)H�)Rh8)^�9)�:2)�=)xSF)_�?)��(F�(b:)}��(s�M)P�E)�(O)f�9)��))P�B)�?)96M)�K)�K)��u(5�@)��(b�C)�͵(�H)��N)�,)K1P)�J.)6X�(�.3)��/)�#E)�q8)+eL)��?)�]<)J�")��4)z>)�23)���(�H)P�R)�3)n��(�N)�62)��A)f")��H)E)ٻ)��M)��{(�))ө�(��4)$mK)@OA)�cI)��D)�oH)��)��L)�F)J�E)�SD)��3)��9)��)�/I)W�-)L\�(�
4)yg)s�C)㙛(Dn6)��.)�A)�){�E)�3�(�:)��.)�W6)�<)��)]�@)�C)��6)�{;)�F)�f(���(�N)��](��(wZB)'x=)PM)��D)v��(%��(��)�K)˩5)؎6)��(��1)�])u@=)5�(�)H)�zF)��K)�F)��H)w/D)ٴ�(�H&)t	)���(�({�')��-)"�L)��A)V;)E(I)A�")~�-)$K9)'O)3(!)�3�(��>)�J)�:1)IG)&�P)�C)��(M�;)�cJ)���($�+)pW(�?I)��;)��E)Vn(��(
kK)�=)Id4)�@J)��G)�nC)�F)㘌(~(M)ۚ+(I+5)H)-)��<)��L)�_)z�0)�C)�SD)e\;)c<B))�)�J)p9G)s�(z3F)N?)��!):>)��L)t9K)<�Q)�D@)�+�(�pH)�"�(��)�W)��C)�:F)��C)7�4)�9)���(7�7)k.5)��(���(*�(C)A)vWA)e30)�O2)�x)Rb)��H)�9E)�M)���(f�H)�Ɓ(�5(@)�(o�E)K�:)q�4)-�)փ<)�3�(�z)�>)�*)�xI)�fJ)*9)�=)E�D)(�#)i��(�D)��=)�f;)m6))>)�*)/��(Hq3)��L)B�}(�;')��M)!V�(��0)Q.M)<SK)�u ),�))J&F)�-u(�mJ)��I(��3):�/)��%)`�M)��)&�;)�G@)�(�(��b(�H�(8�I)M��(m�)�RN)��G)��(�
)�m)�T(uA8)�(Kq).h;)ch�(7(�i�(��=)cO9)\E:)b�()^�;)L<>)�u(l\?)W�)��(�
B)H��(�H)D��(��C)0(1)k&�(�p%)��F).�(��=)�4)T�J)L\H)k.N)�>)�&E)�>G)�E)*�N)�=)=�R)�zH)��J)��?)G�Z(�61)_72)�C)�.I)��%)_Q)�1:)h�H)ƁL)R��(O�e(X^C)E�@)�69)H&�(���(CO)^6E)T�:)5)h�=)E�8)E�7)-r�(��)�I)MH)q�){�@)a�2))�)��,)�2)>��(\
M)_��(C()�9)ޕL)N�@)�r)QEC)�oP)��D)wP)%0)&k+)�)�1�(�	F)��=)[�')D�6)j�5(w�B)�Ի(ݤK)jkN)�F<)hT4)�t�('i�('�F)��9)4�G)Δ5)F>5)�B)�H)3dG)Br3)QHF)6A)�֕(BwJ)��*)�z�(�Y()w�C)��$)�C)6s@)d�3)O�;)w_�(�H)�@L)i5)��?)�uA)� /)g>)wqj(��9)�KN)e�A)f(F)��2)(�M)M�J)��?)��) ]B)�FF)�D)x!)�/0)��.)��A)��(-91)�4)�*�(� E)X!K)�t(P{E)3rE)�N)?VL)afF)��9)�H)���(�;A)Dc7)F�(ߛE)�0)le*)��.)^^B)�_=)M�&)�UA)i>�(���(L)"�(��/)��-)��I)��3�M�3�)�3���3�:�3PJ�3I��3I$�3�0�3���3���3Z�3�U�3ޞ�35A�3��3';�3i�3�A�3�5�3 g�3J<�3�=�3~��3o�3���3Ժ�3R:�3�V�3���3D��3��3]�3�)�3���3�5�3���3��3��3�4�3��34[�3ɫ�3���3�3'9�3=�3��3#N�3ݷ�3U��3x��30(�3&0�3{�3�J�3c=�3�3c:�3��3��3�:�3^�3�4�3zG�3��3���3��3A=�3�k�3��3�0�3�$�3���3E>�3)=�3F0�3�L�3�3�3�)�35M�3���3�*�3��3g�3�	�3ܑ�3�K�3;!�3vO�3�]�3��3"��3)�3Te�3�9�3*�3��3�%�3���3rx�3���3c<�3���3�H�3%��3W'�3���3�q�3�>�3]+�3��3`�3_��3���3�D�3H;�3���3֙�3��3�H�3�1�3���3}�3�3{��3�4�3��3���3���3�5�3NQ�3�2�3�!�3��3o'�3�:�3���3���3��3�0�3Nd�3 ��3�@�3Q��3���3&M�3�0�3%�3�'�3���3S�3���3���3y<�3wi�36�3�#�3���3
X�3���3�M�3z��3��3���3���3�3a!�3��3�'�3�8�3���3B[�3���3��3���3/��3�b�3���3�*�3�&�3���3�g�3j��39Q�3�F�3���3�;�3)�3�4�31r�3M�3��3 �3���3�<�3�'�3*�3Q�3'@�38X�3O�3���3W��3���3��3'�3�3�3��3�7�3�$�3g5�3g;�3(h�3�!�3A��3�l�3�9�3W��3�M�3U��3���3'6�31��3�$�3m&�3�F�3��3:��3��3]7�3��3.�3�3���33��3I��3��3�"�32�3���3�x�3z5�38�3�.�3���30�3f�3`P�3���33.�3���3_��3�l�3��3J��3]�3=7�3/�3���3\��3���3$��3l5�3#��3�z�3��33*�36�3��3`�3�q�3@H�3���3T��3�L�3t;�3+�3��3.�3�1�3*$�3���3'��3y��3��3���3rd�3��3��3���3���373�3���3���3_�3��3E2�3F�3��3���3��3��3L6�37�3?��3�.�36��35�3�E�3��3���3��3W��3�,�3j�3��3�.�3���3(w�3�A�3�4�3.��3|>�33�3n�3�9�3(<�3��3e��360�3P��3��3�C�3���3�U�3���3��3���3��3f!�34+�3���3��3*�3�!�3i��30�3�Y�3���3�:�3���3��3��3��3���3��3�D�3K�3��3�N�3Z�3���3�4�3�4�3D�3a��3qn�3�W�3��3N��3w��3s��3���3/O�3�%�33��3F�3��3c8�3;C�3���3%��3)]�3�3�3ó�325�3Z��3���3�Q�3�3���3���3��3::�39��3AK�3�K�3�
�3�B�3P��3�&�3�s�3Ж�3��3�J�3�-�3>9�3�	�3���3���3���3�3�3���3FT�3 n�3y2�3h�3���3��3��3�^�3�
�3���3 �30��3���32�3��3(��3
K�3\@�3���3,�3��3*�30�3�9�3�E�3I��3���3�#�3=1�3x�3���3��3tF�3(�3�E�3G8�3��3��3B!�3&L�3j.�3��3���3���3M��3e)�3:��3c��3�-�3%��3���36,�3?��3���3z��3>�3FU�3y��3���3���3#��3Y7�3E�3�4�3��3��3@C�33�3�?�34y�3&��3�U�3��3)-�3-�34��3�D�3ٍ�3Q�3B�3rC�3�I�3�'�35<�3��3���3n|5x�{5Ǟ�5���5���54~|54d|5���5V͂5NUz5v��5��5�I�5���5���5�[}5��5v#|5���5��5E�5_�}5��}5���5`g}5x��5�}5C��5	т5s܁5�'�5�v�5G�5c��5�.�5h�{5rQ�5�u�5G�5��}5Xt�5J7{5�y}5c�5��}5+|}5�Ё5�Ɂ5�ς5&j�5��}5��5���5ы�5I��5��}5L��5���5���5yZ�5O �5��5n�|5�}5Uʂ5�(|5b��5��}5��5'R}5�^�5-܂5ͫ�5x�5��}5�'�5B��5g�5��5G��5G�}5{�w5I{�5��|5l�5���5�z5�}�5�w5�؂5*��5&i}5O}5)ւ57�5�Ƃ5�3�5?�}5���5y��5܉�5;�}5"�}5���5�̀5��5��}5�}5S�5-��5�}5j�5'�5��55��5`҂5�|5�{{5�=�5���5��}5n{�5��}5ӂ5�k}5�W}5S5�5��}5~��5�}5�͂5�̂5E��5���5�{5�}5���5.{�5%��5��}5�$�5:+}5$J�5h�5��5�{5N�y5|�5�x5���56��5,��5�5v~�52�{5��5	5�6y5LՂ5�~}5��5��5�y5y5�5~�}5`��5]4}5���5 ~5���5��5�O�5鰂5���5-��5: z5�{5��5K��5���5{+�5�=t5�]�53+}5q�}5~�|5���5	
}5�}5��5��5%Ȃ5}5�E�5��5���57�5�/�5�ւ5U#�5��}5�}5�n�5�v�5&�z5��|5N˂55��5�8�5`܂5��|5[�~5��}5=�5�5Ny5#�5k�5���5�ǁ5O��5�=}5��}5�56}5���5x��5��5=��5���5��}5�ۂ5H�{5��5T�{5a��5|��5Q�y5l��5�Z�5��5w�5{��5��5S��5�R�5��}5g��5�G�5y2�5�5z5�q�5���5;؁5<@�51y5�}54V�5�y�5a��5���5���5P}5s"}5��5Y}5k�5�W�5=�}5���5R�5��5�]}5��5�F�5���5�}5�K�5�}5���5��5̀5P��5�^}5D^�5�5۔�5,͂5��}5Aہ5�ׂ5�Ow5�S�5$��5<1�5.��5���5
��5��5��x5���5��}5�4,5v��5æ�5Juy5�}5�*i5 ��5Jg�5�ew5�K�5��5㯂5xπ5�}5�2}5 O�5~5�Yz5{��5ꡂ5s��5�|5�}�5�=�5�͂5���5��}5��u5!ւ5���5Ԣv5�t|5D�|5ę�5q|5��5�u5מ�5�z�5�}58�5���5x�}5��5)��5S��5���5~��5\��5.�5-�y5�c�5�D�5�R�5��5W)�5�~53n5}�54�}5�K�5~��5t�5�$}5�݂5��}5Q��5��5�m~5��{5�؂5s��5�5���57}5F�}5���5��5�$�5�=�5���5j��5j�}5�x5���55��5k}5�$y5��|5ͦa5�Â5@��5�t}5+��5{5��5QC�5%�y5W�5~5�
�5*��5ۂ5|5�`}5���5�J�5d��5���5���5Y8|5\��5�l�5���5_�{5%��52}5��5�ǂ5��}5��}5�I}5d��5`��5x�5��5az5΂5K�y5Y��5s�5���5��|5y�|5�}5�k}5u�5ځ5U��5��{5(��5�9�5ܽ{5�k�5�=�5��|5�{5��|5`ς5x�|5ˠ�54��5LZ�5��z5٠}5:�|5�|5�
�5��|5�h}5��z5W��5˰}5�Ѐ5c�5|ۀ56�}5U��5��5�u�5"��5G�5Nq�5��z5��51��56�|5�ӂ5阂5{�|5�}�5DĂ5?Ƃ5�ł5���5�,}5�<}5�%�5�;}5��5�z5@��5��}5��5j�|5:e�5&��4˱�4�`�4�4�X�45��4�,�4b{�4�?�47?�4q¢4�4q(�4��4߂�4m�4)M�4��4��4���4��4-�4(l�4襢41)�4�	�4�&�4���4���4DU�42-�4;Ĭ4n�4oK�4^#�48�4�L�4M �4T��4�t�4e��4�;�4��4?q�4`H�4���4���4拧4�{�4�?�4�6�4���4%k�4�y�4=�4�C�4�v�4v��4�C�4�[�4Q4�4ܧ4sٳ4n+�4��4�ç4W�4_˧4��4߫�4m;�4;n�4�0�4ӳ45�4�4��4D�4b�4-S�4�ɓ4{�4�Y�4AU�4�4z[�4�Ȧ4 ��4f�4�s�4�Z�4bX�45��4�Q�4�ݳ4d�4S�49�4db�4(��44��4G�4�p�4�G�4ߋ�4�l�4�Z�4� �4�
�4�o�4�e�4�B�4��4l�4��4�7�4�l�47�4��4�{�4�Y�4��4�9�4$г4�?�4�E�47�4�b�4��4�4�T�4ې�4%�4v��4	��4�$�4Q�4 ��4���4^�4N4�4a��4���4�M�47�4�6�4�y�4/s�4A
�4��4/ś4d�4�b�4]V�4�|�4�?�4�§4а4a�4�w�4��4��4Ħ4�߱4L�4�ɖ4�m�4u�4��4���4;~�4��4��4I�4��4�§4H?�4zc�4�/�4���4�e�4�h�4Z��4���4���4\}�4߱4�Μ4�/�4*M�4�A�4�A�4��4��4��4�<�4��4@�4}�4Y��4c�4��4
��4:��4茧4Zݧ4ks�4D�4���4���4;��4d��4���4�ǡ4�٧4~�4eg�4 �4�1�4+��4KM�4��4��4�٦4�1�4$�4�H�4��4Y�4���4�4U\�4�Բ4a&�4��4���4|��4P�4	I�4�h�4���4&س4É�4���4�@�4�4�4�4�Ƴ4���4�O�4�|�4X�4�Z�4�H�4<h�4��4�-�4�8�4ᢧ4��4ּ�4W��45=�4 <�4�&�4C�4�ç4�^�4F��4F�4��4*߳4�б4;��4��4A�4ϒ�4�̧4���4۰4�=�4�l�4k]�45��4���4���4�I�4,ڤ4"�4O�4.>�4��4�j�4  �4Q�45��4�Z�4�w�4��4�å4���4PA�4�s�4��4��4>��4�ȧ4��4�%�4�"�4���44R�4��4�m�4\J�4���4�4*u�4ͦ4F8�4ο�46ó4��4>��4�q�4�}�4�]�47+�4���4>i�4m�4]��4/P�4,�4E<�4�N�4�R�4VT�4�"�4�4�-�4�l�4�x�4wD�4��4 ]�4ft�4�>�4!0�4t��4��4�q�4���4�n�4M�4Ǡ4���4芧4��4�˳4^�4��4]:�4��4�E�4�3�4�E�4�γ4A��4���4���4"��4��4`z�4 j�4�u�4Wb�4�o�4fl�4�|�4�m�4��4V�4���42�4���4ؿ�4�Y�4�<�4���4T��4:�4���4`��4:6�4���4�l�4o�48U�44�4搲4$ɐ4���4/��4���4ا4ˋ�4��4��4⠧4�ձ40ϳ4SȢ4ۙ�4���48P�4���4�W�4U;�4V�4�a�44��4���4�4�U�4`��4�R�4e`�4��4--�4���4/��4J�4N�4�v�4I]�4r��4z��4��4��4Q��4A��4�4R��4�4U%�4Yҧ4�Q�4���4���4���4̦4:
�4���4�4�F�4 ��4��4���4�k�4Gץ4t}�4+�4��4\զ4�B�4R��44��4׭�4O
�4j�4�=�4qo�4F��4/��4���4m��4Χ4�8�4��4Y��4S��4���44 B�4ϵ�4�@�4�k�4=�4�{�4{H�4�Z�4��4�o�4К4[�4�ԧ4�i�4�M�4u�4�/5),5K�5���4��/5�(5��5;�'5��+5b�2515�{25�05��85t/5s=.5�T%5��+5h'5�8!5�"5|�5}� 5٣!5qt15�!5��(5��95$!'5UY-5[�.5UK 5dp15�1'5�P*5��+5 h75�5P�5�"-5�E-5{�$5z�)5�75�Z5;4#5?l-5Ft5ݯ!5U"'5~~5n�/5[y(5�05�5 �+5Ȼ/5�5/�+5��!5q�/5h%5�%5>�$5�:!5%�25�H.5ۦ#5A&5+�!5�"5f�-5�5%5�)5�w5H�15�Y$5_5�65�	35�(5�Z5�5��(5%5X�5R5R�*5C5�b15G"5Ww%5��5�5^:)5s�&5��35ߋ25��&5)�*5K�)5�Q"5��-5Ŏ,5�>65��&5x�05)�/5�:5[W'5"�!5�`5Vf5�<,5��,5�&5�h-5�F5Q %5�E/5T�.5�/5�M%5�%5��-5��05��35ޙ(5�%5�5}�&5X'5�5B 35S�(5#)5+5=F,5#%'5Y[.5!*5�x 5Q�5��5�,5�5_Y5�S"5k�*5�?,59(5C$5d(5=65}�#5�!5K65-�.5��,5�05��.5��.5p�$5߃&5��05�6!5�m*5]�!5��5j�5��15(5NT&5��.5�+5�-5�e15b�+5Ɋ!5�s.5e�"5��.5,<%5��5�)5��)5Z5/�/5�5~&#5�5(5 5��5R ,5U,5��$5�N75?c15y�35q
5��75�75K�%5�+5b�!5.�-5�'5�"5ː5��5\� 5�35�#5rm5ۓ%5 _ 59%5�/5��5��	5&5�.52z-5})5��(5�-5��%5އ.5��15��)5�^5E�5	�$5W/5��)5�&*5Ơ(5p�'5+�-5I�55D�+5�-5U�)5;�.5��(50� 5e�,5I-5S�'5&�#5�+5��)5�|%5g�25��%57�-5F)5'\)5r�05��.5�125�*5��%5u)5��#5��+54@35`"5��5d�5�25ӹ5M�#5?/)5gZ5m{+5��15�-&5�-5b�+5 �35cU5W-35(�-5{55��5,5\e5s*5�z/5��)5E�!5��5�25�B)5}�5܃%5n05��85y�-57�5� 5<O55Ż"5�65�-5�+25O235��,5��#5IW5X�
5@�25,k%5�5'5�&5�5�(5��#5V�/5��%5Ke(5ڢ*5x25��:5ڏ5��'5��%5 �)5<$5Ј-5�8!5:�!5�35*e55��15}�+5�235��5h�$5Y�'5��5��&5��05�>.5 7+5},5o95��,5��#5y&5 >05H�&5v�5 �	50+5|'5H745�#5��,50�*5>*5tX55C�05M445K�!5�+5��&5G�5V�&5��%5��(5��$5�6,5��35 R5P225�5��-5-\35�
,5�$5��5� 5� +5��5`5��45�#/5��5�+5<].5�=/5��5�o35�	35�45�q$5�*5�3550$5V�,5��-5�G(5?�5�'5F#5T7
5�c,5��*5�35��5f�/5�$.5T�(5�A#5E,5Ш+5��"5�E5��5�|'5��5^�,5�M5�� 5�[!5n45&.5�%5�5��'5tG%505ې5=�#5�z.50/-5pH5l�5��+5]#5:�(5Yr5�6$5"t%5��5n .5Q 5��15ɒ05�B&5<h5�R#54� 5O+5̞5�H 5�M-5d�"5� 5�.5��$5Q%55�-5��'5� 5�)5�h05d�'5��+5�U5^�25�-5�!25-�-5��5�#15�2&5:�#5�]45F*5G�&5�%5�25�05ݕ%5�s#5�E5�5��*5Y#5�1#5><*5�5�-5�-59�55�R4�N4��M4��14ز74�<4�N=4uf@4W�G4��D4��E4+;M4�Q;4�lL4_H;4M4��A4Y�C4�KI4�]K4��O4��L4�I4��F4��J4�N=4w)<4L�94��74ºB4݈F4�;4nzF4�6P4==4QE4�ZI4/DL4n�I4�"G4�MM4�J49BJ4�bI4)�4�PN4��74�I4��44M4Q�N4a�L4)�N4	lP46YP4��C4��N4�v4�=4�~D4R�J4�H4�4�bF4H�=4�C:4�NJ4(�O4d�E4�L4�J4��F4��J4M4E14"2M4�m>4�S?4��P4P�H4YH4�qG4j�B4�&4G4��84v�>4�?4|>H4�3H4�J4��I4r�H4�B4�-4�G4;
S4��G4b�M4��O4�4��I4�L4��F4�qH4�!46�H4��K4-�I4�>P4��N4�4�G4�MI4y�F4��I4�C4�'4�f,4�4Q�H4+H4��O4�L4,64��K4�@D4p�H4��Q4�4uM4E4�'>4�}L4P�24��G4�J4?�F4��K4�M4h#4 'I4�F4�K64�,H4ЌG4*xI4��K4k�G4N�H4��M4��J4�N4T�D4��941�G4GK46�Q4U�74{484�54�JP4Q:4$�,4yD4��I4��/4��F4�4:5I4�.E4H��3��L4�pI4�k34,�I4�cG4T�D4�!I4��F4,�G4�]M4��-4¼@4*K4s�I4�94��F4�+4{4I4�QH4�F4�/C4��54dM4^=N4D�=4��M4UnG4j+G4�~D4��L4��H42�G4�-N4�L4P4>E4@�L4�4�E44#4�RH4)H4N�E4��*4�*I4�K4� ,4.�G4�4��*4�/C44�/4ίH4�=4^C4�N4a�H4��I4��F4��I4��K4q%G4��M4�4@�G4֏@4��F494īF4�>4I4��I4R
D4��P44�L4��94��J4TN%4<cD44�4�*4��D4_bH4�O-4��L4ڢL4�^M48}L4?4��H4IE4�ZM4n�E4+, 4�I4�;H4}�F4]�I4��N4F;4�G<4NyJ4��=4�q<4eJ4%�C4�hN4�<4r7F4��E4M�R4{I4�iM4��J4�]D4J�74;|�3�uG4e�;4�24~�M4%�I4��O4,_4D�4��F4�?4K4n�P4�D4_x94��N4`�N4	�G4S�B4��D4/;4�rG4��G4k I4חQ4P�F4o}H4- 64�;4��44�VI4G-M4w2?4��J4avD4��H4��F4@�B4ߞK4�-M4�
4��.4DI4]M4�BI4�74^�M4��=4�I?4/uA4?�=4�v:4��E4�)H4�Y74;�F4��94�Y64��94�aI4�lI4��%4a�F4QFH4�;4zO4�'64LE4��K4oD4jxF4 �P4h�L4i�-4�I4ժH4EG4��C4*K4�~48�G49�R4�=4!PF4��M4��F4PgE4�NC4��F4��G4��D4I=4�D4dC4��K4�sO4Y�:4��G45X<4q�H4��F4}[J4�J4��>4"I4!H4a�F4k�F4_�S4 H4T�M4�-L4�~4�D4)@4��G4%�E4�tO4?uG4;�.4��E4@�O4_�94�e>4� J4�0:4��H40�O4��4�A64HTF4/ ;4I4/�H4woA4��I4E4�4a|H4�!14Y�G4e�I4ϺC4��K4�B4�%4�_4��O4�34��:4%XI4%G4��N4D�N4P�H4��D4*�H48�F4��=4��M4cW;4�M4p�/4�kO4��L4d�K4-TE4��-4�V-4?�74�NA4M[H4�D4�TP4N4%xH4&E4�:4��14DJ4�f849�H4�E4��-4L�4�>4qBF4�m4�64�zJ4r�C4-�H4_�J4X[L4 B4�M4��G4��O4�;
4��I4/�I43�H4��J4��94�rF4�[64Q�Q41C4%�I4#�E4�nL4�SH4:�4-�4L؀4op)4�#�4�U�4���4���4L�4N�4���4��4h	�4���4�w�4��4�4�4��c4A7�4�4�w�4���4���4��4��4�C�4i��4�!�47�4wv�4�|4@��4y�40o�4'�4Ĺ�4Mu�4;��4˄4���4�4@Kt4��4��4�1�46��4�4� �4փ�4�ؙ4�0�4�m�4��4��4q:�4��4�O�4מ4j��4l��4牙4A��4���4x�4E��4�d�4(|�4��4"��4*��4�M�4�`�4*r�4�'�4��q4��4R��4lh�4q�4�J�4���4�.�4��4�4���4��4|U�4H�4 љ4q��4���4;��4�d�4�,�4���4�&r4�v�4�K�4L��4.A�4�ə4@�4�<�4�6�4��4��45%�4�4;��4��4a�4���4F~4��4���4��4]��4���4���4L8v4t��4��4�	�4�{�4v(�4آ4J̨42��4���4V��4��4��4��4��4���46��4�!�4���4�͖4!'�4�;�4�<�4]��4��4G��4P�4��Z4`�4q١4�l�4��4�_�4q��4T�4$3�4ay�4�4���4:w�4���4ZL�4�f�4?×4�q�4��4�4���4�4��4���4P��4N�4�Ȝ4�4f�4�`�4ppv4vɠ4���4t>�4�>w4���4�O�4�y�4~��4��4/�4��4��44���4NQ�4"�4{��4�ޝ4.Fa4@��4�$�4
J�4c��4܋�4Ʋ�4���4<M�4Q<�4pĖ4S��4�ג4ҿ�4�@�4'�4ܒ�4��4\.�4>V�4�;�4��4 �4���4�p�4?�4g�4s�z4+R�4(7�4dS�4���4 �4y*�4�'�4(��4��4rU�4���4{^�4�9�4���4̑�4?d�4��4��4�/�4�n�4�4K��4�)�4��4=�W4��4V��4b��4x$�4AR�4��4ܒ4b�4�p�4��4ǻ�4I��4:ʘ4aS�4I<�4�v4�~�4�f�4ߝc4���4�̡4�֕4ȗ4l��4�;�4���4|��4�B�4�:�4Fu�4_I�4��4�}�4X��4��4�D�4o�4���4̫n4���4�4١45��44��4���4�I�4�4�ޔ4f;�4jK�4��4&�_4��4�|�4��4��4��4��4�{�4Nt�4�4�4� �4���4Q�4Rj�4��47��4�P�4�:�4GI�4�4I��4��4�D�4#D�4N�q4R��46ѕ4j]�4ō�4�~4�I�4HՐ4��4ME�4�'�4��4�-�4�r�4(W�48�4w��4뽚4G��4
0�4Aw�4ښ4B=�4	��4�X�4{��4�d4��4c�4vӡ4�m4��{4?,s4/�47�4��4��4b��4捠4��4��4�B�4(-�4+7�4���4D*�4�f�4�0�4��4Q#�49u�4<?�4�h�4K]}4���4���4۩�4a
�4'ĝ4�Ȗ4���4��4�4���4oO�4�	�4��4��4Uy�4�>�4$��4��4~M�4�"�4S��4=�4=\�44N�4��4h{�4���4��4t�4 F�42a4���4��4#�4I�4�F�4�К4.��4�G�4�ލ4���4e��4�]�4k�4t�4I:�4Y�x4!��4N>�4���4.-�4��4U��4��4w��4č4�B�4P�4~ڠ4���4�4`�4nՕ4��4��4d��4��4Ɨ4{U�4�!�4�o�4B�4B��4Fp�4ә4���4ݖ4v�4嬞4]a�4>��4�ԓ4� �4�9�41�4/��4��4l��44�4"Л4v�4`P�4"�4��4ah�4ܴ�4R$�4�$�4FP�4\+�4�^�4�v�4�K�40P�4��4n)�4歚4���4l+�4��4���4u��4=�4ڼ�42ޢ4�{�4�-�4p��4�ˢ4��4i6�4z�}434c��3���3f��3�>�3w� 4#�4�24)�4m�3r�4��4 y�3R$44�[4� 4�u4�k�3�|4h44I54�4-
4ͥ�3��4��	4ɸ�3��4�4��30H�3��4x34�� 4�4.�4�k44�� 4��4��3" 4��4�r�3,�4t' 4��4G�4��3[�4|434�~ 4��4�O�3E 47K�3��4#4U@�34 4�/4u(�3�4��4��4N�4�u4�04��3�: 4��4��4.,	4�~�3)c43�3�4f�4a74�ը3J� 4�4U� 444�4T��3O�4�P 4���3ʆ4�F4�4D��3=�4Ĩ4T��3	� 4)b4��4+�4G��3;�4�+4
Xa39�4��3۸ 4��4oB4��4N48�3��4q�4#4�I4�43�3�V�35�4�p�3U��3�4���3u��3�4�E4��4�Y4��46&4d{4B]�3h�4	I4U 4^G�3��3�e	4�t4��4� 4�m 4#]4���3�� 4�v4S�4�?�3��4g�4�44թ 4��4�
4V�3��45`4�H�3���3/�	4*14�4-�4�.	43x�3�34~o�3�X4�q49��3���3�S4��4���3�� 4���38��3�4#�4i�4��38 4�c�38��3�
4F��3*� 4`4?��3�4���3'�4���3��3d5�3_45X4{(4�G4�) 4N\
4sV4��4^��3�� 4��3��4?�3s��3�U4ac�34S4��4���3��4	�4�4�,�3)E4���3X�4�0�3$�4ǩ4�Q�3M�4)� 4�4�3�J�3�N�35 4��4[, 4��4�i4$� 4K*�3FO 4@4�+�3?=�3m��3�[4��3�� 4�4--4�4�4�4`:�3�A�3���3��4�4I4�D4��3�I4(�4<E�3��4��4�N�3��4e��3���3ك�3��4�w4�A�3Κ4w3�3XE�3E4+�4� 4W4��4���3���3�t�3���3,�4D�	4]� 4�j4&��39'4�l4� 4n�4��4��3���3�Z�3 4�|47;4P�4v��3��
4:~�3y�3r��3g��3��4�{�3r� 4M4&-4A��3��4��4�54��4[4?�4���3@�4���3]��3��4d- 4��3S�48�4��3 �i3x��3�44��4���3V4�C4B 4���3���33�4�U41C4ʬ4�\�3�<�35��3��4F��3{�4�l4<N4���3�4�3�d4�4�m�3շ4�v 4���3�3�o�3-4�,�3��3��3�u4cq4}74G`4:��3�� 4�4m#4e4�L�3q;�3W481�3)l4��4q4�	�3~�4�R�3��4@{�3]�3-4�|�3m�4,P4P4��4���3�4_�
47�4�24���3]3�3�X�3�545��3#�3f�3H��3�] 4|� 4"4v~�3�u4s�3j 4���3#��3�4T�4-� 4~��3'� 4��3�F�34��3�r�3�k4Hk4o�4iU 4��342�3� 4&H4��3.#�3�4� 4 8�3s\4q�44� 4��4p��3+y�3�4�R4��4H 4K�4G� 4�X4��3
4)Z4g�4���3�4�`4��4��4�4�4�3
Q4��
4��4Ʒ4�4ʤ�3@��3�&�3�4���32v4,� 4/�4��	4o^�3o�4kX�3T��3��4Q� 4m� 4�4�J4��3�4s|4�4��3�41�4H�3�"4ef�3�,5�]*5�*5�l5�55��>5',(5�k75j�25U<5�s45�:5U7+5Q0�4y�+5�495��45�
95�m25#15�/51�%5��*5�!5��&57%&5�35X�,5o~'5�o65p*35�95�55��4_;+5�@75bl65<45ni(5Il/5�',5�@45�$95�$5��25��,5�k35��856�05�H15I��4��25��/5aG$5`y+5� *5��!5��65��45=�65[�+5�5�85M|05|�15k�65}\35�745e+(5y�-5��35	:5(.5��/5,�5�85;�>5�� 5�D*5~�55\�%5Ln)5T�/55�-5P5��'5~�,5hd:5�@5Դ+5��95�q35x�5�5��:5T�:5��85c�%5�{/5̀75��35�05iG/5�s(5�R(5�t/56�-5T�65O(,5O�5555D�5R255�/5��15џ,5R�#5�~#5~4-5s)15��65��+5�75+/5v�55�25�<5-�05�/5�M,5&�$5t4/5��:5z35�5q35z�5u�05�O25e55>!<5��)5)"5K5�05�� 5��55M<5�F-5�4585��55>,5��35{�/5�)5m�05
�05
�$5��45ӌ(5�a,5b�15��15�55u�&5�'5ud25�#,5��*5��-5�Q?5*5�/5��75��65��#5�c05�/05jY/5�j*5a{85��$5685�o,5g�5�h05�55-'5�45�e5��15��5�85 o.5�+5�j75�&-5�q25�;5�L(5~65��5��,5!,50](5�m75�z75�F(5�5��5�(85�:45��.5M�45�/5��%5�25�-5;�#5;�5d�$5!�75�-5�75�D45��-5�25ϩ&58%5v45��+5��-5,�75h� 50�05/58�,5�15w�35Q�;5q15=@+5~�5��15bM75�;:5o�45��-5\�?5HB&5�w45�A353�25_:57}D5u*5�:5��15��"5S�.5�+75�45��$5J�)5�e#5�65�'75}X#5[w65��57e/5ߥ!5Q9,5�85�495LI25$5-�65��55�651/>5o�75�_+5|u;5�/54"!5.5�75�.5�Q85��)5��95�Q75�*5�7.5�>35�,5��#5�05v�75�k35�N/5�o25&�95��;5�c)5\n-5v+5�V 5�55�u-5k)%5��25Tj;5d�5�)5œ65�!5}5�"75F�45��25Վ15�t+5�	.5DG/5515�55��45475�u65�?/5�T4555M�*5O�75 �55v�;5��35�-5�B)5<J"5Ƴ5o�.5:!15A85V7;5��-5-L55�@35�#15��05�95Y�15�15�5ۨ%5�'5�!5��75Y65��45{�85F�25,5+�75�+5��15��(5r175kk/5l05S�05��*5.(5�15w.5�45�-,555��15��25�K45a�15�/*5k�$5<.5�+*5�m-5��25ۂ:5S�85��05�25�,5n35��15��75э%5�05v	25i�(5��25��35�:)50�(5��05cB.5A�;55!35i05��15�&5C�:5�05��65�$5L}35��/5��55M�,5�?05m�158R25,�5�( 5V�)5��.5�45�"&5Jz65�� 5�}-5j(5!=5$"5��75~E55�d:5D.5X�35%Y95�/5�S5oV25��+5��/5F�55�]5��75�{ 5�,85��/5�85��5��+5Y*05�e15E15�*5]65S��4R)5�5ӓ15��#5s�'5�25��(5�H65j05�$5j^#5��05�.5�S*5�q'5�i55�15d�0525!�65�N45��5\55��5t�05j@55�e5*254!51�=5�)5S:85.z75چ*5�k05��.5�;5��3>�M4+~K4Y�Q4�!H4::Q4
|L4�J4�M4�B4 4��F4�~>4dC4[D4�-4�iF4��K4i�=4��N4�H4�K4'�Q4+L4�Q4�tE4a�J4�\L4ViI4� A4h�'4�^#4H=4��D48�Q4ӹK4��M4 aE4��K4�(4>T�3C�A4�BI4��H4�J4�Q4av?4�kM4ǙL4<	F4�)4��C4w8D4��R4[�O4�!M4{�L4��M4�pL4�qK4_�L4��L4Ne"4�3%4��O4�fP4q_J4��O4zb!4��54�/C4�54�O4��I4�B4�J4��F4q�$4@FG4\�L4bP4;�B4�lO4q)P4��J4�E4��<4h�4v�M4f�H4/�%40�O4&N4��E48I94��?4��A4�*N4#�M4�74#�F4�#M4�?C4\�E4�?O4<rI4��L4D�O4K4��4�gK4
(M4��T4�C4QpM4��L4n}L4j�D4�>4߼@4�E4��L4L I4�H4��F4�.G4[M4cjN4K4&rC4�:64�gG4�B4�#&4}!D4h	A4�RL4��M4G��3��B4!�F4��I4��H4�C4�-4�L4TTI4k�H4PcO4��,4�G4'r<4�e�3Ѩ4yI�3#6>4w�Q4icE4��K49M4֣F4`	G4��@4d|N4�C4��K4�=C4[�O4��L4�-M4�L4P:Q4K4FR4;@K4��64��G4[�*41�N4��I4#�K4�/94�7J4=�E4Hw,4B�'4��H4�M14~�T42�I4��O4�PA4��O4��J4��F4J�P4��J4��I4.34ӮI4��4�IO4��E4�M4 L4ǃJ4 �D49O24&eI4M�I4M4�N4&4<�M4�I54k�G4A+P4ͺ4!�N4�N4p�J4"�H4f?O4c	E4ҢQ4cF4�T4�9D4�E4vM4�K4�/4v2447�E4��F4TqM4�M4]B?4�dL4��64W4��D4�[;4,xD42{T4Iu�3y:F4�AN4��E4"�>4"+;4��4:2>4��J4�G4TBK42M4�=H4��N4x�N4R4ˉE4vL4�L94�wH4]�L4i�K4�,N4oH4SLG4��.4Sj4�(4NcI4u�<4�EA4Og24�NH4AG4j0 4G�G4�J4;nF4�G4��K4":4m�4��F4/�I4��E4��D42O4�x)4�� 4�P4f,4Ni44��O4/�F4��C4��(4jI4�#@4��M4�>M4ݑN4�zJ4,�P4��L4<L4��I4��I4h>4��94�O4ÜN4��O4�,4�'E4�4��L4�EV4IM4V�M4c}@4�'I4R�O4��J4�d4�K4|G4�G4�BN4��H4��14ۿK4L�E4!�#4�pN4*x4lD4jyN4�J4�PL4��F4[�F4~�Q4ǰG4�M4��N4�N4�!@4�H4ïN4J74��L4|sM4[WB4�<4D!J4m�N4&�D4a�A4�G4PhJ4kA4�E)4j�C4�OF4i�M4o�M4>�H4E4dYM4�&74�Q4F/Q4�M4�N4S4��D4
aM4MBM4��L4�W?4!�G4QL4�pF4p�L4�SR4O4KN4�DJ4"74,�4��4�G4�J4$K4)x-4c~Q4��G4R+?4h�P4�L4��?4IN4�
O4}mH4(I#4ON4,aP4��?4�= 4/BI4ޮK4��)4>��3��M4]fJ4�Q4U�P4��/4b�J4�9L4�IE4�B4[X64�mH4�I4�VD4��P4K�)4��G4ҾQ4��D4��B4'=4�O4�O4ΊN4 E4�YA4L�D4��I4��14;M4eG4�
A4��A4��M4E*J4�W*4ǋH4�@P4wI4X@4��N4��A4.	G4�S=4��"4��D4�834�yI4��=4��@4oFL4�cF4�?H4�R4e�N4i I4�A4��O4~4G4
VN4�'4A�L4�H4��R4L�G4�(N4y24��I4rOJ49K4��H4��N4��G4�-J4�I4FNJ4P+L4�&C4�A4�L4>qL4��Q4+ O4�(�3s�4��-4�74s�-4�e54��.4�=4��24��-4��4�:4��-4��(4�%)4Eg4430344V�+4/�-4��4�(4fl4�54�1;4V�34P�34o�04Z�94�24���3d49�34O�+4$%*4P�-4j�)4#�14��944{A�3lq+4�i749`;4	04�,4��4`/4�)4��3s�54�b44l�(4�34�%4�':4wb"4�+4�-44��24'34�p44��+4w.4�84�g�3Ʒ64?��3TX%4O�'4jE/4n�844844&a(4��.4
4�O4464��84��+4i�:4��64l�:4�y24��64�_34�Y 4�?&4�44'�4ak34�!74VA,4-�4Z�24�6%4��24r)74|�!4n64�504ˎ94��04L�-4��24�54��04�04��34ϴ04�x04Q�;4�-4�84Vy)4�64G.048�24��94[�&4�f%4��4<�84��44��'4̉04U�/4U�74��/4z�34�n04S
4>N4��44a'4r�/4N�14B�3x�94�d24�"4�v54޲24�4�54�:4;�4zS4�d04�e74x�14h;�3Ρ34S4L]4� 04��4�M14�"84��44��34�4�>34�C34#�54(�74��84�C54�24��+4F 44��-4q�,4�(�3t�/4
�04q�/4|��3:M"4>24�&"4�14n�4;�4�)4�84�504�4F�&4�n84q94]74�54*<(4��24Ɛ14e_84�46;4@j+4�*04Wg/4;54rB54��.4]J14� 4��94�:4O�74|�+4x=�3T44��#4�614E�44�4.,.4D\:4�d24��4>�14�t64��:4��:464�J*4:�44��14�04���3a�4v�4��54J�94c~14@0�3��4k�44x��3��34�x44F�24a�44=$74%�14�4��94\~%4�k#4|�84�(4�4!44Fy24�C;4�v94�.4�<4��4��34��4�)4��-4�94�I84]�74�+4H/4�84�_24���3��84��04��&4�4�74՛(4�E4N)4"X.4%-4+
64��,4�c4n4�I;4m�4½:4^s94�;4��34s��3�$*4'�+4گ$4��/4RL4�t34�C$4��14ԏ4��34�04��$4!�:4��84��4�554�b14414��+4eC4��*4��,4n�74K�/4Mu94��4?e34�.4�34��14�|4�?54�84��24>z�3@+34$	14+��3'�(4<K041�4V�/4'�24~�
4y�44u��3��4]�24E~/4�)/4}�.4�44�Y/4O�34o�'4�l.4��64�:)4��-4�i/4�4�?!4��64.�.4��-4C[.4#4�14�[*4��04ð74A)4��*4z�+4�V�3�R-4��*4� 64�64� 04�4�224�R84�g04�_,4��.4\04��94�24��04)u$4�94(�$4c -4>_94�n/4�b14�44��-4l�64���3�"4ޔ04n�.4z
14��-4<8:4�@94 P4�/94��4��4�.4�54��14�"�34M,04��'4]�54��04u�54�V4�e�3�w.41�44U�4̷-4U�"4�04zX14E!4M�'4�b4�'44�v�3i�/4ױ64r�!4��24��
4T(44��44��)4D�14��546*�3��44{�+4��+4�z74��4�Z/4��4B�%4:
14�+4�@94r�04�!04D{94��3L4v84�U14��24�4�y4�-24C�14��34��*4�,4�74�/4-*24��94u54 H54�i14���3hQ74Ai4���3��-4p"54�B14*�64�4\i'4l4.4�)/4�L:4/�:4�e24�a/4��4r��3FL)4�s64��&4�S34@�04|�,4�n 4��4.x�4�4j[�4"��4c�4먿4᫹4�6�4�#�4Y�4�q�4u �4���4��4���4ݼ4-�4��4���4)��4	ʸ4v��4�x�4�@�4�о4W�4�z�493�4�=�47��46�4�V�4�754���4�
�49��40�4fԳ4���4ɩ�4�K�4B�4%�4���4R��4k��4\�4~�4~5�4x�44䵺4�a�4#�4���4�F�4�ʍ4:�4�D�4A-�4+и4�O�4�_�4� �4���4�H�4���4Z��4pҿ4�8�4��4���4�=�4���4��4�s�4?z�4���4t��4k��4=1�4� �43F�4K׾4}��4fE�4!b�4u��4��4'�4U��44�y�4a��4�Ͷ4�;�4��4$K�4w��4R��4���4���4>��4ʚ�4�Ի4���4��4�ʲ4��4��4�d�4Fڪ4F�4t'�4$��4B��4�k�4pմ4|�4���43��4s1�4ۡ�49��4�c�4ͧ�4E�4��4UF�4�ù4�Q�4+D�4�d�4.v�4���4 �4�Q�4S��4�C�4�&�4��4��4Q��4���4w�46�4��4�M�4���4�Y�4���4�4�P�4U��4෴4���43��4;�4�Ž4�@�4⤷4�	�4M��4ԣ�4c��4jx�4R�47W�4��4.�4���46�4��4�ڷ4�4�4,��4���4�.�4 ��4~G�4H��47H�4�,�4���4߅�4�׶4���4vc�4b��4Ų�4��4���4F��4��4y>�4%��4ۜ�4���4v��4覞4��4�4�q�4կ�4^�4��4���4�4˼�4�>�4���4U��4.�4N_�4�7�49"�4J��4}��4"a�4̾46��4��4�׽4.>�4��4��4y
�4��4��4݃�4�ø4��4'r�4���4�s�4�{�4��4�*�4[�4���4��4Q�4i�4�/�4���4�a�4"o�4��4-��4���4'*�4*��4#��4	2�4���4��4�ϼ4���4�4��4R��4�ʿ4 ٯ4n��4Ae�4��4���4��4�{�4o�4�k�4��4�49ľ4��4+ܺ4f��4�-�4|)�4�=�4@�4��4R]�4�ν4a��4�N�4��4��4
@�4u�4���4"$�40�4�?�41b�4 ��4弼4��4V��4{�4N��4wƱ4���4:��4;.�4���4^�421�4B%�4݌�4�2�4�c�4��4
�4��4�4?��4M��4C��4��4���4Uy�4��4�I�4���4��4�O�4��4$��4�X�44��4`e�4�:�4�#�44,�4��4���4m6�4	�4�4�F�45��4���4���4�4s%�4���4�^�4���4C�4�F�4s��4�w�4�^�4���4�{s4�r�4?i�4�7�4���4���4.m�4$%�4[�4�n�4̾�4���4̫�4��4��4��4tL�4ǁ�4���4�ؼ4"��4���4��4�a�4'�4w
�43�4���4і�4.˳4)�4��4{��4�c�4���4��4�&�4B��4�P�4Ծ�4`L�4�y�4Ӂ�4/ݯ4���4���4$�4���4mx�4�P�4�G�4��4ؼ�4赿4���4E�4���4��4&D�4I/�4�d�4vY�4pG�4�5�4_��4J��41X�4��44{�4xj�4i��4_�4�4��4�*�4h��4�P�4��4G�4Z�4���4�o�4[��4Ka�4���4~��4qG�46�4��4��4�8�4_�4�+�4-�4d��4��4#߰4�l�4�>�4��4��4���4���4O�4�J�4p h4	�4F��4<C�4�8�4���4��4_Y�4s��4�y�4[�4�?�4�@�4�/�4���4$ܻ4�g�4�m�4wd�4�]�4��4v�4�P�4I�4���4��4�6�4��4{2�4��4�H�4&��4X��4��4�4��4���4���4x��4D��4~�4*^�4���4T�4��4�<�4���4��4���4g��4��4D��4��4�G�4/�4���4^
�4��4��4�f�4��4$��4�k�46��4��4���4��4押4���4���4�V�4i�4Vή4ߺ4���4�'�4W�48�4F�4�G�4.��4��43z�4z�4Ԟ�4��4�4j%�4��4a��4=��4��4���4H��4*Ǩ4S��4G��42޹4x��4�n�4I��4W��4Kk�4�]�4 %�4X�4��4!��4��4*�48�4��4�{�4J�4���4���4��4���4c�4��4�o�4RB�4��4�R�4���4ӻ�4���4(��4�t�4��4���4�[�4#��4�`�4 1�4d��4���4�z�4�I�4� �4S��4��4I��4q�4��4#��4��4i�4��4%��4�W�4�h�4G��4�!�4:O�4TZ�4��4�ܽ4:��4˔�4�G�4�c�4 ��4��4�B�4�S�4
H�4�C�4'��4���4�5�4 ��4/��4���4�5�4��43E�4L��4���4���4o*�4���4���4���4O*�4m��4��4�4R��4��4j1�4�Ė45q�4�X�4�F�4���4��44�4Z޻4摱4�4���4(�4ҟ�4di�4w�4��492�4���4L�4��40��4���4ʿ�4<��4��4Z��4�4���4�u�4���4^Ѳ4�6�4��4�׹4.��4C��4��4(��4�b�4�/�4���4��4�j�4o�4p�4���4Ki�4/f�4㈾4�>�4�G�4Q��4��4`s�4��4SW�4��4Y~�4���4�L�4φ�4�X�4���4��4�4�4W��40��4��4o�4�6�4.E�4�r�4��4��4M/�4!�4Sҽ4�W�4ǰ42��4r��40��4��4�h�4Ar�46��4�n�4��4�Ͼ4	��4���4���4��4)�4��4��4�P�4y�4v��4=H�4{��4Au�4�l�4���4��4��4�r�4R��4I+�4!�4��4u�4���4�c�4���4"��4��4	�4'd�4yX�4�j�4�C�4���4��4e��4�߫4>��4��4�x�4I��42�4l��4��4��4�c�4�e�4(4�4���4���4��4�4��4��4��4��4��4���4�7�4]�4ȷ4 �4�"�4���4���42��4&�4?�4���4<x�4�|�4ٴ�4!��4 K�4e�4MS�4���4�ͼ4qi�4_�4e��4���4�Ӯ4��4T�4d�4��4��4c�4$��4���42�4�د4S��4��4��4��4�>�4��4U��4Uk�4e4�4Sh�4pl�4c��4���4��4��4�_�4��4 ��4���4}��42ƹ4�4�	�4DA�422�4ى�4�?�4�8�4�z�44|�4^ʱ4�l�4���4�N�4�j�4��4���4y�4-��4�ο4�N�4A��4��4��4��4�վ4��4G��4�F�4�5�4���4T��4��4&j�4�n�4qL�4Ê�4��4�X�43z�4>��4�H�49��4��4��4]/�4�~�4��4'��4���4v��4�4߄�4C�4���4$�4���4\4�4J��4���4Y��4���4+5�4<e�4c��4���4���4�3�4�F�4@��4^�4�(�44��4W�4dʰ4B��4��4q��4�
�4W�4��4���42��4}�4��4J��4��4��4���4�5�4���4G8�4��4�.�4��4��4��4n�4���4���4K��4��4��4RE�4=|�47b�4��4���4�&�4|��4G4�4b��4���4<��4�B�4�Y�4/a�49��4�d�4 ��40��44�۪4$��4]%�4�v�4���4g�4K'�4�n�4%��4+��4���4>.�4���4I�4w9�4	۹4�4�4�Y�4r��4���4��4 @�4�b�4���-�r-��-���-	��-��-9q�-;��-Q�-���-Vr�-%�d-ȵ�-?�t-���-���-�d�-z>�-�k�-��-�zK,=!�-��-�t�-�~`-`d-W�-���-2H�-d�-Z��,_I�,/��-��-k,�-ʊ�-Ц�-�'�-~}.-���,�Z�-SC�-u�-���-�w�-�N�-��-?8�-���-��-�s�-;M�-���-w��-�Y�-���-;�-Z �-8/�-���,���-���-*��-9R^-���-}�-?e-<�-Z[�->��-��-r��-��-gU�-���,41-�*-��-#`�-?��-_F�,>�-с�-�Z�-�1�-�y�-F�-5��,,��-w�\-|��-	��-2S�-�-�B-t��-T��-���-���-xA�-f��,�r�-���-���-�f�-���-���-j��-l�\-���-{m�-�L�-���-M�-!��-(~�-0N�-\,���-��-e��-��-���-ΐ�-I&�-��-���-�v�-LV;-�G�-R_e-
-���-���-��-q��-;��-_|�-^�a-��-��E-2��-}g�-Ra�-O�-�m�-���-��-Vb�-IA�-�L�-�a�-��-;��-GNo-�t�-���-}��-�(�-��,h_�-�q�-�>-��9-��-|��-��-
��-��-P%4,���-�l�-��-g"�-�C-J��-/c�-i6�-�f�,�f�-��-��-���-�H�-<ޒ-��-µ�-���-v{=-k��-dN�-�:�-1l�-2%-�-J��-�*�-Iz�-/0�-$�-�H�,��-t�-kE�-���-�P�-���-=��-<�,�s�-���-���-�/�-���-z�-f��-^�-Y��-�3�-҉�-�B�-��-���-���-R��-�}�-��-7x�,,�u-[KL,6�-��-�z�-x؄,�y�-�2�-m�-�J�-���-��-T��-���+���-���-l�q-���-~v~-�,�-�ũ,x��-m��-c��-[Ƀ-Y)�-�B�-���-I��-��-9��-�.�-��-�w�-���-lͥ-�G�-�R-��H-���-:�-?s,���-Z��-B$g-A	�-���-R�-�z�-���-���-O}�-,��-d+�-�r�-S��-�r�-k��,���-�A�-[�-�T�-�D�-m��-�;�-�-�Y�-&�-?��-K��-6�-5�,���-4�-�}�-ܽ�-L��-���-۰�-���-x|�-�-��-���-�~�-�)�-�r�-�-���-��-��,w!�-�cw-1J�-$�-}V�-Ֆ�-��-;5�-���-���-�9�-N��-�-(r�-\t�-���-�̡-���-z��-��-���-v�-8��-�.3,���-ӻ-o��-(@�,"h�-�-:|�-G��-!�-�+�-u�-���-tX�-���-�D�-Ui�-v��-Q��-��-«-�	�-��-��-S��-���-�D�,� -V��-�-�%Q-��-���-C�,�^�-'��-��-�`�-���-	�-���-)+�-�V�,��-��-���-u�-���-#s�-�'�-[G�-د�-�`-���-�R�,�^�-g�j-���-Ӳ�-@��-�+�M�-��-@�-ދ�-���-� 8-�%�-� -��-c��-� �-���-�u�-��-�M�--H�-�y�-��,|O�-���-�~�-n��-�G�-���-�l�-]��-���-
��+Ի�-��-���-���-���-���-q�-%S�-b�-	K�-V�-�[�,+i�-���-���-�C�,�L�-�t�-��n-��-M/�,�b�-l�-S&,�\�-�y�-���-!(�-��-w��-�P	-a�-|H�-�O�-�J-\��-���-�w�-��-��-��- b�-���-�D�-Z��-�-�@�-��-I�;-�T�-M��-��-D_-T -��-P��,2�-�s�-�F�-C��-���-<�-'=�-mWI-+��-^�-�j�-k�,�~3MG�3B/u3/�3R�y3�(3��3��3�<2�r3��3�?23��~3���3y�3�3̫h3:Y�3:nD3��G3�A?3�x3 �x3A�]3w�3PD�3�F�2�t3�$}3�Q�3{S=3��3�|~3X��3%��3X~3\":3�}3��}3�gK3iy3�/r3��3i1t3���3 B�3eY~3��{30hp33h�3ٱs3�"~3i�3n�$3�~3�m3��3^�3�s|3k��39�w3ʁ�3�v3��|3_m�3!�:3�M�3�&�3�́3#�3�V{3%�}3w�}3)M�3��y3P4y34'|3(Ry3�jz3��3���2��2+�}3���3���3��w3Ǔg2Rr�3�z3uy~3���3dw3y΀3��}3��3kx}3�3��o3�^~3̆�3f��3*�u3��s3��>3�[z3ȿ|3k��3C3'9�3�~3%�z3+d�3��3�s�3'�3ġ3Ҏ�3�~3�t3j.�343�l3d܁3@�E3I�~3��}3�v|3�*3��23��~33
z3��n3JC�3��u3��3�3�~3{�Q3=T�3�w3{3Z$�3�U3��3�ǁ3g�3r�}3��3�}3�Ky3��i3a�3�׀31��2�p�3K��3rDz3��~3��37��3��q3t�3�y�2�|3�ƃ3��3m{3<�|32�g3�d~3�M3l�3�jt3�G�3��y3'.�3�~|3% �3��n3?>�3,�}3��3�3�z�3Sp�3gK|3\!v3��a3�3N
3��	3<6|3-�3��y3W�3;�u3|F�3��3���3���3���3�s3L�~3?�~3��3��X3�q3�n}3��3�36K�3��{3�{�3b:�3}U3�[3S��2��3Gh~3y}30	�3R�}3n7�2!�|3a|�3�vo3�>x30�}3֬b3V�3�3N3m�~3�`�3��j3YI�3x��2�F}3=V-2�Z�3�Ԃ3ZJ{3��t3(��1Q�y3��|3�c3!{3ӿ�3CU@3A,�3C3)�~3�{3���3��3��3%�z3��{3��|3��k3��s3�1�3��|30Y�3S3L�s3V��3�d�3�Ԁ3@��3;�~3U�{3�m�1P�3t^|3 yH3��3�}3c�}3i�M3Da3��31�}3hJ�3�3�3��3nU3Df�2�{3�߀3��3u�2�v3�my3��3�^z3�D}3��u3�f�3^@�3��z33��1FӀ3��3#�3�D3z-3��n3�3��3�q|3�}3�3#�3Vv}3�~3��T3O�{34~3�΁3�o3�'{3��|3oix3�l�3��~3�~�3��|3t u3�Z3w�|3S�3�|3Mv}3�}3-̀3u�3��2��3�33X�3�ۂ3g~3��|3��|3�Ձ3���3��3C�3YLy33��3X�z3�!�3�E�3�v3Qd|3��|3U3��~3���3E�3���3��w3k�3j�3)Y�3ۡ�3au}3�V3�L�3��~3z�}3�A 2�?3�(�3��34�12��l3]y�3>��3N�d2�3�~�3�!|3���3y�3�т3V
~3�|3�g�34�m3��y3Ԣl2ws3��u3���33�3s�3��3ww3dwH3�ȁ3x�{3�M3��h3��3ڤ~30��3*�3�Qz3e�y3�"�2�\;3�C~3��E3�L�3*�Z3�E�3�3�`�3�R|3��}3��|3TЁ3;A3o�3��3 �w3�2l�m3¹{3��z3@Ki3LG�3�\~3��2�Z�2��}3��3כs3��~3�L�1�3�w�2]�E3$d{3��3Z�~3��o3�L�3v�}3�v�30�~3Ҕ3w�3&2�P|3M�z3Nz3%�3v_y3(I�3��3N��2G��2|��3d{3���3�pq3X}3V�}33��3924�z3��3�ȁ3�}3�y|3U�}3���3�Fs3Hz�2��3U3v�u3�gz3�:�3�b3��|3��{3�V�3X3�Hm3oz3ș3B�m3#g{3��3SH�4�P�4���4��b44��4e}4�V�4��l4-�4bD�4�)]4ac�4���46�v4�ڍ4��4}m�4�$�4�G�4��z4 sz4L�4%,�4�j�4�k�4��4��84�&\4fC�48��4��X4|��4A�4��m4�4H�4Fp4�׃4�4��
4{݋4_P�4��4���4qa�4�Ȇ40�4h�4A�4h��4)�4D��4{j�4���4��4�q�4y)�4l"�4K��4�g�4���4���4�F�4�V�4�'X4F�4&�z4Ç{4U�4��l4ί�4��4a��4�4�/�4"R�4�w4F�4lY4��4>��4��4��A4ϰ�4#Ɓ4(�4�R�4�x�4#Y�4���4�*T4��V4X��4�Մ4��4���4J[�4ʄ4*�4�d�4:�4���4O4��4���4� �49i:4���4N|~4���4���4��t4-F�4A4)�4c��4�}4!�4~�4
��4Cb^4~�4�H�4�ـ4�B�4(4���4:�4/�4��4�"�4Q�4R�4�94�3�4�4��4�x4zt4P�4�_�4��n4<�y4��4'�4�~4n�N4��4�r�4�b�4��'4D!�4��z4g��4��4z�4l}4؋4���4�#�4f�4���4��z4��4��4�7[4�ő4+�4Y#`4X4ĸw4���4�E�4]�4>J�47�4 �4���4~�4��x4��e4���4�6�4�4Mc4ʇ4U$�4��4�w�4�C�4���40�4 ��4��4�A�4���4�}4|�4g�4hm�4�Wq4���4!9�4&Đ4jt�4d��4��w4j{�4l��4���4�~4	�4w=�4�4挌4���4Ȅ4.�4֎4^��4�:�4MG�4l׌4�4L�4d0c4,4�4-M�4��4�E�4���4��4��b4-��4���4U�4��p4���4!�4�`4.�4�O�4F�4f<�4���4���4��4 ��4?�4��4��4�Rx4Ȝj4a�4[j�4Ѵ�4v|4=��4���4;��4Y64���4I�4�L84�4:�4��{4�?�4X��4��{4�K�4�{4���4���4 &�4$�4�s�4�>4��4m��4�V�4?G�4�949�4?ݏ4��4m�4<�4Y�4��4얌4C@4�֍4祝4tKr4軃4���4���4YW�4'P�4�D�4�	�4
�4�˄4i��4�i�4��4��4kX4��4eww4�Ox4 �4j�4ޥ�4=_�4?�4 H�4ˎ�4^��4��4!)�4�V�4���4N?s4�N�4Av�4޸`4�!�4�Ò4�B�4�\�4� 4�`x4v�4Qg�4Q$�4�~4WRh4�4��4�$4.r�4P)z4=;�4jN�4�V�4U��4#Ҍ4�ܔ4с4J�4|��4[)�4���4�Z~4��4��'4�O�4yn�4Xp�4�Ґ4n��4r��4J��4��w4�u�4�u�4��4S�~4��4���4%=e4���4�g�4g�4��y4�ۋ4��4+a�4^)�4�i�4�
�4���4F�4;2�3�t4��4��|4�hk4`��4h��4�;4��4�Jh4|4#��4� w44�4��4Z0�4���40J�4�-�4��4U�4�%�4ED�4)�b4�0�4�Ń4�ԋ4�?�4N�4�4R,�4�4s�4��4A!�4��30D�4��`4�Ϗ4y��4�,�4�@�4\�~4�-�4V��4��X4 y�4 #�4d��4TÈ4�Wx4Ʉ�3a�4�2�4ה�4�m�4�^�40��4!�@47��4R]4قe4��4��4{/�4%ƍ4)�4p�4�p�4���4��4`�_4ӂ4��4Ea�4۲�4"~�4(~�4�4`�4�g4�z4�U�4�Ä4���4ѵv4�ڇ4�"�4�4[��4i4���4�V|4}ȅ4g�4��4H!�4�4�c�4��4�m�4 ·4�Z�4栐4���45��4ǿ}4��t4O9�4�T�4Ȅ�4��t4.x�4�-4rЃ4��x4��j4��h4��c41@4�74�y4pz4��r4,]d4��v4��a4�4WL]4(o74�u4��:4�r4kL4��k44�r4"�T4�no4f�l4�,y4t94�W4�Xa4�q4�74>ik40yq4j�v4��p4 	A4<�x4&Nc4�i{4j�f4�n4��a4s4�u4~�v48c4�;U4!�b4�:4��m4jr4-uw4�jo4��^4��b4r>p4ɀ$4g�s4̶u4Qd4�
r4�^46tg4�zq4�o4y#Y4}cs4��n4Gi4��~4��H4�Et4��e4�$b48V4|m4�
94iu4�g|4��g4��v4�Dl4�BL4�Vm4Ju4O�k4�/m49�l4�/4��_4�Yq4G;y4%�Y4eo4�4!*r4�;4g�s4Y�m4C�y4�U=4��t4�n4��24�Yo4�qp4C84{�z4b�T47�t4�9i4Y@4�p4��o4��:4įp4��r4׶l4?�_4,�\4��[4�>u4E�Z4�(s4�;q4/04�h4,Er4��q4�6R4;0X4�`4F�s4�l4|�m4id4BE4F�d4kv4��U4�U<4��q4$�Y42Wh4�YM4�vS4�jm4�vi4D�o4�\4/�m4D�x434��{4��K4v994b?4�vl4$�u4��{4h�w4�x4ۢo4?4�y4x�=4��p4�+?40�p4�e;4n=4 �f4Ypb41e4i�$4vHz4_|X4��_4�6d4Ve4�S4��I4�{4��t4�_4��:4�=4V�u4�y@4��h4u�p4w4�_4�k4X5740�p4]zs4w4�v4_Rx4�Xf4x9p4�W[4S/p4�l4�z4�o4^R`4Aa4�ws4Q�S4��Z4U>K4�Ue4��V4�W4ʭt4�m4�xq4��|4Lw4zp4�p4�j4��b4�Qj4��d4z�p4�%n4.d4Pn4�VL4�b4\h4�i@4�L4Uc4��m4��w4'�e4�D}4�'l47�q4��n4Q�k4ؠ44��w4��]41Sn4��l4�$24��=4��t4�`s4��s4�s]4��b4�P4�/q42�s47]x4Z;t4o�z4qu4X�^4a�_4zNr4��x4��b4?gh4s4e�r4��Y4��p4�|
4U
;4t�u4�7>4�r4wsx4��h4��p4#<w42�i4��q4.x4��x4�qx4i�u4/7W4��s4��64uW'4��v4Z9F4T\4Vw46�d4�	w4.y4yd4zev4�dk4�L]4�7u4��r4�in4�0B4XJV4�
w4ߌ]4G�d4�2w4�z4>�g4~�y4�84'U4� u4��r4��54_�t4�h<4b\4BZp4=Or4��j4�s4-Ej4�ep4ð^44,4w(F4�Ox4�>84ٟ_4�vC4�Ux4%�P4��e4Rb4��u43|4hvb4��o4b&\4�u4 �d4�&94hb4kx<4�A4-C4�pu4�W4��q4 	W4#�o4(z4Z�r4�Ur4�Qt4�AZ4�A4_e4� >4��t4�|y4%�n4�r4��r42�\4�yz4$�84'{u4� c4��t4W�n4��p4�2V4)�U4�m4��74Tp4��r4ދc4�f4��n4��t4 \I4f�p4�5n4S+p4��h4NQl4V&4�yt4A�h4�9v4O�y4�{V4��`4=�s4#n4�54p�t4U�l4.�r4U@t4�u4d�B4�l4�#>4��`4��:4d&w4I�x4�U4pt4 s4Qv{4�s4@�j4��i4#Zs4��u4��q4��-4LG4�No4�:x4ۡv4y@r4�N4o4�0x4,�p4�F4EG`4L�f4��|4��:4�HP4_�4�a4L�T4�AI4�^h4�m4�jk4m�i4��m4�Wt4<jm4Grd4�v4_l4,AE4{k4�(c4��v494�(_4_p4^�k4��o4%�%4�Yq4;5%4Q)4��T4fa4��u474R4�
m4�c4P>u4s�E4>g4�@o4��s4{/r49�64Pk4�P4�(t44y4��d4�r4�R4�`4��b4F8u4+9p4��w4X_A4��k4��U4�q4�x4��j4�\�4�I�4��4�ԃ4DM�4���4z��4My�4`��4���4f�4�7�4+;�4�q�4��4�T�4�O�4Y��4S1�4>�4_ջ4�[�4{0�4��4qx�4SI�4|��4�o�4�9�4�h�4�e�41:�4�?�4���4�/�4�+�4%��4MF�4��4�g�4�ӵ4
��4��4�/�4���4�-�4���4� �4��4���4���4�4�~�4i@�4V9�4q��4:��4�}�4���4���4ul�4�2�4�"�4z��4vR�4�d�4-�4C��4�l�4��4�Ķ4��4l��4ť�4�5�4=�4m��4t��4U�44N�4a��4<�4�¿4�|�4�L�42g�4
,�4�W�4�^�4t�4a`�46"�4T1�4:��4^�4���4�U�40�4�s�4���4�.�4�O�4�F�4g��4�r�4�)�4��4�g�4Z��4o��4�[�4F��4�i�4�F�4,@�4���4q��4vK�4:�4���47��45b�4&ݹ4�S�4�4(��4fa�4�M�4�3�4�3�4 ��4V�4�L�4t��4C-�4��4�P�4� �4CJ�4kH�4���4�Q�4���4R��4�%�4w_�4�{�4��4���4�H�4���4,��4��4��4���41��4>z�4E:�4�U�4���4��4	��4���4ǚ�4���4G��4�A�4�~�4?��4���4�ֻ4W\�4,��42��4X��4�g�4*��4�ٽ4_��4J�4���4c��4���4�]�4�t�4k�4t'�4�X�43�4�$�4���4j�4U��4_.�4���4,^�4���4zذ4�)�4���4���4k��4+g�4IE�4���4
ԩ4~�4��4��4Y�4a��4�m�4���4��4qu�4�ľ4�4�H�4���4˻�4���4�4I_�4���4��4�޽4K��4W��4��4W1�4���4�B�4ʨ�4]��4�M�4���4��4!M�4���48V�4��4��4��4���4�3�4�n�4�/�4>�4��42/�4��4x�4Bڪ4���4d)�4k��4�h�4�Ž4���4��4B �4�5�4&�4�<�4��4:��4�}�4�H�4��4�I�4Vع4�v�4�	�4���4qS�4e��4f�4^�4��4Y�4�\�46��4a�4��4`��46��4���43�4�4�K�4��4↽4���4�v�4>ͼ4{��4V��4K��4x��4��4�k�4�4ϰ4��4h��43��4|Q�4���4�i�4��4�>�4���4�2�4X��4^��4�W�4�4��4���4�{�4C�4�k�4B��4��4���4���4�w�4��4I�4�f�4Q��4�<�4z��4��4:}�4�W�42ί4�8�4ٻ�4DX�4��4�F�4Ǫ�4]b�4F�4�+�4���4&��4�,�4Z��4'��4�@�4N��4���4���4��4���4���4�K�4��4Ě�4V��4���4;��4ɾ4^��4��4�g�4[��4[`�4��4�9�4 ��4���4���4g��4�!�4�,�4%�4�6�4c�4�2�4$4�4�޹42��4���4@K�4��4�`�4���4"��4�h�4�6�4��4 �4�J�4���4J��4��4W��47b�4�2�4���4���4�#�4U�4�ͷ4ɽ�4�P�4恩4��4��4>
�4t��4�{�4��4���4�,�4�֣4���4{�4��4��4�S�4ޫ�4H«4�٬4���4'A�4,�4���4��4b��4U`�4f�4䱱4\��4��4���40�4�:�4n�4��4yŸ4�i�4c��4;�4���4��4jV�4���4�n�4nV�4�Z�4�[�4���4W��4��4_0�4ڝ�4���4���4�m�4���4W�4d��4���4#�4�*�4j�4ZS�4b��4�W�4Ū43p�4(&�4�+�4tC�4���4�!�4K߽4 �4	�4��4e��4T@�4g��4�u�4�4MW�4ճ�4A��4�$�4د�4x��48�4F�4^��4���4��4�I"555�25�[.55,5��>5�,&5/.5�975f�/5��35��55Uu25f�47-5�5)545�35Z�55N�+5��/5%�05�]+5<?(5|l.5�i:5�-95�XC5z�15�y-5�E5��=5d05���4D�>5�85(�35��*5�265�(5�#5#�15��=5w�(5~XA5a�=5Rh/5R_25.�'5��%5�p�4ި&5I?/5]?/5�?5Q�85��-5�,5�p+5�W'5)E5�335�95��)5��75AL95��&515{25�,5�f35�~65-	65!/5�a/5w;5��65$l*5:�65XD5��.5>�/5�>5�W@5p@5�E5V1>5V�?5��-5DW;5�}45
�45F�15M�*5m;5�-5ԯ?50+*5`N35e�;5_�.5��95.^.5/�;5�05��@5�C5s�/5�GC5�m"5��15�85xA@5�m)5�Z;5�.5��-5�.5�+5��)5̸>54�05�J05�
95�n15��-5�F5Ql15E15��+5@0-5��!5-�25ӠD5T�$5�05�75�s65�q 5��55�15�=5��05�'45�35I95��B5^0)5]<5�/45k�%5��35��45P"5&< 5�e<5��$5��5L�752 >5��'5�O15�y45��85޲/5��25?-5�<5�C5�/5r�I5��:5,}85k�/5w+-5=�45�05�+5��$5;95b�35��55��@5�15�L>5�N5R:5�)5%k65��.5�l45��=5�9552#5�!25P�65g�251L<50FD57D*5x*5�.5C_15 �=5'�>5V�(5�G15�2(5z
456p)5�D45�<25��'5�55�?+5��05�}@5b�'5��A5�65�k%5�]5b�95��.5�A;5�.5��35,�95�=-5�w'5z75��15��-5۬,5�)*5X(5�;5��:5uC45�s35��45��.5q�45"R75M_C5�-5�,5��=5P�65�05w�;5B�525mm35�5C5@p?5�.56�:5I�G5�15z_55eo457�05-ID5ݝ*5X�25Th85+e95�,35��:5��65z�5��15�-"5��@5Ɗ-5�(05��5S`65.o5��15�75�,:5$765��65XM45��5�75 �5�SI5�:5��85G+5;z>5�O55JU&5��25��>5
�&5��,5Ek25'u4551�?5=35t�05Z�15%�=5��05҆@5`J(5��252+45��35�<5t75o=5��=5475��>5f8?5�:5��65UA75��)5�>5RX?5w[<5�45�1 5�65lG5�q45&�15��058h/5�Z.5�c75�N65��45	�(5y?5��(5�255>45l35��45P<D5��15rz85=.5#.5�<5*r452�85�25:�:5�D25[85�65��,5F�85[�/5v.:5�e95�75�55`25��5�25b�@5�<5��45�(,5ެ,5d�/5Fh55W{15��85k#5�k25�".5$�75��-5�15.d#5@++5I=5Hj-5�35��:5 D35�4545nF05e�)5w�35J�25�45�j*5��15�)<5��$5�"=5�45��15@=5HV45�y15�!5ɣ5m�C5�45�1656h%5�H@5�#/5�*5O@:5p�65�-5�25ڏ5a�45V�95��&5�v25�j85��:5ˊ5
�05Z65D�75G�;5�#5�35Np5��55C<5�|25z.-5��<5�d$5�2.5��?5�.@5��95s�:5I95L 5':#5I�,5� 35^q15��=5��5+h"5��75��!5�(A5��,5�105�F�4Dm)5ǉ(5�15b?5�45�5�s15N75�-5��05��$5g�?5"5"f 5Ӷ/5щ55ǜ:5�45]�05|#*5��*5Y�45xc;5&�:5,15Ge95m25��45��*5�(5.�253]&5};>5ͩ$5��15h�45��;5㬬3+�3�r�3�?�3~��3'�3Z��3���3��3��3r�3��3D�3:�3R͐3�g�3��3�+�3m)�3U�39J�3��3���3���3��3EI4^@�3\��3
��3J�n3���3Dr�3V	�3�8�3�}q3r�3���3"#�3{[�3�c�3t��3q��3�y�3���3^��3��3���3p�3MW�3���3F�3+�3&C�3�F�3E��3)�n3"��3�N�3���3O��39|�3���3���3��3;��3~ �3���3��3�
�3D�3�#�3a��3��3˱�3��3q��3���3U�3pI�3_�3m�3�@�3+y�3��3��3���3g�3��?3�3�3^
�3L��3���3~
�3�g�3�c�3O�m3<?�3y�3Nd�3o/�3��3���3�u�3�3�3��3��3F�3���3Gi�3��3��3Ԋ�3���3��3���3ґ�3�~�3;�3���3���3Ǫ�3���3K��3���3#3�3���3O�3A�3b��3�a�3���3%a�3�n�3aK�3�Q�3��3q^�3���3��3�|3���3���3�T�3�{�3���3��38��3��3O��3?Q�3��3��T3���3��3���3�f�3j��3��3@�38��3O\�3~Z�3G4�3G��3SV�3��3>��3�'�3�A}3���3���3^V�3�6�3C��3��3
��3G��3B�3�Q�3��3�K�3L�3|��3"��3Y��3�K�3���3U��3JX�3���3��3{
�3V:�3�ћ3���3���3ba�3��3��3���3@%�3�!�3���3�B�3r�3�A�3}C�3�(4Z��3���3���3�a�3x��3���3���3E�3���3���3���3�C4��3�.�3�O�32!�3��3Ӑ�3xx�3[��3,�3��3���3��4�Z�3d��3z��3+*�3I�3� 4�_�3��32��3p��3�p�3��3�&�3���3���3���3��33T�3���3s�31��3�3���3tg�3N�3
N�3K�3��3���3�s�3�w�3@B�3N��3�T�3���3
\�3Ly�3W�3�g�3���3���3��3���3Y*�3���3�L�3$��3>�3O]�3�\�3))�3GI�3a��3�U�3h1�3:�3T��3��3HN�3��3Ʃ�3��3��3���3�s�3~��3��3\e�3�(�39#�3�\�3���3VW�3���3���3@��3%��3���3(��3�\�3���37��363�3��3}�3�L�3��3���3޿�3}_�3�	�3� 4�I�3��3*��34#�3���3�>�3�7�3<��3��34�3/�3�B�3g��3���3�#�3��3�.�3 ^�3�B�3��3�ö3@��3���3���3���3��3���3�3��3A��3:�3��3%��3���3O��3Zj�3���3o��30�3X�3�{�3Jc�3���3e�3�$�3��3� �3S��3A�3���3QC�3�6�3��3F��3p{�3e��3ٕ�3N%�3�R�3��3�S�3���3���3���3B��3�0�3%��3*�35��3��3��32��3��3��3Չ�3
��3���3>�3@��3�d�3J��3���3���3��3���35ڝ3�I�3{��3`<�3���3���393�3���3���3���3�[�37��3V"�3�,�3���3i��3��3���2�V�3Q�3�3x�3���3��3�V�3,��3�4��3���3���3��3S4�3Ԁ�3I��3#��3���3��3��3[��3���3�G�3i �36��3�>�3tt�3	e�3��3M��3��3��36��3���3�n�3YM�3� 4|��3��3�3�3'�3��3���3���3.�3�3i�3)��3���3���3�x�3L��3S��3([�3�y3� �3=��3:|�3���3���3��3��3��3h�3ĕ�3���3�%�3]�3z��3Ea 4��3Q#�3���3�*���)�*�0�*�k�*�.�*YO�*��9*��w*�/�*��*Z�*)�*7�*u5�*5��*�ՙ*+�*(�*�%�*U2�*�U*��c*�#*`�Z*ܺt*n^�*�r�*i,�*f��*�!�*��*@F*uY*!�*�E*�	h*$�*3��*A)�*�i�*�b�*��*�$�*���*���*w�A*4�*s�>*�.�*�L�*s*	��*_L{*�*�l�*&k�*NH�*+ �*^��*�sb*?�*��*�I=*T�B*3�*EWH*e�S*g�*X�*�Ll*'��*���*��*h�S*v2*Y��*kb*}�*�a*+��*�NL*�0�*6�I*��*
�B*Щ{*G�*�Gd**��h*,��*�ϕ*��[*���*��*x�l*pL�*F-�*SƔ*z�>*�J�*L�~*�Ԙ*_Y�*��*\Ò*䗎*��[*���*��k*�l*�/n*���*#��*@v�*�<*?R�*��*t�/*�d*�B*Td�*�1�*č*`Dl*��*{/�*J�*�i*���*��*_�^*8�w*0�*���*^I�*l�*�P�*�_*N��*i,�* �f* YH*��_*�*~S�*s��*'��*$�l*�7*�;�*_ߗ*�{�*���*_�W*�y�*���*?Uu*�T*�ϕ*�s�*^�*��T*�1�*E�o*�ے*��e*�ؑ*Ԅ�*���*H��*䒔*&S�*�*�'�*�̍*�X|*hz|*��&*�g*��u*�O�*U�*&�*5k�*!�A*��*o*yZ,*$l*z8�*�
o*�z�**�F*���*%&N*��B*��*fΕ*��*��e*��e*��h*َ*B�Z*g/p*�w�*V��*�d`*B�z*�;�*�Ez*[�*_�*���**M"*��*|�p*/'�*	�*�"�*��*�ix*l2�*)�*��X*.~�*$��*�i#*N��*,[�*���*�˕*\�~*�E}*��*�-�*��	*�(�*�O*,2�*DS�)��*σ�*�`<*�#�*VnZ*Q=8*0c*�Cy*zmc*�;�*M�a*��Z*s\F*��V*��*
Ă*Y�*��*���*���*��L*rp*���*�V*��J*�T�*�hv*�K�*�0�*-h�*�[P*�Q*��*1F2*rG�*K:9*���*Q�*M�a*n�*��c*Ú�*h�*��*3�~*Ᲊ*Wߙ*��S*M6Q*�Е*�y*�y*8i�*�n�*1�*vʊ*,S*��*�}�*앛*�x�*�(�*,ߍ*#ņ*�ԋ*�4�*��*(5�*5C�*	 l*_@*�O*��*vaq*���*�N�*ܹ�*��s*�*|�*s�*�1*�R�*�/�*[�*0C�*�,O*�9�*� �*5%i*[�l*ﱟ*ۦ�*(��*�'U*���*���*F�e*U��*ȃ&*�=**I�*	 **���*�6�*�͞*}�&*[4�*;k2*l��*�w�*�X�*@3�*Lv*��*�	|*X��*DO}*�*
H*�	a*�*�	`*|r�*R�*:�*Y(`* �*�t=*�Q�*�|*�6�*.E�*A�*S��*�8�*#q*�)�*b��*��*�*ʍ*��*�})*z��*p�*xA*�'{*뭜*��*�9�*�i�*>��*WI�*�Wb*��*5�*�o�*I��*Qo�* �*-C�*FO�*�G�*6�*p�_*E�*�i*ֶ�*1�m*��y*�;�)�*b��*Wa%*�X*9W{*�1�*�R�*�A�*��)��q*�*��t*��*�e*��*��*�7R*�9�*e�X*"\*�lP*j�*���*qkj*�`�*�Zh*�w*[\�* w\*�c�*z�o*P �*nl*�˜*�*&�*�,^*��h*/L�*r5�*�]�*U�*#~�* ��*Gԛ**�*��*��*w��*��*��B*Qw�*��*�K�*���*��*�<�*�߈*	њ*� y*ٹ{*�H�*2�*^*vHd*�s*@��*��(*$�*��*��a*XD�*1r�*7��*��*_��**�u*xݙ*��*��*�mU*a�*��*�d�*�r�*���4�q�4$q�4�z�4A-�4/�4N	�4s}�4A��4~�4���4+
�4*��4�*�4'��4EM�4�^�4�j�4���4e��4"��4K��4�7�4�*�4.��4L��4��4�o�4��4��4���4�m�4A�4L��4�o�4G��4�H�4���4���4�?�4+��4���4�J�46�4�4�G�4�4 k�4�T�4�T�4i��4d��4��4)B�4���4~]�4��4*�4��4P��4�+�4p��4�e�4�J�4E �4���4�]�4���4Oo�4}��4#J�4�a�4���4w5�4���40��4q�4^N�4�>�4�i�4r�4
�4^n�4���4Ջ�4q��4M��46��4���4��4s:�4��4"3�4Y��4Kx�4�4���4���4l��4,)�47��4���4��4w"�4��4"5�4�L�4Z��4���4? �40p�4�y�4���4a�4�U�4�.�4<�4���4��4���4��4\�4ʾ�4�4�4�N�4�_�4�^�43�4���4��4�u�4}�4C`�4���4�'�4 ��4���4��4�_�4d1�4���4L4�4	��4��4J�4�z�4�$�4�x�4�[�4��4(y�4G�4	��4���47��41��4�ʼ4x�4\^�4c��4���4]q�4Z��4�4��4?�4��4���4]��4���4#��4�F�4K��4���4!��4o:�4
��4d�4��4�'�4�`�4��43t�4���4:Y�4F��4Ԃ�4���4���4[��4���4��4���4;��4���4���4�:�4���4o��4�}�4�^�4�f�47�4ք�4 ��4���4�V�4���4C��4j+�4�=�4���4r��4?+�4]	�4�X�4���4w�4���4�4���4\t�4���4LY�4���4%E�4(��4�(�4xH�4�4���4��4��4@�4���4�K�4���4<�4���4б�4�2�4Ж�4~�4L��4r��4j��4_�4D�4���41�4���4e��4�B�4r(�4*V�4��4�S�4P��4G��4D��4z�4�Y�4���4N�4*��4]�4��4o��4 ��4���4�%�4s�4Y��4s"�4y}�4���4�#�4n�4��4\��4�4���4�B�4:E�4͔�4�4t;�4/w�4��4�1�4�.�4��4�"�4��4���4��4���4˫�4���4~�4���4K?�4���4���4�i�4��4�.�4��4���4A�4O��4���4��46�4���4�v�4%�4[k�4Nb�4��4��4$��4���4y}�4�˦4{V�4�(�4���4��4�1�4uJ�4B�4�;�4��4!@�4�d�4Il�4���4q<�4U��4F[�4�P�4�|�4�-�4�c�4��48��4>Z�4 Q�4�-�4Q�4LF�4q��4�q�4�]�4A��4���4-U�4��4���4x��4ł�4���4Ab�4c!�4�E�4���4@ʴ4O��4!+�4N?�43�4�b�4إ�4���4ً�4�j�4��4=0�4��4�-�4&�4��4Wc�4,�4���4}�4���4��4F�4��4;��4��4���4_W�4���4p��4$��4G��4�}�4O/�4���4��4\�4j��4ym�4l��4���4G��4�*�4���4��4��4���4d*�4[��4���49;�4e�4�j�4���4���4�c�4L�4�4�4���44��4���4���4i��4���4=��4pI�4m��4"��4i��4U��4�Z�4��4.�4���4ij�40�4$J�4�p�4�J�4]S�4f��4�:�4�@�40�45��4���4���4���4�t�4���4#��4�W�4$ �4��4R��4��4��4!�4��4Z��4���4���4.��4��4�=�4�J�4���4.��4i�4�X�4�N�4���4%�4���4��48��4C8�4��4��4���4m�4-��4D��4)�4x)�4=w�4���4>X�4/��4W�4iE�4L��4���4�15�C95�95nNH5^�=5N�D5��)5�'J575�H5��F5��75��)5;J;5O�:5c)?5}�<5��<5��5/e45�nH5��E5:b75�25��Q5�15�t55��=5O�C5�8,5�U 5ТH5��@5�;5�0.5H�95^�=5�@5��C5��,5��;5G�15�IT5Ș+5Ez:5�w@5��?5i�;5nB5��@5��I5��=5��25�A5�>5��@5B�?5�6@5
j@5}x>5e�B5cb65�C5)q05�<5��B5�P45~>5J95��>52�-5��R5��5�A5]1K5'�N5B�955b55�^:5��F5�W,5L�65׷65!�<5�85ox<5�!35�	*5��M5MJ-50�"5Ĉ45J�@5�:5�5G5�.53	<5�0>5�0E5�)5U=5w�95p�?5�SD5��>5��65]@5&:;5��'5$�J5�G5��B5K*75=�?5@�@5��*5W�J5��15��A53%5�B5^i<5f�/5�H<5\B?5�^K5��K5.�?57)55z!95�\95�R<5�)'5�G5�_C5�RE5��;5߀?5�KA5��=5�?5=�%5��D5ħA5d�-5�}H5�}A5@�@5�II5�A)5�p95�A5-"65!15�5�:5*�%5-�:5�J5`1G5�t451?5(�E5-�.5O�)5HC5H�05a�X5L.@5.:5 �:5`N@5��55=�@5ϋ,5Pg75�|P5��15x�P5e�-5H�<5�E5n5@5��;5�uB5�>5W�55�05J�S5{bF5s�75im=5/�<5��G55�D5�55~?5�;5�;5��I5tI@5��H5'8I5�V75�W65(:5[J5"95��<5.�?5�I5�>5D�H5ä.5[I6595�05�45CA5��?5J(5 >5�/5s,E5�{;5�W05�6R5��<5q�/5{m65�/5=5�*5?�>5�45��85�U25�!5u$H5��25?�;5��:57�A5�(?5]�,5!95�[45f�75�(5
B5�U$5iXB5��*5W�75yi05�&25iRF5�3-5�95fz$5�w<5��5�/5��'5�J95�55��H5I�A5{�E5�)M5��85wr(5��:5�55FB5�05
55�k75;?5��<5y�65��=5�	55p�K5�CI5�]*5fs85y�&5'r@5�95 �E5�;59B@5�+25��B5�95�65�85�nC5/�E5�65IA05�35��5�055z65!�.5C5�,G5^�!5�F5�n>5��N5r 95I?5��G5d:5]�05(`I5X�=5zA5|"65�%35A�95[�45>�L5:] 5��=5(o?5��@5�$5D�@5�@,5*�'5OI5�F5x3I5B�@5��@5�6-5�K35��B55�@5��U5�5��)5]:5��;5:5C�+5�X35>7C5��#5T�*5�SP5H75�a45�55��C5�15]H5%�85�05�.5��55jB35&�O5��75�V75�85�^D5�4D5�r?5�X/5	�N5�)>5�"A5�25Po65wBA5�_D5��55�35��O5�S-5h�-5AbB5X"5�o:5ԉ@5>O=5��K5��>5ZU$5�C5L�A5�8!5J�D5��-5��85w�<5yB5U/5�{05L)5j�45��5?�:555�>5� =5��45j55Y|;5K�E56�*5	x@5��A5F�N5535��@5I�>5�|C5/�:5z}95�735q�55׸05$�/5!�25��95tQB5_�=5�U,5��@5�PD5��$5=�75Δ85F�/5��+5�tB5�2$5ғE5H!:5�*5Z025��=5խA5��?5�X53�B5Y�35�EC595e�35>%5��=5`95�m!5!a?5�s95��B5�5�'5��<5��G5FL85��E5�#J5�m=5ų75�F5��5l<5$�35��75�)@5�-5��:5Y(5��25c5;�95��95�65��65�.5H�@5��<5zE5�(5m:5��25�E5I�15	";5q!P5�*5l�#5\5��85�52%5�:5D-57!5$.5�5��&5΅51=5��"5��5�F 5��+5`�'5�d5�E%5N%(5�C"5c;#5#5;�.5Le5��5^�,52�25F'5G�.5��545I�5#��4~�(5e !5d�5��5� #5�j#5�[50�$5&5�&5%@,5�K-5C�5I�5w�5Ɠ+58 '5�
(56*5$I#5��%5%�*5f�5R'5g�"5�� 5�$5�D5��05_�'5�.5*�5�Z$5615�x!5Z#(5�(5O$5ِ5<O-5<"5�\!5w%'5�#5ӱ05}S)5��5�5zS+5)L*5� 5��5��35��5n+ 5vY&5885�6"5��05��#5�f!5s�(5�$5s*#5L�'5 �15h}$5C�&5�5��$5��%5@5�*)5� 5\ 5�T5XR57�5� 5v5�($5R�"5� 5��5��!5O�"5Q	5�. 5a5&&5s{"5l)5�{'5�U)5� (5j�5�.5�x'5�D'5`v%5��-5�'537!5K�.5G�5^&5w�+5�(5�� 5�s5y� 5��5�V)5U�'5fA"5�J5��5��5��#5r;(5��"5|�55'15p�56�(5�5"5�5�z5�N+5�0%5�%52�#5��"5޶5,�!5CC*5Ō5�,5��5/)5�)5p�5�C5��5P$5*�51�5��"5�25d�*5vS5��56�5f>5<c5Ǎ5/2%5�"5��5�S5 &5�5ͅ5fi,5SU�4��)5�%5��5#� 5_$5>�)5$5<T 5h�)5�7&5�m5�"5%�"5�5�r5�)5�*5�&5"'52�35W&5�(5MG5��5�-5�_'52�-54Q(5.}$5b�(5�I/5F�.5^�5x�,5�h%58b*5|5HG,5�5i5W�'5�*5L�5Պ$5RT#5��5��(5�I5�I5z�5�%5#$5F�,5�A,5h�5>�5�P54
#5T� 5��25�1"5K� 5^5��&5^�&5Q'5a 5ϭ$5޶/5ɖ'5.k5��5Q�.5��5��5s|%5i85��+51�5��5�=$5��35�!$5r%5��#5�i-5J�"5q�/5� 5�'5��%5@�5-�"5�45~^5�^#5q�5��+5��"5MO+5�|#5e�-5s!5=�5�3�4
>$5� 5�"5ar"5b$5��5�X5�{#5�(5w&5�"5f�%5�k5��"5z_$5�T5��!5��$5�V+5�~5�F5�%%5f5��-5H 5Π+5�.'5j-5�5a�5 �)5y35�k"5]85Є5 �5��.5��-5r=5��5V25Wy(5X5�l'5*H5$�%5�P"5$$5$"5�(5�(5B�'5�\ 5��5�05&�5I0*5G�+5,�51{%5�5a5��*5�x5	5�{5�4,5�25Ko#5�#5P�55��5ss*5;�%5��5��5Ec5Z�-5��5&�5�'5o'5��15��&5n`&525z�5��5Lg&5�)05Ҳ5�.35]!5$�%5��5D=5�Z)5�)-5�.(5�o 5s�$5D�5*�%5T2#5�3)5��5I�5n#5r05�R5��#5e�5�5 5�"5�M 5��5�Z'5�K-5�Y5؃5\�5�&	5�n5�&55Y@55Ʃ5{�5�%.5b�*5��)5,�5��5��"5�Y*5b"5��5
�)5ї#5R�+5K�$5�5ag5�5(S%5�/%5^�%5��5J5�#5�#5H+5�)5�G"5��5"v&5BZ'5x�5�D!5�5
� 5L5��%5#%5�5b�5��5��!5�� 5Ɣ5�5�r!5<5�s 5v\%5#5D5��5�S5Y05(5ư 5��.5��5��*5 *5�+"5g�,5]�,5 �&5��,5{�'5�%5�L�4�94D4��:4϶�3�m.4FN4.v74��<4�`?4E448:<4��54?��3�>4]� 4�A543k	4{C4[�+4�B4rcG4[43�54��,4̱84��24O�4�VC4?�>4�C74.>4�cB4 �464T�:4I;4J�94h@4�*4�tA4�.4��44�:4�H@4K�4�I74o4B4(4v�74"
>484K:4/�E4L�54&4��74��74R�;4f,34+�44�X@4�:4�"24&�94Ol74��=4��)4��64_N;4��64A3?4��<4�,64g�84x� 4X]�3t<42�94`�:4��14�64,��3��:4~24^�?4��34��=4�54��64�B84�"@4�n14 �,4� 54N1944�@4�4#�=4�*F4ҕ:4G.C4N�54��<4�mD4�54��:4P�64��64�s94�N64'4�r
4��=4��3~c;4ں84�:4�zA4rO643I54.�74�74|�;4

>4K&'4/�148^44�C4�94�84B�84��;4��74�a44��4�N
4Y94��74�14��;4U�34]�04��34l�<4J�84}�<4�h.4J�%4�w$46�E4<4&JA4?�;4|9-4�=4�h94�f;4K=44u=4�g<4�/44ts:4��54��74�z64^�4;q@4٫A4.�<4�4NA84:g&4mEI434պ>4��64�34/:4�=4ƽ:4��4�64�Q?4&�:4��4�64HQ44�84�C94��;4�4=4�B4��4�k84ۉ.4G944/��3,74 �;4p<4�F4�f74a�94jO:4�D+4v44e(54��34^�34�q<4��84e|4P!4p'64��84��=4�84E�74�<4c�24�44��84p�94�44p�@4ɇ)4�<:4�5<4e�74r�,4��24��?4�^4:�:4$�B4��,4GC54S�>4Ұ54�674g>4m	64��=4U�+4۔4�(=4��04�u@4�=4�4� 4��14'>4�=4�54:�%4B
>4�%74��64)A4B�94�=4�N74�RC4��<4�:4OjC4�84�84�$<4��>4aE>4h[4��4��<4i
A4�y@4K�;4��84�d24 ;4 �94�<4 �74KN84�&4)�:4��=4��"44�74�
41�&4�j74x�4�A4�4L$:4��E4��=4�44�54r�74M�:4��;4�264��:4�B=4s>>4�@<4J[84�(84�@.4O6;4Ń84,�454��94��B4-�3��<4�074r�<4`bC4h84��;4�I74��84!44p��3�a�3`�64�A4Wg4�')4�i74�-4&�4V�54�'4}�?4�-4v	4��84�V;4��?4��44��4�m44�z/4��	4�t4�>4�^;4�)?4n+4�N84�<4@�@4v�24�94�)<4R�!4�84�I4b�<4�@4>v64�r14H�24K434��34>%54�;49"74,�54g:4��64	 A4T�=4J/4:	;4��>4�$=4�,94�O=4C�24�54<4�A4�`44�84�34��;4�4�o%43�04�?4N�4�4��94�y,4��?4{4��,4W�=4��;4ˏ34�-F4�]24
64��4�;4��4��?4p*64@>4�Q<4�A:4"34�:4LR;4x��3];4�K-4�"+4�(4��84{�645>4&%-4@�*4e�4�94�T4��54� 4
�64��24�m;4�84�x<4*R4�+42�54��4H�94�74CU94�a<4�>4,94��@4�549�=4;h84
_4�^64uD 4,M74lT	4�BC4�54�34�=8454��-4��47@ 4ض4�:45A�3�\	4S�24>S=4�^;4�824<4�+=4?�3�{4��>4?V;4}�4�74�64��44�*64�v)4�\)4�84[<4
?4=4-j54�;4:L64�+74b@4?64q?�2'`�2bm�2���2�-�2j�D2+�2~]�2(Q�2�Y2q�w2�ߜ2~72oc�2�1v2hߥ2S��2���2P�?2B#�2a�`2� �2
�2@0v2�Ú2���2H0k2Ɍ2���2:�s2���2H6j2�U�2D�p2�012�i�2��`2�V2�I�2|4h2�DC2�2��+2�2�؝2���2h�j2 �o2u��2�{x2{�u25�Q2C�W2ݲ�2�q�2�2��2p-s2��2��2u�2�e�2wk�2�އ27͌2�(G2�̀2n�32j��2؆2�}2{��2���2/�r2�3�2q2eY�2�k�2�Ƕ2m��2�l2"�l2	}29�2~��2���2��g2�g�2K�2�q#2C�2��u2��A2�H�2��G2dg2~�k2=�2	<2Pg2B{�2S�2�;2�F*2���2N�e2u�j2o�q2KLb2
�@2-\}2�2�#�2<��1Ns2��2���2���20�2}�M2;��2�ȏ27?�2iv�2J�2^2K��2��d2�L�2볌2��_2c�A2��)23n{2|��22�2Ո�2�]Y2�ı2�O2}�$2��2�j2zȓ2��2M�n2 �u2�$2�z�2&�2�2�Sr2���2��2�ù2F�2EI�2Fw�2��2$�2�-2+A�2JU2��2�k2Lrn2�2���2�ט2��2�׳2��~2 �t2���2��2���2��22j�23mY2]Q�2m8e23I�2�Ym2�`~2�̟2B��2��W2��K2-P�2&}�2x��2��2=m2mn2:�d2���2] }2��r2�.�2�wv2���2鉣2v�2�Z�2�q]2 ?E2�YK2(&Q2�P�2+k�2�{)21gZ2���2���2?2$�i2���2�=92���21�o2kUk2�u2��c2S}}2~!�2�K$2Fzz2�52�[�2�ʬ2��R2�X�2{e�2B�t2C�2݄2�h2��\2o��2�s�2�j02��26�m2Ji*2@Ձ2x�2i2e�\2Z6�2�;�2c�:2��~2s�2�R2�h�23M2�M&2�j�2�;�2k��2[�]28J�2ɽn2Z�2a2n�}2KX2ߦ�2[Z/2d�2{V2���2��2�27�62�T2�2��p2o2�	&2w�]2.�U2�њ2��n2���2�)]2��2�[2`�c2�G2��k2�O2p�2ۉe2v�)2��P2Ӭ�2���2MK2�12OS�2D�s2�h�2`72�:�2hс2�s�2��}2��2�.�2O��2Md2,jI2��%2���2�9{2J�)2旁2��2�`A2�B�2��|2A2��C20�R2��O2sS82R��2k��2�M�2\�s2e:�2�;�2��J2d,x2�[2�q3��/2��]2�mG2�J=2f�d2��52w[L2�]�2��}2aw�2�L2��2�Jr2sll2X>y2��d2oY�28�2+=2�.2̩P2M1}2ML�2}��2�m�2.*2ٟ2uE2�2�2�Ж2п�2x��2��o2��2FmU2��2��2Qv2B�|2{�i2�P2@ -2P�623��2vҠ2���25(B2(�i2�ub2�t�2��82J�i2r^2���2o�|2�4m2�h�2u�2�~d2͵K2.��2�M�2�u2�+2�x72��U2��2��2�r�2F�!2D2�g]2J��2�2���2���2Wf2���2̭+2��22*�b2A�2���2�G�2=62	h<2q�|2p��2�2g��2F�2K��2��f2�#2k�v2��F2'�f2��w2��92�vj2�C�2�Lg2*6f2J��2�Z2��n2�2}�2�2E�2�M2]d2S�2k�N2��2S-�2nl�2	��2 ]�2�I;2���2�bu2$b�2Y�2��E2k!V2,��2�n@2��52%H62�L2./�2�n�23+�2�T�2}Bi2f��2W
�2�Q2�H�2(��2�y�2 P2��R2`�2]�~2m4�2��T2s�H2��y2�(c2u��2�d	2�UQ2��2��2ф�2�4�2'�2I�l2��2�I�2� �28uE4n�@4p@4�t?4�94�:4P54��F41�@4P�%4m�:4\C4?;4�?4�	84��E4�A@4�nA4�i
4�I.4�?4�bG4��C4�1941�B4�:C4��#4\�?4��=4��94UNA4J�64�B4E;4��4=-4_�C4 xF4�J@4�WD4��:4��?4*�B4�B4+YA4�E4� J4�>4�B4�4y�:4A4b/4!�@4��:4m$4�1F4|QB4��C4=C4��D4�D4�HH4+�94u�A4�aD4� H4T�@4n�F4	>4�4�G4�6(4!-04wU>4�5-4�04`�,4Q�>4X�A4��A4\�4�V94��?4��84��;4��@4F�B4�84�B4:�A4:�A4��@4R[D4tpC4,4�}B4_�D4�gD4�ZI4C4G�=4�TB4Z]>4J.A4��4�4�BA4��C4k�B4o]F4Yo?44�B4V�@4��A4;�;4Jg24�%B4��;4�{<4w�B4�?4:]B4f64P�A4�P=4�!E4�2G4E�94�@4t,4&{94�@4F|H4��B4�UI4�z94�CK4�K4��:4:FB4��>4:�H4��C4ǯ=4+�B40�/4y94�cF4�K@4'�<4��,4ω@4�>4PQ<4��A4�D4*�@4_�H4�J<4�D4U�D4��E4��C4;�?4��B4�=4�?4��E4̵B4~�G4w]F4L�&4lNA4C,C4��E4��>4�p:4��(4B4�!4hG=4�-4>?4�n:4�4%�84�<4_4~zD4b]>4�384��@4ЌG4�;"4`�>4�C4*�4f�B4"z�3��B4�WD4$�;4hq=4�94$;4�K4`>=45�<4<�B4{B4��G4��D4&�?4 4==4yE4m�A4�G34}Z14�cI4k�>4�H4�54ʿ:4<�@4�=>4� F4��E4v�4��E4՜4�%=4�>4��H4�#<4�d94%G4�=4�A4z14�PJ4ҿC43;4	}J4�C4R84 �94��A4u�B41�24��&43�@4ay;4�D4'�>4�?4�K4*�,46�4߼54�`G4+G4��?4��74t�?4n�@4�K4�$B4�]G4��4 IH4	E4��54�$ 4�:4�LA4��F4yr>4��;4�]K42
C4��F4��B4�m
4!\>4�C4��E4M�54?g?4��F4�84*>;4LG?4��4��F4`i:4e%D4��?4Y�>4��A4�K4F�F4�:4�&�3ԺB4�J?4g94(#4��=4ҕG4�NE4�d<4Ϫ?4�\=4�=H4��84�I4�F4,�:4�� 4��94~X=4:E4��B4�rE4�fA4H�74]�24�SG4�94y�:4�k:41�4ݳ+4RA4܉E4�r;4@_E4��74_74�K=4I�?4��?4�UA4�@C4�84^�C4�E4AH4�d&4�Q/4�w4b�4��>4Hh34MH47�74�B:4��C49�D4�JG4�U>4JI4V�-4�f:4�K4��C4R�C4t%4�T@4*kC4H�84�246*'4	�?4&s@4�`F4�*4z�?4��4knF40�G4E�E4�+4��>4�B4�;L4t�=4B!C4�B4�P94�:4^DD4m�B4b�'4�=4�TC4 �<4g�B4�?4V�A4��G4��4�84�64+";4�A4H}H4WB4P�D4R�4(N4 �=4 �=4�HH4�C4�6F4��84�/@4��;4 �=4�3C4)WA4��:4�l74�B<4.�?4��;4�@4~�;43�I4.14�2A4}@4sH4�=4��@4�C<414�EA4�5D46>4��84&C4 I4�842�4��4J4�>4��:4��:4D�F4U�94��B4+~<4�yI4�?4�@;49�
4(o@4�;4=�C4P$@4TC4)�?4�F4y�>4�@4Ŏ:4ҎL4�:94��!4gQ84�
4J�@4O�D43�;4%�4�P74	�4�74�Z�3� A4�N;4��D4��94rz?4�74,$G4
�;4�?4��C4��G4�>B4�s?4�I4�&H4
�F4YC}'hF�'�r'l_�'��'��'�W�'���'�?�'���'�`�'�g&���'�c�'Cݕ'd^'n��'	x�'3�':�'�#�'�*'㼕'<��&qۚ'�,�';��'�3�'�&�'��&Wؑ']_'%Œ'�i}'��'�ʔ'�b'<�'�ǌ'�V
'��'6ϗ'��E'�W�'9]�'�I�'(��&�1�'��'̆�'���'��<'�܍'�Ɍ'��'ŋ�%�y�'(ӗ'2�'�Ř'��$'|K�'��e&���&�,�'�>�'.r�'�u�'�S2'C��'6�'Z>�&�P'��'��'�x�'��;'5�p't�'��'�T�'f.�'.�K'���'^��'�0�'nM'˾}'�'y�'w8C'°�'�v�'���'���'u�&�'�4S'��'}�&�f�'�r'�b'��G&�Ӏ'$�'t�K'誒&B�']7�'x��'{�'T�''���'��'��'8�'/0�&UD�']��'�l'�@g'��&>V�'Ɗ�'cp�'f�&F�Y' ��'BS'8/�'�&�^�'���&�ǜ'Y�i'��'���'��'R�'hvl'녙'�m�'#�&V(�'F�V'V'j�'�Õ'%'�&�Y'�	�'p��'�|�'���'�'���'	�'y�'�@'$�8'/�'���&��'���'�k'5��&}�~'y�'n��'w�'���'Pr�'zŅ&��'�'+ �'���'b6�'�Ģ'�c6'[�'ᄁ&�E�'2��&Kې'Q��'Y�'��'w+�'�')s'淍'"�&$��&�6�'|�'	�'k��'Ju<'N�p'2ߜ'P��'�z�'���&a�'9�'V '>ԟ'<1�'Y��'}��'��')��'�''͜'P3�'P�'�Ϋ'�Ó'^e�'@2�&�J�'�O�'�ߚ''�R'x��&g�'�'	'�9�'�4�'�Z�'wv�'�,{'7��'��'*�'���'�O�'�g�'�g>'�a)'=�'���'��J'%Þ'�e�'�N'�؞'�H�'̅�'���'��'�
y'ח'�!�'��w'�?�'Ŵ�'&�'��'Xϒ':�'��4'���'���'{��'�y�'u� 'a��'�$0''�Ȍ'R��'og '#E'Z=�'�U,'&��'��'a�v&��b'���'ʒ'̓'���'��&Qk�'�b�'젒'N�A'��'Q�'���':ߐ'��v'�u7'V��'R͠'���'a��&70�';��'�"�'�'�'��`'�w�'��'�'�'V�'>�'�&���'{�&�d>'^~�'��w'ű�'���'LNe'O�'���'�[�'�&���'�Ñ'`��'�K�'х�'TI9'�'Ŵ�'m�'��'���'�?�'���'\��'��'R�'�qt'�'�l�'k{�'N�t'.��'Y�'DY�'Y*�'��*'���'B6'��'i)�'���'%�'֊'}-'�(�'ZΝ'���']	�'��'�9'B+]'\)�'���&�ߓ'`I�'�S'P�'N_�'���'ɕ�'P؞'V�B'��'W�'p�'��n'c�'�@�'1|�&k	'(K�'�/�'!q�'��'+!�'�0�'h��'�Z�'���'5'��'b�i'���'�̃'�ؐ'c��'
��&���'W�' 8'{Ul'��'D�O'��'���'���'��'�p�'Cs�'��'V{�'��'j5�'�y�'��'��'�z'�A�'���'̠'tΜ'Q|�'!+�&|#'�(�'���&7r�'��'�ڎ'�y�'��5'᪑'���'��i'��'�u�'/��&'�'���'\w�'hp�'���&�q�'�܍'N�'-'�]<'�:�'�1'	�'�%�'Q^b'��C&>�'pQ�&��_'&�'���'.v''��'�a�&᳊'m'�'�ƌ'ߛv'!��'ݚ'
��'�u&��'�'�{?'��_'7X�'�m'�'�t�'w'BD�'�>l'�՗'i	�'
�& �~'y�'!|�'�K'��'��'�c�'���'d1�'[�b'H�q'��'��4��4P9�36�3ԗ4]e4 	4	!4
M4'42W4{�4�w$4T<45�4��44�4��3�84���3u4j��3�14��4�P4ǩ4��4؆4��49�4S4�,4d�3�-4��4�4o�4��344T�4
44��4���3��4���3Wj4�Jg3f�4�,4ru4]�4|4��4>�4C�4�s4�5�3�t4"�4�#4^S4A4w48f4�@4���3�4v�4x�4w�4]:4�47L4� 4� 4��4]�4?�4��4MR 4&44O�4�\4"4Ό3�V4,�4�n 4Z�4\4�64��4��4�(4jA4h�4I�4V�4+�4��4�)4��4cE4>4��4@�4x�4�4��4��4(�4`�4K/4%�4�"4��4�94L�4��4Y4��4c4g%4��4�m 4��4Hj4�w
4��4 �4,K4�!4Y4�`4��4Hd4y{4Y�4:S4ҳ4b4t�4��4T�4`w4��3�4�A4�q4:�4�z4��4K�4�4I4Ќ4��4r4��4��4��4J4�4�4��40H�3s�4׋4AD4��4�B4��4�4K 4 �4v�48M�3&�4��4+�4���3F�4`�4�4��3��4�
�3�O4�4�24g�45D�33�4|�4�b44�42/4��4,�4�t4�4�t4Y$4O� 4Ka4;�4�H4a�4V�4�\4П4�7�34Q��3XB44�4U�4 �4K�3W�4n��3�,4�{4�44 A4S�3]c4��4K4|�4}4N�4,7�3:x4* 4�4;x�3��4q 4��4�.4��4��4.�4�X4�a4t�4>_ 4l��3Z�4��4�N4+R4��4�~4}w4�4>Z�33��3��3��4��4��4��4E�4r�3B_�3� 4���3��4��4ͥ�3xI4'Y4�4k�4�.4�s4qn�3��4�V4 J4�.4�4��4��4�44�� 4�:�3}�4:;4�X4�*4�4��4�O4���3r�4�]�3��4p�4/�4�~4=4a4)Q4��4��3�64,k4M4\�4�]4�4B�4r�44[a4�{4��4C�4�(4-/�3�
44e4�84>4ڃ4��4/�4��4*r4p�44�4�4>{4�-4f54�4��4���3��4nJ4�(4*43�4�^4+4�4�E�2�4+44�4_4�4���3��4��474��4�42$4tB4��4� �3-�4M�4��!4I4��4/�4<�3B��3�4D�4��4�G49�4C4��3(4y4l4QG4��4`�4�	4�4�>4�w�3hE4��4�n4�4@��3���3r4_�4D?4�|4*�3�4 �4���3�G464��4���3Sx45��3^�4ε4+x�3�4�4��4�T4W41��3�4���3��4c�4ַ4�k4%�3Q�4w4w�4F�4);4�4<�4�14'J4�D4=L"4T84e�4�΢3k{4��3乘3�4�(4�4WM4�=4&��3T�4$x4ɺ4*�4]�4��3��4P��3��4���3��4/H4$�3�4k�4��4`4�4W�4H`4
�4nq4��4A�4k��3 4o�45�4��4F�4ĵ4�42R�3m�4+�4��3�4k�4�4�3��4|�4@�4/,4�4��'3Fy')�}'�8m'���&�H�'�M�'�>z'"�C'9n�'��{'ȏ�'3�'�6�&l'	�^'��c',p�'Q-|' 9�&v�'���&��z'=�&���'Ȟ&'��['[j'��R'.Y�'E,C'u9{'T҄'	k]'�'ްz'�2U'�x'�k'��`'�!�'��['��y'՘�&��''��'Ie�'�9Q'e y'�փ'S��'o�^'lm#'?ij'�ɀ'ZV'8y' j')�'	zj'kr'*��&���'��o'��c'��'��&� c'�\�'�m.'�Y'6t'>�{'�2N'�O'�`'#"�'��5'��G'�n'X�i'P��'�t'�Q�&�&��m'��t'JP�'�_�'�P�'�v'r�i'��'wÞ'$j�'��_'�hK' ��'c�i'�S�&�)�&�׆'<��'�ѐ',�4'$+U'}�'w��'A�d'�9P'6�z'�x�'ylL'||d'"i'���'`�'6�'~�&�f�'�:�'�5m'2�z'��x'[$�'�0y'�B`'|��'���'��o'���'�'~�^'�d' ��&S�'�%`'FXu&$�'�uu'���'2)~'���&UaS'��'��'w'�D�'��'+�'N32'qpt'�>Z'��}'���&	�'�x'90�'�h'd�s'8�<'9S�'��4&�-Z'�q'+�b'3�{'�Ij'l�j'�`�'�m'vlh'��v'Uk;'�Mf''��'C#4'�t'{jJ'3�&�rl'�:@'��u'�4r'��{'�i�'{d'j:f'X�t'��j'�v'��'4�r'kt{'��n'{�&�o'���&?~'��`' i�&�)d'��d'I�\'��&�#q'�%y'��*'PYc'�&UV�'S� 'y}'
�'��&k�s'�I�'��a'.�'�a'��o'(\'�Au'0n'껄'Ϗ�'ld�'�b'v�s'���'��'���'�iZ'�i'�w('�֊'�j'x�x'YL�'�'s]'��'7i�'/�0'OL�'�l&<��&ڌ~'*n'�k|'��2'P�'��&'�5W'��'�y�'R'a��&8��&�ŉ',ێ'�ۼ&i�|',�j'�e'�^y'�H�'��&�'��'��'E��'_�}'��{'�J�'	'�Xb'�?|'�%'�7'�>t' '�)h'"��&l�t'�ߘ'�V}'��q'�{u'�l'�w�'E�'��}'VX^',�'��'��L'���'܇'��`'��v'm6R'm'��K'��&�c-'�i'�I^'~8#'�@'���'h�j'H' �Z'*�V'"v'�\e'>nt'��'N�x'�j�'��'�#'�#u'GQz'�I�'��b'�b'gȋ'�Ku'�O�'�vR'�`�&f�|' kf''�J'Oe}'�/�&��='�j�'r-�&��='@Rj'��h'yW�'�"}'�� '�[b'_�i'5=n'/,w'"Z'�4�'s�'�Ls'$('�'hЅ'�@G'�7Y'bB'���'�x'Ĳs'�g�'�x�'d�' �'�wl'�w'/�}'��'�=f'�Ǣ'F�_')v'�'�j'�{5'�qy'�f'��'�m�'%D�&�ޢ&���'{G�'o��'t�O'�^b'��'H|'Eqm'���&��'&M�'�W�&k>t'�&a'Fz'2�
'���&��'ıW'?�n'|_^'�;g'n(w'�P''�ݟ'��'�v'H�q'�3�'/�t'&r{'Ts'��M'�qa'a�u'�6r'_�t'���&���'��`'��'�Xr'
��&�7'޾'P�k'z$i',��'�6�&��o'�mK'��c'Z'��m'�fj'8'Gѓ'�K'��m'|υ'��v'�m'>�r'!d�'S�J'Dn�'|a'hZ�'d�&q}l'��N'ż�'o��'a:~'CEq'.2�& �A'��W'���'�g'��W'Ivp'ʔW'��'O�3'G'"#'`L='�v{'�qP'��^'D�b'bH^' �o'iW�'�T{'-��&��s'��z'��9'�%+'{�6&�B�''�s'�!s'�Yq's߁'��'��'�4i'�Þ'��:'PKA.C�P� P� PK                     1 checkpoint/data/3FB- ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/30FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/data/31FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ0��1XD8�^7�7����!U7%`8��&8��7������7^M7�*��G�0��6��.}8��s8���8�6�0�v�g�3PT
�W=��t�0�k�7<�7�M�v��1�8�_r��ָ��G��@ŷ��$6Ho�7�z�8�&x8f虸l`����ӷ�U�1
��5ܧ7	��<�A�Tc�7g�f8!p/2���7 �8s��h�8�>4��8i�0KA�6�%1PK����   �   PK                      checkpoint/data/32FB ZZZZZZZZZZZZZZZZZZZZZZZZR�4�v�5ن4���4�f,5)N�3`�4�/�3d�@4�`5B�X4�!�3�,~4!Uy'�J�3���4:Br4��-5B?�'j��3�wb/b�4�TG4�D'Ε�3���46�4��^)mO�3���5���4�95r�I4I�44�4�<5�S4kk;4<��4�w�4q��-��3��4��w4z��4�{G5YM4��*k��4aqF53A58�A4v��2N�I4�,(��4��'PK�y��   �   PK                      checkpoint/data/33FB ZZZZZZZZZZZZZZZZZZZZZZZZbG>��5?�2n?�̫�`�<9 ��h��W����;����>�C3��
�[�k>?>2ǒ?RA?(�>E�@�>F�/��ee� 1�����!��>Ξ��ND���Լ­����#?a=C�R���p�?Fp?�[����=?�ލ=x>?�����~��Ws�3�Q��)�?��R>�:�>�ˆ?"]H��/�d�Y?��0�ѥ>	Z�u3�F2�=� �?t��?�H.@�P;�8�~>
�L�@��<�+�?_:L<�?���?��3�1䂿!⎿6˽�b?��4��E��e;|>�.�?�>�%W>1IY���ƿl�>�7��Sƽ�v�7G��ɿo�h����=k�M�"��?��@�D�?Ct?��=��?ɴ�?mj2?U`?�;R���/�ÜU?c�=W���-@�ԾvC����?G����g?O>?���>�X=��y�K?q��?i��?|n�<��.����?c`��x���˥��@h?2�]����	�L�9aۿW�?)�E��g+����]ӡ�Xc�?eX��PN}�E�`?��������{=7�����ҋ3�� @�ڱ�������c?�
�?Wc?5f�"�8��Dx?è?q�?�J޿m��>+�?&�?4xS"�N�K���w���վRx�f:�?^[1?|A���4p>�w@B���SLa?z�A�L�?�9{��A�/���*@��R?���?�7i?ՌE>R�,@>�:��蝿�˟?�+?���>��s<���=>�Y�?F�>|�y��;�œ_>< ��qM�>$1�atɾ͎�:⿏׽Rdk��������m��^c	@��?UmG�R�?�y��H4?(��>��?F����>�r&?O�{�'�?��F����� ?���?:5$?��=��L�E��}>��?�LJ�H?��=p9>~��?����r��j�ľ�pQ�}�>����?e�a�%)����I�4���t������?���?|�??3�s���41�?ԕu�v��?�a��!����w?��r?{���4�?n���,����;��rI��?���Ӊr��j@̱�x���̔���@T^�?�m�>=4�;6�����c?^��?�a)����?���>C�?lr.@��@��ν��?1a�A���ʗ���?G��t���֟���I�?�J?�x� ��.���V?���??/�>��ֿd��U}� L1�Z��L�G?�
@{�"?H�#?�\�W	f?.MH>�H�1��x��?��?�>	�>?����w?� �k�,=��?��s?r#y�ß��-n���#����a-��X�?3.��>��;?��2>��w��?����g]��=ca���*?�e�pVK������:�?��#?�Q,?#����wg?�D?���>��.?u�>=�>��U?M�o?C�x�
N��6콍?h�*�٪�)���������=�!۾�d1@]�D�>	;X?G��?E�>�����
���'t$?/u��&�S�y?��&>��r�5�>r�[��a9@ )2@f��?'Ĕ�3@�5�>�H��O�W@kA�>�%�����7:�~�*��鑿B�#���>����?צ?��=�2�NX��!�]�%r>�,@?�_L=Ap�>�4 @�Z��9D����?�;�?(궿�n_>�{�<���������?����\1�&�5��=�?��*�����C�}%O���=�R?w�y���>��(>M��)b�y	�����(^ؾ�m)�}F�?9��>�)?�����>K(?b�Y3�G��>;dx>�?�r�A|���l�?�|�?"|����?J���Ί>��*���/�n
l?�܂?��.����>�v��uG���C� e���3��,��?x+��*�̿x�5=b���] c?4�?�>kG9��%>�AV��+F��ƾI���!D�>�8-�=&�?w�6>�N�CH��9��Ƽ?�uӽ���?�6���F�QR�����>�u�ٻѿ(1��d���o�@��t��?Μ�#Pؾ+]�>L��?��)�{����?H���k�d?>L��\�?:f==� @ S?E�t��K�dz@I��?+�$�����A�?�$�>�C���;?2#�>�l�>�J�?���=8�?N�g�a�/?2�a���p# ��>�?��	?jA@=�)��E@pn��{�'��6۾��ӿ�Y?f�X?& 	��UA����>�+ʾ|2��ML¿��?����Ղ?�3�>������=�ͯ��l���$�?�Eʾ�zl�55@�oq���� �O��?��S?�[@/�?7��������P�v�Q�U?��@����|?��6@
 �.��A<?�F�
�N�Q���Vl����?m��>�a~�~�s?��k?���?����I?R�N��WE>Dծ?=Կ��'>�����c,��¹?�þ�6�P�xO��]�.>�z�PX�?Vk?''�!JN@�N?||���`?T��=��Ӿ���m�G?`-�?� x�6��z��d��?R��?Q	L?
A�?J^Ϳ�,�����?����A�s�����
B��\@u�
?k2��n���.?c�*?!�@�:? *�>���~ǿ��?J]���M���^(�� Y?�O�?�S�>b��-����>�ܫ��ޥ�7%�j(�Io����?�6��a����>��F?�;##?�V��	M�#����0?�P?'�C>"��Q��u6�>ӝ�I�M>G@&?�j�=��;?�R��L�6��a�?��>XM>{?B�۾$P>sҾ��J6�h?T���_�>��>�*�?�
�>��=´O�4�?��G����?Y�3��m?�Xe@��>�½�V'@�y��2�O�v�3�+=��N$J����?�mX���V��&"��9���(�?jw3�-��?��@
Ӧ�COϿǱ>��?[�<�R�?*��?#��>�����}�HD��-��"��c":���0?YJ�����c��>�=��[�<(jt�W�4>��Mr�8�s�3�}?­Y?����"��e@�^r�a�_��͢��m/�$�X=������"?�zݿE�=��?�?;���-�?�A������0~?�=�Q�ML
�j�7�N����c�0�?�p�>�	�?G�?�K��<���>�:��0����?��?��T?�����	1�?�ü?G�`�5��wL?F��>Vb�<�ھcd�Z��z=��Ͻ��?K�?{��>CNW>#*	��6�?e�'���?�B�m�>x�[?�g�?���>*�9����o�l�s����?9�.>���> �?ʢ_?j�>p>׾��?�y�?bO�>���?6�>�q�\'��!־�CL���4@��1?�)�>�g�?�L��#�f�0F�?H����]�E2����?s?��0?Cq��3ݡ����?�
��n?�?��?�����q>��Y朾aq�?p��>J�7?!��>8;ɾ�Տ��X������}Ǿ�*;?E,,?�(-?�/�?�RG??�[?t�4@SM*�aG���l��\G	�HB
�Ɋ:>�;"�f�?��=9�>���M�?�a�>mh�>�
(?!M�?�d>�[q>��d?>����R�?B�����>�?��>��-?�n�?VP6?X��W>"?�C���0?��#�a:?&:?���=j���e�������t��4�����>��
���C�?|�>�y?�L ��#�a��x�
�~�j�{��%?���?��N?�Az?�P�> �R>��?��!@\T�>���>-l�?Ф"�� ����=py�����>���m�F?�J?v&�?G2�=8���/>y�>�[�>���>̧�?���ԑ�q�=��?{�@��J����>:�����>"��� �>_z����>�N�?v�?�+��R���w'?��>�a�T�0��4��?p�uߙ�P�	�8��?��?>̕��g���	�?�?��T�3ҿ,F�>��?'{R�
�?��>��b�u��?�ח��|�?0�(?e{C@���zG�7�u>�%�>�?T?�=@g&;�"�����<�[�?"�׿�h�����?���>W�O��h���
�?A�u?�羽����#��e?�\ȿP@=�U�<���?#�)���>�>��?7)�?X�ĿY��?=���N�>)�q�ټ�?9d�������?��?��?�hо'�>=Ң>��¿��?<��>ٶ����=��,?uX=���?e8�?>q�?3�i���y�J�a�!=&t�=`����?=�@�zg�>��>N:����<��	�p�?d�2 w�����]�����?v2���>B��=)x�?��>&$�>J~���Ya���V?8�?��?�u�?h��=����9����?F":��U�D�4>}���1���_gJ>��?
����>�B�=p�;��i�Űx���)�*H�� �>�TN��4�:�\ٿSi�>���>�� ���=���>�� @�p�9�=��?�җ?�P?q�4?��X����>�?�B��~���$��la=&�>�Y4>h @�e8���+�E\��[$�>������?���߾�"�?�>�Q��7%5@2?�ܪ�u��?[?��m=���?&i�?��>�q�>��~>u�S?97Ծ/|�?4y?-�1�>��?i�^=�q�>8e��kJ��a��6��? ��>"?����Ϙ?�#?�1��q>���'���ت@��?]A羿-�?�?_?�:�X���]hƾ���Ŀ^3@@��?��P�'����$?w{S?A#��n>�?杖�ʵQ�F?l��U?�5��~��`Ꝿ���=>!�>�<��`�?ㅟ�f�+���?{���M���v?�M���^?Dp�= �0D��߷>諒����N�#?6��>��>�_���?�Oa���?�?���>R���;��c? 2?�A�?����::�>q��=��	��?�9���־�V�?5N?J�?Գ�?a�6����?���R��gĥ�S�v>��?��Ծ6�?���� ��u��?bV?:�i�]�?���>��j��У?G�?o?�o�>D?&����7�>Ƈ���ko�ӈ7;�|�Ҕ@?����[@"{#�M�?���>����оߩz?G�տ"q�>�?M�m��>�o�?c]>��>sA����>\�Q�	�?��ľ6zǽ ��?G� @�I���)?|fn�dR�X�D?�r�>�ʾ��<?�@��X�?|b?��@2p�>q�?=�ؾ��*?�}W����?�܄?�t�>�?Iڿ����>�i���п2 }�5�>no@�-����1�?.�~�؃->�B�?��׼��H?�O�� =6O?/^���@vӿV�?|y���+���۾�פ?������>fX�=�E_�y��?E�<@���=~a:��l�=��q>FB˿4�>��ƾ,���+P�?1���y?�����H0���ɾ$o�>6�X@���?�J`�ɧ˽��ſOP�?v���Y�B����?`LH?�?>s?�%�>���q��?<�'?�0<?5{�?52$?����b,?ݒ@C�-��L�? _�J!�����]�>W�{?ė�?ul&�r�>��a��{S�O�?>,*��Ʊ���>0u?[~�����^��� �>�@?k�{�6E��Ꜿ�&�;�M�?���>
�5?d�οSX?θ�>PK��ED  D  PK                     < checkpoint/data/34FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ/�$>�I�=��o=�M(>�,�����;9�<���=���d��=�R�>5G�ҩ־]D�wU��4>1@>�,�>�2�>%W���(�����>�RO�T�=Gݜ>!ԙ>e`���>.�)��|���xK�����bp�=�̄>�0�>w�>k�w�����"��+���g">r<�<��w�Ma�= U�=ϐ�>ݤ?=	D����>��>`�>#o�=�UR>x��>��}��=,Q���=�̼�F�I#�� �@��9v=�ɾ{�">,pȾ�n�>�9�>4~
>8��>g>�>�L>S���Y샽s�=(�>Ѭ�9@�>O��aHȽ�O>=d�>¹���B�t=l>ݭ�>�ԗ>��X=h�H=�h���QE���
~;���>?�>E���N�M>�.��Ի&Ub���'>j�<[���R(�=��>�M��T�J>vX��6D*��g>���>ٲd�oB?�cI�ӊ�;��K>��G���e%>	O>�=��]=��Ӿ�y=�_�=M$>�+9)Nx>�qϽ�@޽�?.��
��u�>���>����=7ġ=�nL>�;>Α?���QeL>Mu���=�z>��<����(k>e���\���1E>���=�Hw�SG�>�%�/�b=����$O>D�p��K�P8>�涾/{ݽ��7��n>�{1���>`��쉝�7��>򛮾p�J�v>Zr�������9>�<־�"�/3���
�z`þ�X��M��=id��T�<��'�>�^4�L>�!�`l�m飾��=PiZ>�|�L߰>UM��i2�ke��cὌ��>E��=z��;m�;�h�Z�*>�>���>"��;M��<nEd���a��0�<#�>ߨ`>��=�>.kϾ��R�ё�:�=|�8������､/$��t��^�;nN��pe<�4>�@;�a_>�)>Z3����~>E8�;ql�>�`X=j"�=G�����.�B� �@��F��>*f�='p�CŽ~�پå��#ٽ+�<��>�S��Z��<S�<>� ��lAb�9�$�4s��;u��v?�>$�?>5-�>-=ؙ1>oT��)1>�$A����<�%��ٜ�>ᴙ;u�_�<�y=L��>����b@��Ž>o�+���L>������>@s`=QxF>��3>Fk�(2�ɧ�=����	u��:>^[�<�Q=�ڽ=ѥȽpv������H�>̷�����>��5|�9��#�_��=I��=L�/�9
[>�==�{b�H&>Q�>�&���>��>��S>�;C=`������o���M>����Krb���4>��>�1?�J6Y�\1>sԆ<�`>�}k�M2�=h��=��p�����>.��=�V���߶��ޫ�f��Z�G�?����ڗ����v"X>�z뽍�m��齀T=�fh�����Ԡ�������$��XN�xl�>qYȽ�H��g��=�I=b|��^�*���c_c�H�<�5=;�ż���>�'�m���s=�==۞<W��>��J>N�>Ԍ���+C��Y�>`>NA�=4�Խ����z^�+�p>��H>��)���r>�>�>���?p�>l�O>�,��%E��ߨ>
ݽ���v=HBC�+�������=��	���?��۽x�>w�<B7�=� �>l�>�$�<�p�UE�<�f<2�7>\K��L~��7�� �>�K>��J���D����=Pv}>~E�z��=qB=r�b�A���>%=�>�n�>ln���s:���3=4�>Tҭ�A<H�굽�������J��7�F�G���|>�~�=�U=�R(>�Q�<���<���Qq>l{#>
ӥ�v�>ZfL��8�����/��x�;d��>���q�=e	��c=٫Q��>��1>l����0�y]3>ߩ_�{1.�E��=i�:�Z��^�<�9�=0��{1��m=�?2>�%�n����=r2������ ���RĽ��;:��>9�?>Ҽ���T�=NY���<1>�ξՌн0�F�-�h=�>�M�>>�=!�!>f��==����=��{��/�<��Ͼ�<p�m=����,Ϛ<%��>��u��a�=�"޾�:��Uy��Z~�D���牾B�����=x�&�o�"���$Q>�S���UB����=��>�8U�(~>�@>�򉾡}�;$@e���3���>Φ�>��ֽ������>���>�=YD=T�>�r�>���=� �>N�=4μ�ߪ>��+>�E��=S>�l�>*��>�椽G�S�}���ҏ�\2��>�ϋ����=���<NW/�R@3�ӱʽX�F�C�>��G>���������c5���1>�rԼ� ��p��V�=�uF�T�k�`�:��5ɽ ���7��>�y�>�rF���=
|�>�{A>��ȾU���r;-�
����PW����Q�P:�<��&>���>έ���rX�̉����>��=���>�1��)x>ϕ�>���-Ǽ=��~�)s.��{}=<\�U>��������CF>��c�F��>����H0>������;(�=�Y`>}�N>|��=��-�=��>𭻫PD�p�:��q��
n=L>�>�=9W���z?>^�:*�<�})>z�<������=mM�Z�/�>g�=��&�%ؔ�n�=hN�C��>h��>ܬl>N�u��9;>_�p<�B����>X@L>}eW��BQ>�2���#=f2>*�q>��f�ͤ�=\�F�����ր>'�#=��#���?�DC��	>W��f�@>GE�>�җ>��<4�=�@ݾ��;��j���[=r�>�"��
\�=3�>�%i�yU��EU>�w���i�ܽB��N1�~Z1>\7����>Y����>�k>"d�=r�J>�v�>pԾb��=��>���<�D���ɸ>G��;��=�Q���>7� ��̊��ھ�.�����|�f=��>oK��<B���TL>��]>⃾��>�8	>�@�ûw>�[w���)=��=��.<�H���邾=�3>���=��>-�5���>��s>����϶�>2��=��>Q'�=��[>�q�>�K>w��=�޼=9Y��o�>�a�>E[a>8W�>!�~=@�i�.�>�QT�i�C�.z�>al�>���=���?qR=9_
>���=���=�>��>J�,���=u���塦=�ۧ=q�@�[P �յ5>؉��Nڰ>Vʻ�aw4���z>���f�=z\�>�x�>(��݌H��<�<`�	�{7X>V��-�<�w<>�R@�j����_���<�{d�jF�>�ҏ�%�ۼPmv�.�;>Y�1����>�D�>�>p�Z>D�V�V�����>ij;ݧ>���	vX>v<��a7$�凥>�M�>Sme=�2I�G*�=r7[�h���f�=ޛͽ�� ���2=��<���=<Hr>��)���E�b:>%.�� .\�0>���]�>@;�>���읾Y��<��&>pq��z�F�>[�����>�;4<m!�=�5$>V蘽G����>�ĽD�[þ�^Q>8��=9]a=�F�9sr>2i7��;.=���B�>�=3�$��Q�>S>L=��">�m�����>Q��4�=�J־O��=�ǚ>Qo�>0�<���>T`ھX ��tn2>��4�e�=YL��5t۽Mc��4�=�I��Z�!�,91>�n�>�=$>s�\��y�=���>��=�M(�x�G��D>SR�=�/�P�=6f<�CG�ʅ8�n������=��w>J�o�[~Z�pLZ�y�>��=�Ls>���]D��*�>ju@�������>�V��=�*�>�n��[�����>�R*�� >���7��=�V>�Ἵ��½�Z��5���j�B>o>�*ý�aQ>�\�=� =�H���Ѽv9:�LR�o�T=�½��u�D��=<9��M>�bR�7:�=Ht�=�製���=`!�=Yx>]�����,��T><>�
J=R2 �U =�hw�e�������q�=�m><9U�A3���s���*���=�V�>���,;>��W���8�'��%�->����'ߡ=Dc=�'�>� ?��>̢'=g������R���Ҿj��>��=sۆ=���]��m�=>;�>~����V��QT��e4����>�D�>ES�"n"��9�>�7�}����v��I-�΁=[��=�[�>���=%dM>^G>�tk����>�O�>����P�j>�}��9�+>H�o>`g>Un>�ض>)�~���e=�轄2F>��>��>�И>�=,8P�4�e>��{=��:=��,��ɼɬ�>��g>�$�=ʼ=#��=���>T�P����t�����T>T�=-����uҽ~����^>R"?1hO=�8>�e>�a��@�E=l_�	�>���?���ɽ�����JϽ�w5��\�<�>1���
=2��>~uԼ��y=�#>v��������i>�K�>ss>�!���~ǽ���>ۢ�;�!�>�����{��<��>��>�p�Jn�_���Fd�=4�5�w �<�=_>��>]�t<I�N>6�a=f<�dy�>�/���>	Rڻ�o�$�;>ƚ�>ۻ>� <Y|�����gl>)��>��.�h�����s�x�3���>��>ֱo����B���b�=e6M>���>	�>`��=���>1�>����Ͼ���>������T� �a>E���/�G	�>, ˽�S�=2�=��s>p�t��<�u"�UҨ>?=�� >�;��o��:�s>�V޾t�5>�T��X��	0�=F�>���>�_�<�F�K��x}i:��=Gg8���x�E�F�M��Y8>��=yv���_>sg�=<?��_����cĪ��U�>���>�蕾
z�<5i���4>��轳qO���8E^��ؽ˴�蛐>�堽YO�>Œ�3����>Ǟ�=�ۖ� ��a��k�X,E=�����>h�T>s�=3M�=��>��%>�|R�n����Ѕ�$�>�>1 ��>K��=6H�߯d��ݭ=������=��>�>l�=�B�r-X=ދ>����\>w�����OMϻ"ro����=R~S>�ո=�9#<�)#>6d���y>Px�<U� �����P�i�[9w>l�O� ����W����=U=i> ڥ=Cl��Dd�v�=�ۡ�E=��i�y�<�b>��O��0>���xy�>��<��X��k	�����Â���5I=��=��1���	�i�:X/>�a����>XҚ�B�Ƚ4>�����?j���_�7>,#�T�ϼ1U7���<�1?>���>��j�j[�
�>J�K�/�q����=Wϡ�F	ٽ�U�=��=�%>�_i�)�;�ｘ��:��0�\> Z�ߐY��O�>�$��+$=�6>4�f�-O�>`�=�G�HG���;�=�О=;K����r�޽!w7>�g��"=��l�-�-<��=�#7��5�=�_�l䳽<# <	*>r�I�`�>[�>>�.e<�i�=S�>&K��G<~K�<�Ⱥ�o����켽V����S<�n��HZ>�>Y�t�b�!�"�ҽq�w<��1�����E���Y�@��>���=B3��Ȥ=⫵=���7��������<�=S�.ҳ����=�+�tVb� 	��c}�\;�T�>�[�>bҰ=�-�=i�>��>�'սj��=����3c����g>�?ٽ�.j>5�d=6�<Pk��k���>��Z=�5�͐i�ռ��>R�%�8D�>~��^G�=��=�y�����>��I�U�;�K� �4^z���.�慘����<%�/��m�=F�p�n�Ƚ��<�:�=(��=�R޽�o)>yms��2��ڒ�Q�=���< E:��>ݳ�>.|�-�P=�]D��1�>�����=�<��I�HN&���v�,���{��=�C�r� >]��<H>��m�A�A�s�&��R�=r9��>B>�Gw�-,-���U�6`�=9�j�d#>�yl<3yz>�����V����>� �;���=����f0�6.>�f����=[Ȃ�'KQ�鑤������9;>rmo�� ��b>�/�>e�>n̟=
])�O�齚h�:l���r:�>�O"��t���>q2��T�=��=���=�M>� <�醾A#�<Ԙ��� N<!��=��t��y��d��4���1ӽ�u�>2��� �=�I=�a%�z� �f�=�l=:���"�>�xz>�Q��A\������[�=Q�e�6l`��#i��1�7׭>�z�=k+��������>�9c��}y>��}��=���>���=�ږ=��`��+�>����\>��ݽ���>k����5�y��#.�;�1ڻ�s�>���<���=��=��[�RUB���>�:�C�E>���;�'�=�HQ�W�=���=":Q>�20��a�����1R��X�;|��?2K>ԣ
>.�3t1<P@>�F�*Ћ=Wg���q=N; ��i
=[��>$&&>)5�=]�>;g�=��=>��'M����S>��E>3�H�{�A>���=��o>�(��+��6m�=į8�VJ=��h>�Å�o�����K>zL�U_H�
��<��Q�HS�Vm>��q>@a���<t3Ľ��;N#C����j~Y�VG>'�>yp��6����<��>����y����
>��T>�Ľ�m�=�ʼ�n�8��rN��{���?�������<�(>�/�<TF=�4\> �=�.�|�=�m>6q�dͽ��S���#m��C�m@0�@\<���=M��=SĚ�&�=���R�k���_>-؜=n����>�>/�v<ʆ���t>��~�ҫ��"�I�֣=�����=��+>0���8>뤆��K�;���^����<�y >+��M\�=�����c=�����l��ؠ���y#�m��v@��^L/��Ƒ�붷�8���4׻X�r�tM�>#!:u`�s�3�L�b=Lu;�6��=RB=JA>�Q>=n>��߽�9u=��F��>.3�>)����<߭Y>vD>dڊ<���`���V�I<7�"��eܽ�\=Ma+>�<�=��^�]EF��5>:l�=T��=����is�a�̽]'�=P�c<n3�=�J>X�:�������y�3��x>^�ռ�>�H۽1Ť�: 0�q���&Z��j �ژ�=�Lf>pX�=���=���>�ZW������a�	Z���+��C)���)<��=@Ib�v�Z=���=�z�>ة!>w=ò�x >�.��%��>���x!�S�J�����=p���ݗ���e>t�I�@�e�0J��o#"��r
>� �=���=��@�+�����=z����
W>x��'����K��ό>
W='`n�P��=�n��FB>�<>��O=�5н�W�=r*�� M�D���ׯ��\a@>�+[>ƍ�=p�=�Ww���;��	���>��3>_PX��A>"FF��UQ���ٽ����[=�膾w��=�hL>۽@�d<�s,>PKV���L  L  PK                     4 checkpoint/data/35FB0 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�*����ö�=/=[�Z�^���QL���=�"=��ż���=M� >,K =YOG��!E��<l�ʻ�M�2�<�>�Zw>������&;�ʆ;������w'̹����qM:b��SLE�
�:����v񀹋)�� =������9@:�|���o���l����͹��������"99��,�����`:il��i�<p<w�	:�=�}�=��K����<5�;���<o�<�L�5f�Q~�� �<T�;�\�=Fv�h?/>-_нА=(*���^�M���#=n��s=PK�,  ,  PK                      checkpoint/data/36FB ZZZZZZZZZZZZZZZZ3�>lF����=>�)��a��W3>d�=��.���<r�=_}����)┽,�=�/5>�F�=-NF>}��Z��=��<'�&>zL=PBM��	�;h����(��x�=�|S>F�׼ł8=��W<��K=�dm=�=��V>�5|=p�>�ݽ��4>��=�U�<*�u=$�� >k��������.��;!�_�p߽ʟ0���=����Rb�v��=�V׼�%ƽ9��r콝�>�����''>����՘*=f��=?�?�n<��0�q�0��t�=t+>�!,>��+>ߣ��_��>Y p���;@��b$7>�)�<s}�K���
�	5����=��/\�!�W>�b�5��=���;�%>����1@=��`=��">B���a#�=㢇=�~>�X������=��<��ƽIG)�[g:�x��5>CC]�x����ػ"0>>(�n����w�>�( =~������R��=���=�J��Zr>�;���R���M����	ϐ=Q\�=��=��=6�V�n/ǽ���=��>vt�=.�=�mΫ= �G����=�x�=��=�!>k?>L�7��Q�;��/�� ���B!�~���k=ν����>T��=:o">�=��)��y-�ƞ�=�s
>&�����Q>����C>�W�C�>�N>�[>���=?�=$��o;>�맽���Ĭ.="]1���=m��>]�L>�Q=�"
>�u�$��=�ְ=�W�<BO=Rt>*�O+�<�0���=��+�	�S��T$={.���h>v<�>��Ľ�>������=d E��k[�y%��>��񙽹��=��݈�<�櫽W�=��<�#>'��Q�s>U0���ڢ��G<��E=��5>��>#1��L�C=2p�=��v>��	�� =���:�H��妦�]�N>V�j>\猼ZdW>���-��.�%QY<
�6��Sb��-q����=��<�'��>�ǽ{n5��S:� w�%��r2��TU��m<��4=��\�
w	>���=X��=ek�=��=~�?�
�A>�6>�/�=����=�k��]����w��/Ⱦ��7i>���l���ؽ#3�`��=5Z�;���a�>#���0��+>¨�=��^���<;��v�<�E;� >�~F>�	q�;v;���{�daC=%��=��B=�����u����<q�>3� ��3�=�i<=ca�3<�s��i�
>�ѽ�V��#���'��2�=X�#=y��=Grm<Q~�=��7���>�ߏ=Kz*>�`��v��>:0�=`���3�>���TY>"��=�M���N���=Y��=�O۽ٍ�
�ͽPyR>ⲙ=d�/�v
<�o�X��=����i�-�N=ԙ7��J�;D���a#5�E�=]E������R�X�O��=ϭ˽�=���pg��D֥=�ɻ�>�=(�<k�E=�{��41��C �w$@�[HG>�Cw>��<�d,>&��E>�������a����=���<�ѕ=�J�z�=�k��:*�'�m��16>�T=����H�L���>Xm���*>�5>���Q >u���甽A�����Vg(�z��=D����н=F��uϔ=�ܖ<%���(-�����t��<��)=���=��L�`�ռ���=�L�=���=h�
��5߽��7��>N��0�j�͢=��L�Ǽ�,>\�K>^͓>��g��$�=_[��^r����=��>T�>�!�����M���ƞ=2=9�>�r�=^�A�-�->A�E�6GC�9�#���\��h>�J>�oD>,s=v)A=�o>�i�=*8�>	ND>��D=��=V (�l��=���d6�xX#��������|��;�;���=1��="��=F�=񮓽 �;�g�>n�c=���<bP�>!�P�G����<��F=�Ｗ��<�J<-�t>�=���:9���=�#�b��=4�7>H5 >�s(>چ�<3���u<Sc�=�!�<"󞺭@>	����l���~��Q	>=��=+n ���L>>Ʋ�=4ѽ1(���
��&�<�!G�r`>�:��-�=��9>)��>~9���:�(�$�\+5�T��=��U���=��=P1нkK�-�ν\��Â>��>'��=�s�Y����Ǽ@� �<9>���=��>ڭ���	=$�>��~<�ऽ�JQ>x��=��M>	�8�`��=��½N�=iU�<��b>y�A�	>���3R>�-�E���g��<�L�=�">'9���1�<=� h�E#�3Kq��&�=��>9讽������V�;i1�<>��~>�����!���A��,�D�=���S��(<域�~�L>�����i��<��=!g>�3�����ݜc��2������*�eC#<���=^�=Jo.=o~�<Y�t����=+�G=<���X8�/�>z�V=0�E=�������e��)B�;���Z{���>��qy >�iV�PKY9N�	  �	  PK                     < checkpoint/data/37FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�*���Ƚm �=���< Ծ=L�=jV��E�D�`��=���=P/������UŻ��<�����!��U�����\�������^<^ч=�v�Yi�����PK$�Umd   d   PK                      checkpoint/data/38FB ZZZZZZZZZZZZZZZZZZZZZZZZ�?�=i��<'�<`��=7K���-��$w��{�=�G]=�0�=�>=�g��m�=�Z�;��������Eq�;T�]�������7����=Dz�riԼ�:=�W�<�@ۼ7a�<�A:��z�Y��j�;�t�=	r|=a%
�+ȼJb=��v={l�=p����D=	;Ƅ	=��V=^�C<(��<v��� л��=<緽��4ݼ;����"��=���cܡ=  @<X�wU����<��=ő<=��5�F�μ0wO=q�}<6�<��=k×=�b��=<J~1���\<�Y�<S"\;n�"�F���%G=߅<U?�=.�9��I%>���X���6�:�i�/><�D�C��=�r�L=�=m�$���H=f��=����!�=Y:=:R���l�<����H=h1G�+��=a�>2KE=*�ȽOQ�=��=@a<xB̽�#��cwN<Ղ�<`߽���=��<Hf;��=x�=E�%�������#���=���==s�ѼN䌽{��<�u{<�nY=<��<�����Ž�wλ�U�=d�M=U��<��׽��<}0�=f�佰i��)o�<{c�:���=#F�<�\�=�9~�����Nd�����=.�=&�=+�=�-�<�н�f���n�;RR���<�=�\0�̨+=����S��(>o7��9>"�i<�B<�" �N��<��>�Y���G��ц�E6����=��<&�3=�׌�U=i�����=�(=ϟ�=���=9�|�O�8�!q=���W���JvW>G�=��R�_��>�f׽�߽w���+�;=�L=zG�;��R=�����{��AS>�-w=ʹٽ2�0�� ��/�7|)�H>��DŽ�l=_�G�+Ͻ���Ӑ.�� G��#�=p�D<�ժ:~����܈= �߽��;)[-�g�^��b�"D�=$�[�抄>�{��ˡ�gm�f��<�>�H�,���R�����l�<Aʋ>�F�=��<E�==R��=y�R=����L��=��Z�1Ӗ��>��G=i�<(y=�1b�<�D�=��=޻H;�x�=𯳽̐νpm�=��<(��9IR��=�7�=(�ԖĻYC�S������</�@=������*������y�<��>�Hؽ.J�<�Օ<)�=ތ�=&f���<�c�<TI�;���=x{f={�a��p���*<���<�-<����=>�3�0�S==���K�1>p�u=���2���OQ�=�<I�
>'�<�˽�I<F�=��O�#>�#��e=�*���j=�歽1�gOs=�D=S?�=�-=" �<j>!:%����� J>+�'��;X7��+��c�O*->�f���=�d���)<C�J��խ���<�q�����8s��ڼ�=_�=��¼�瞽ģ��=��S���=���=A_�<�Y<�/e=��J��<�TK�=_�~� R�:)>W��=�����f�=_����Q=�Y�=�����v=���<O�;��=��=؉޺�.�o�^>M�_�1�=5I�	߼D#<����<ܑ��<%2G���������>=s�L=w㼝}
<-�<���i��<sA	��Ml<���=��<aG��k��8��׼��
=�e"<G��=��<=�i=�<Ô��9ҽ¶���Տ��r<Om�=�n<�$��|ø��<��2�=�A=ր�=}V���{�=��@<�F#�So�<� �{;>���=R�#���=M�;\�*���u=�--�u��=0���Y�`��Ύ>�������<���?T�=
�O���t��+���e��Wo�Z�3<z�=���=�{�:���:bԟ=�g���od=�	�1��=hgJ>���l�b�eZ����=M�𽝙�>�Y3��"�=�<��x�B�I=�s�� >�b�=�m<���g5Ƚ*����Y<�D���:Լ�1>���=�@!�	8�����|V��:�P��<�:=9��=��f=����֨�>j���":�=YQ�]+�=�R=\"�Ai-��=t�6����E�:=	�=a/;W���A=��;[K���7߻maR=Cm/=C��=P(�=�7f=��ǽ!쑺���<��w�={�������>�t��=ٰ=c��=�J�< � =�mj��}<<"�v��1ü�?<j4����A�ϐ�<��f���&=������<t�=��=k���#�R >H�Z=*a=K�_<<*�z�ߟ�Hꣽ�7����������<��<����'a;��P<�ԓ=d�����=>\=����z�=B�F=`�;�ϩ<;�6�n$�<�̴<4�,೽|/�l�s,�=�5�=̱=��=�%����=��d�Bd�=<�=\�=D��=���=���eּ�Nؼ4lX�[ժ=���<�q�=�Y�E�6=�����0��z�����h�e-=�;���6�=�d�=��ѽ�0>�V?�;N58��,�= Qx�]�_���>�!�=4/{��z��3/|���=�P�=t�=�)�<F���=~�U��ŷ�?	=����"�U�=:��=/f=N${='��D��gAf=�!����<26v=_Ez�3�3�-Ƽ�w ��l=T����g8>��;�O���o���<+��<G�=�]�<�*����`=(ZC=F��=�����=����~ݽ��#��ʱ=Y~�:����}�=]�<�a�jPü�.��[0I����=`=�#\<DM[��:��~�<��)�����ʟ��� �<�:������A\=�}�=-s�=��=���"��=�<4L�=�F<i�ý���<�>� ��5��[q=���=+�>�0�=��½0�Ľê�����*?��Y�=�p�=[(D=6m��J�#<:��9�=���< 5��bX�����=$��<鳕�lp�>�F�=���=���<d	z<vx&���/>!����Aټ���<�C�=W�O�,����
>��ƼŎ���s���#��n9>/b2�br�k=<C0�b�>;�f�44�������<�\e=��<��=f�&�����5	�@��<��[��-4=v��h���}1��ӽn�ǻat}����=)[��XM�=��=<���X�=5d=l+���1Y�Ǎ�=̠��H�V|�=���>�=�5.��
���Ұ��?�<DJ�o�>o�}��R�;hn�~�F>�?�=�=��^�9�����<73;c2�=<�н��=jVM�N��=��f�ի=�'�=M�=zj�=\�N<��Q=����/�I{ǽUK=�֙=lOi�|�����_��� ;À��4���%��'��=�&�=Hr+�0��̵�<,>��<J+�= "<��Y�ȹ��X�B������+��(���z#�S��=y�>��ｾ��;N��=�:=)��@q��~F<t���V<�h�����)�K��Ź=��.=(��=b
r��z-�?�.>�@�=S��=ݶ��`���p6(=��u�Z��٭c<}�=�P�<*j鼐���=*>^��=m
>���)s\=-8�Oa�=Ui�;�C���%=[�_��۽c5�����<��7��k�=o(߽��?�8��<���=~���� �!��^�0=2�<`���3�r�N��Q�<4��=��Z���P�
|=w1���.:=��H�(]#��թ��ϗ=�=�=h0������=>�.�=��9���<�J�=�<��=�Ќ<N܈<(��主��=0��=�/߽��=�q޼��q=dҞ=��a��۾��vʽ~r�.�>&�����)>���<�X=ɩ�<^���X=���xŽ8lW=G[<��r�~��;�y=3꺽n��Kf;�b�L>�M�=�Q����<L�2���=�M0>[��<*��<�^�=^�l=�}j�lFŽU/�<Q�K�#=�T}>��7�}����u�=*g>�z�=�+<��;�R=PЌ=���Z.�v�V��>y1���2���)6>�tr=�F��8��=�x�=��J���}�n��2\O>��^���	�:t�RX�H��z�=,f8��g�9�wB=Aս�@��(�<I�/��V��*n=}��<��:��i 9�'���5 �̏<��.�.��<�k=uS�;�%w���<9��<B-{�|�v= �f=�
���[�����.{�<�m�<��E=������U&��(,�;��x�b����x���ؽlĖ=�����S�=��|=�
!��=��{�<=P8p=>���󓽙�Ի̻ۨJ$�!�<D��<Z�=j�<~$>��P����:m�ռ���4r�=�;E<|���%Y&�Sd��m��n��=�)���h@����=(��=����Q�=�����6=mb�=+�ݽE��=��=�O�NIf� !��k>��M�<�'�=I!�<�S�;U>9{��楽/��<֜�˹�5���$�;Qr0��O�1m���9=�9������������{�=O�>�����<�I=�&;������={췼����t=� ��k ���y`�Gn���"����k-(>��>�T:,=u�弣�S��5�=�>�ͨ>,!��%ý&���#q����ʶ= �&=x����%=6��=�}��I�;�ࣼ������<��>P���i�<��4���ҽ��1�s.�Y�&��2;�*K:墪���ս��6;����ϼ厽��=ż
<�z�<�!ɽ��>�)�OV|=W�q=;<->h:⼾_�c�=,�F=c=�]Y�ƾ=��ڽ��#>�[�>��=�1��3�콥c��p�ڼ�'>�q��oн&!3���+=��Q����<�<�>�=��=��<�=���<����reJ=p�=fܻ��$>��7�>�n)��S�=T�>d�w�cs%=�1�Ӏ����<��9=��;=�/V> ^L�_0�=za/>���=Đ�=ɔ����<J6+�n��<)fc=ǘ��*la���=��>X༽��_>"�=2����Z�A�|>Z�O��z3=��=iM>UՆ<q�����TQ�=����~"�?�ݼ\�=隴���D��f->�R+�������C|H��
�;��:=�:�=y߬�!輤�+>7�������<{����;�����X��>�=xE��BN��}�,�d�$��<�|�=VO��'l=��<�T=�@�=����9�J��!��OK=G=R�sZ���-Y����l�=��ٷ=Fuս���@x����?>����ǻ���ԽE�=Jk*�{��=��=h��a�[l�<��A<�C���գ�ﯢ=��p<����g��E ;�[=8���pLp;�=M���[G=���sG���<��	>d�G���:=��>$��R�Ƽ�t=��+���Y=�P���d���;�%0>2�B����k�Ļ��C���8��<m�,���~�ⵑ�ƘǼ����^=��U<�n+�V���X�ݼ3�7=�a6�+�潫uܽ^�:>�+����=��p:�)̽�(ؽ;��=d�=���́�<Q����;���<$&�������|�q�ʽ�	�;�G;�*�"�7�ۄ=R��<�9�p�\��ʘ�m��;�Մ�)��=��s=�a��4����<�I-<���A��eY_<vc�=g��[�=��=�$H��&�4\�������pP�3��=)E�[��3ú=�����@�=���< 	�=��彯P����= ��<� ��&;V����.����V�ֽDM����<១:dn�=H-�=H��=g�=*=>ҶP�3_�<a������=��(>ڿü��̼�����«�ׇ7���1=�f=>���<2����<��Y�)	�=\=���;��9�I��"b��#j>KU>�u����=D����`���=��輬(��C�#�=M5E����1="^+���5>��<�2^�N�w��&�<$U���O<l�g��=1 X=�*=
�y�Q��<վ"� V�=��R�;��=�'{� �=l&���*��1�l,I��?�=%V�u>���P��X�<�<�qj��G����ؼ��=e�������3	=iẼ���;b�<*=qt�=���u}ռ��O=o���ޑ�����K��K�F�'%�� �=߳˽�w��@�>� ��$�P&��K��=�L�=�:�Q~�<�]��a=�Y뽵����ꗽU�M>+��=	�����`�= �<���Rw=Q�0���ؽTY�=���=|�7<�#���[-=+����佯ѳ�%uS=@S�ҹ��O�<Opn<��#=�j���h�=�<��/��j=Wl_����=E��=�)��|q�<�ג����=Sؽ��q=I?	<��=3 i<;=�4�n=!o*�	�G=/�Ἕԉ<EY�Iký��=�!�����;�g�/���t=[��=_ȼ�r*<J$�<�
�� 7�9ô����=�7�;���*�Žk�=;�<$��=v�#<R:�<2���1�Y3�=9t��E�=ƴ>x���_,�W5K�#�;�:>v� �;�='G�<�=.=T��<L���&�7��R�Z�x�&���<AK=?ņ���=)��`�o�<!ّ=Bj�=ͥ*�A��=��ؼ�p�V�=�7�=�f�=\�������8�=�G=�	���
�i$�=H�3��=OE�= [.=�q�=d$���?�<2:=)Ɵ���3���T�2a�� >t�-�Kǔ�z�R=�\P��	<�J�=�n����=z�<:C�����`�i�ʛ���=)ZZ��܋�d��=9=aI= �2���F���:=�W;�AH�<R����ǽzd;KK/=�>x]=�ݤ�J�Ľ�U�=���=�޲��\�z�):�Z>f�`=� ��X���[�=��������<4�߼*Y<Ǖ�:L<ө��N�W;E��<��˽ao�iį=.7%<}z�=cW�+J�=i��=Td�=�MN����B�*;�^���5<�T�<��\�;z�>�\�=ʾ���ǽ=�]�=�3i��F����">-����=�Ƽ��&�#>��>)����(���3�=��#��J:��v���F��G�=�2G��C��Y�9�Н�<K}-��ý�/-=�Q��r�˻M�r�
�=�*��g����i=9���M��}h�Y��=2ܜ���齊��=tM,>���=J�=���ݱüQ��=.J�=���ZD�&���|Z���}�;R7<�۽�k��S�c<e ڽ�ZQ<�P�������=��=���;��P=���<Q�Ľzm;�Wk�=f޼�����&���=�� <W�;��D�ؓ<�D���Ͻ�*F=�=%P�<�Pv<�x�=���=���=`���%ʌ=�R�<W�=��<����!E;=�A�^ڼ�����e���<"+�=���=��#�!%�=U�>J�P==��D� �=5q�>�՚=��M=��˽���MC="MU����=��/�렍�5>�=��5=$_�=d���v�=�$��n�S���5>X�<{8�fϕ=n��8�9���ߧ=��2���<�������^<>ۗ�m=�`�=LZ>N�#����b��	��S����v��G��<Z�2�����^Ga>>����1��<�V��yt<�#�=_N=��=N��=˂2>�x�=�_=��⽸�
=}�=Sy>��<�l��=�*�=�Լ4��<.Q޻l���8�M�ܳ޽l�=����_�=�p��m�=� 
��^=vA<�������<?��<�?�%=��=�-��@f���9=��=pӵ��#>��5���&�j}�>�e��+`=z�=����ԥ9=Q�3�L�F�����h�	���=�P��̼�]���=.�=g� >����g=�	����=�Y-=����Q�D=n7=fD=����p$����;�@�=x��=�=�1��Ԗ��p:�O	�<w�<:/�"��h#=�i�<�o7=N����G�=���=��]�!-��[=��I=]?�=��">Y�N�<L0�=�<�='3|��Z=�����{�=��:�D�8<�s�="~�=ٽ�D�=@)��� �c�H$'<�I�g���_�JKy�q��=(`L��<]��=�&=Z>�u�=,u��x>y�=�~�=�����2�;�>���=�ic=��Q<�;�Ŧ���=��_;?�;XM�x2��)b�ѻ<b�D��̘=�n,�n�<wG�=��h=c@=��L��֑;X�=�i�B��`�ϼ�b=<�<�Rn����0�>�V#�k��=/�R<\�=J�=����o��;����%���<-JL>SUe��+�F�3�-�P=�J=uc;=�|�����<�����CĽ,�h�f��=���<�+�=��J=K}$���#��:�TY�=q<�lJ!��=#�P�4��y��;T¼z(B�t�C�ATA>ӯ�<��'<�M�HM�ٿd<|�=��>��v��ݼwU���ݱ;g�2�ɽ�fy�bl@�a��<w�<�,�=E��=�n��kA�=�P�o�Ͻfh9�/1����=c�=�
e=�A;�禼F��ۜ�=܍׽bf
�S��=�s���=����A~�<m��Y��<�&�={�1=Jf.<��z���>�����-ؽ����6Ҕ=�7=�>pЬ<i��y��*k�=ń=M��~�;7�{=$;x���=pb=:Z�=o1>��5=ئ��^J0=���n��j��s.�<؇߽��.#ͼwdV��j&�*q>&���/ئ=�	�V.�Y�����,=)%5=6�%��҉�ɾV>�ޑ=q�����&��.��}�*��'<�G��� F<�T��OH�=���5(�)�(>�T=�$�u��;��ǼL������=
�7>;��=���=��Q�U���s施�L����=:��=;��=B��p�ݽ� �=ꅃ���j=cH�;� ��5>_!>u��;�5�=�g5�)A�=A@E=̽=�����y��x��<Q�+�:w(>J�?=,4�=E�&����<3�*�>�н�x=w�P>oS=}���⹽FD>�0���4���2㼸�9Ιȼ�
�:L�=��/<�^�=y�Ľ *=���<�\0>�f�����=MҔ=�B�"�<P@Խ	������K��_y�0�N=q�-=�"�2�<J�������w����`=`�9=|��;��i=*|o<�I=:�"�t&�;i_��1���p�<��c̛��ԣ���^��^= ҁ��Ͻ���<�h]<�����=�d;�MŽQ�=y�<귴=O[�=Pu���Uh����O$����=ͨ�=2U$=|��=9�:�5�=��\=/H�<��ռ$�ݼ��=d�<��T��+�=���;�)	���;0����=����N���=YN�s�%��g=�qo�}ɝ��a�=j
�=��~���r����<��>P:�zO�u�����<�������=]�*�>/0�=̟/��Ž��DDr�ǈ;��7�ٗ=$��=���=��=�Z e�b~i<��q<�6���>��Z�B�����9�v�m=�J�<�=�=�(�j�p<K��=��p���8,������R��=½�Ă=D���̾I=�O��H���;��E��r����=�a ; \�c5D�!$>BE�QӲ;�,������=�= ��V��V����=̨�<g��ݒ�<�5>BC��y�=���7��=A<tb��?ܽE��#�<s�U��+�^��Y9->��	�=|��8
��B�ؽ�;=�������;ǫG<I�=����` �h�=���;M�>��gE�'?=!�<��=q�<H�v=(v���r:�>W��������<F���ݽ��g��$3����T{J<�j���I9��yG�߾=�S��m��<�
>�G�y�>�*:�g�<�>Y
.�?Wٸ���=�μ��Rɽ���Z���E4=Ԃ3�T3=���=/�Ž=�
��C���K=�Wx<w�>z������.>��<g=�ը=�u;�ϖ=��1=�_�[N���z:��┽�������x66;oٺ<o=r����!�B3)�V`a=�%��uz0>I�}=y:�<�7>Jn�<�{�=o��=��<�V�=O=pS*<w㏽���åۼ(��= DG<�P��6h½.����p���M�"d�=#���=nx��:�����<�G�;q������׿����:�ƽkKA�)��<�_<Ε0;�X�=k��;�$=}���X �=��=�=ƷS��K>w�XЄ<]=�=KY�=��t�J�>ۜm=�:'>�T�=O�н���+M߼�۳��!�����x�=��M�������b:��<㫍��r�=c�������j{=���G���Qr��l�<B�E&޼12q=mże��=w:���H�v����9���=�P�9�=�س��;(>�z�<<%�;EF=����tE�<�P����Z1�=�C��$>��=>h"���D<���U�<=8O��w;1�^>]�<�)l��>��d��t�����=�l���nh���g=�7/=nK�=(�>�Lk�=�1�;Q2�=M`>J̈��������W8�id=���<����!>�����=!ų��5�{�ݽ�^z��'�=]4��:}.>]�=��`��KI=�?
���j=]�x<�R ;�i����=���=G���"�=Az-��t�=!�<jZ~=e��=�� ����� ����)>�=!��FM=�5=]�����˻�U9<��=��Q�E<��OY�< %½��-�0u߽� =�΅=�e�;�x��@n=j��=�~����=7B�=�*�=p��=1o�fx�ӊ��X�=��Q��n�=Nv<��>��.�%�2>��u�%$��>�������><�����;��=1�3Y�<��=��NW��н��{=M�/=;�j�,��	ꞽ��=If���]��jn��S:�=����D=�"�%>�4�����0̘=�7��JD���G��X >_=�нP�[��Xn�"�=�&��m��D��=e�.=�Y�<u�< =:c^�{$z<S��=��ſ�=9{v=���S�S�{Z=X*�=T�W���z;�D�<_;�V��#=<Y�<VQ�����^�<�;s�Y՜=C��=u��=Hs��Z�=l;y=p[�=�D=z�=�I��C��V������=j��K��3��H��<;�r��>��V��<��{<�{�<?��=�?�6O�<�?���;����佱�=M����[/��]m=�����>T�=�1=̘�<\��:�ً����;��#=*�=cܺ���G�ľU�e��,F���ü+�<�$ ;8�u�Bj����8=�7=��G= �칀!M>�?6=/Yս,2B�g�=�G8<�>ҼQP� 5��=\�2;|ƞ�p�ѽ��>Օl��E>=0`��Ɇ�f��=&��=L�_=I޻7E��"��;�T�<[I ��k�=��Ch�<�ߨ�ALi<Zk�<�1ͽm�G>�E;�)�=xqT����F4<��[<�)=̍>�X�;���>����^.��R�<���=�=D����ս"�=��=�ӼГ��E5j=7S<J�=	bc=�K
<�yu����|!]<������<I�Z�L��=�PH��>���&�	�'������=aF7����H�@��rƼ�k= �n=Q�A�\
���3���]O���F�<�5*>��<c:>ekz�M��'H�;ɑ}�fc���<98�=�}��z=��x�=1�>8l��nj�=�놽��7=��z>0/z�!�=.�黝=>3�:�}�U�+Wz�(�=�.=�������2�vj���m<>�A7�F�z�ӽ�r��*pĻ�#�<r��<e嵽�7R>���=@�<�>�k>݃=�QR���g<��<=(�A;k�=S!e�g�Ϛ�=Ĕ�<Q=隩=s�j��B"=��M<��<ϖ�;X��=;0B=Z�	�&0�=(��;et�=�dd�-+��O�=�Zi��P�=j�P=����\V<�ꢻ�E�=4%�=���d�=�����QK=F�y<�!Z<h���5�=/�`��:�;�"��1������/R�!�]<`'��I�<��7<.L���R��x���=I �����fE�NO=����𔽸^����P�����"=�:<���=�������='��<ah����ő�j�=9�Ľ�\�=�󽺊�k�=;B�=��=A��=^�D��1�=�@�=��<u��<�v���T
��
۽n*f=�d�ڂ
>!�=&`�=�S�=v�����=�K�=���;'��=�ݼQ,>K(�;����?�>�+q<ڵ��5!>d��=`w��2J����/=���;����cI�g�=6b��ך=(�$<��6��%"=~��	����=r�C>3�i=0����<\Gz����u�=!=؄<��.���>=�F�HSX;�.��>������U���ͽ�5̽�S1=D�9=��=4�6!���	>#w;����U�=W(X�k(Խ����97��&�����~��x:<`b�=��<y�4��Kl��D/�/۽�=x�̼ad=['����c;+��==�<x��	�>���&��D=�,-�=Ւ=H��<&eZ��8����\����<��>(���Q�=3���ϻ�5�[�=�=��>��|���;�ͭ=�(�=L�仐ƞ=�˻=⭖�&�>�o�<�<�=�������(�k�̽6  =�?O=�p�<�9�=��=�뽽�YL=�r�=��~���=s?�����PrE=����C<��`�=NC���<;g��X�=Jߢ;��ؽͩ':u������<�D��Y�d;~H�=q�<�RY��La={񩽙ع���Y��@^=���=��ܽ=t�����$o>��=_L?=��=����3	>󋘼m�Ƽ�1">x`��g3��4.<�sq�$>wcX��NT�A�x��s�f�A>���1�;��ý#��=#|����]�N`�=����J���=̮s=��<�h_=`#���l�<�H�����W��=/�@=}�����ʼ�J5=X��=]� >nb�wʎ�3.ɽŢ�;�$��Dk�kڽ�!���#=W��;��=)��=K��J��=/@��0.�=m�<?�=��߼�=���_��  �=�'�����=�{=��<#�^�֩˽�z��_d����J;F؁=��L<��<l���ߎ!><�w=���H�Y=$L��f=a��=�1�<p�L>�*�=в����u��B����=e?ѽM��Ή�ݴk;}T����<<�Ľ+��=��\=�<
>H���]����r�q"[= ���lI;
������=F��=�����꽨�Ҽҽ��D��<IO��ϯ=y=1>������
̨����Y��<(��=�8�.H=��@�	=2��<J1g=`�۽�>���Z��ӽ�=�U�=��x=Q0��=����:YM=��^>hY��ż�� ��g,�7H����b��<t_x<r?�<}�z=u�>���򺼞�<�S�=� �=\U� i(<�SL�aE=Y���W=���!t(=s�:�g�=��ݼSd�Y�S=� ����R�]���m��Z���φ=M���ٮ�_m�=���:��>?C�\0=���=�P=�'=˯ƻn���=����F=��=b����{Y���i</p=�x�=]��<�{�=�Q���7��)��z�=�� �=�Ƽ�J5�pm���=���<d�&<Ƙ���,�q��Ӕ=���<�J"9E��X�<0F�=�">g�����[�g�N:���ݽ��{<M?�<���=�ހ;dr_=���p�"�ڬ��lZ�6�`��ݽY��G���u�;>����u����d*��G�؞��=�4=�g��Y1�<I>^�ν��>3����xj�&zY�����1�<�Z�<_��렽�~<ښ�>??��(�=7�� ռ/���C�ڥ���=$H<'�����^�=�<$�<&���X��ģ�1�3����<(��y�=��j��y=���)�b���=����v�=T��S)��O:�]w�uz=���L�b=;�2�6��=A�[;l�=�N��X�>[`Y�ڑ�
�&<6&=_��E:��O�����'=�鍽�+��uG>����=�:=͵:��N�<\᷻�b�<#�)��g�=�8�=s�ͽ�`�<W���Mf޽��M�R���:�S��&̹G��=�	���<��Ch���
��=����Žq��=�t�=�А;E&>P��<bGĽ"g >�̂=��?��P�<?Å�$Ԩ=*A�={��=�>Á����3=Mo콘��0�;���=��.�s�	=u����������g>k�=�	L������E�<W�=ގ�;�\�=�N�=Iv*<���=�*���S �����j�=��I�(<�nf�����
킼r{Ž������*>}9�<2�Ƚ'~�; �p�=��5����=�?=��4T伋8�;i2>j->=�i�;�8<���=8D=�J�x����9'=}��=�������<������D�-ތ��1�h��<`� ��ˣ�AY>[� =+R�'�=�
��l���v%=��)���Qz��x>qͽ*�z|��2>��ɹ"��;�#�:����ר�<[|�:?q=� "��p�:�Jr����< 9Ѽ��<�b���O>�D���Av<^%��Ì���F>�,���vD=�]=V����=�]=ˁ�<ax��΅�="�ܼdE��=.ʓ��?<��L�V��=2p�=a�<�����	�;���m�=����)<7���/�f�=��L=�Լ=2Rg�ǋ��
�@<�����b<�h��W��<KT�<��<�hI�\��="�Z=��<A��=,3.�C�RP��QO=�>"V=˪��� D>�M�=l	��@r��=O=tj�=�I�=x-K���G>���<�B*�S�bJ�� ^��c�?=�Ί�M�=��>>8>��K�V>$��m<f.�.�[=9"ۼ
�=1I�"�k<��J=���=��=+�;��<N��</��!�</�=%��X ��M�=e�~��mR<�ʒ=�?=�6�<�~ >�޼Q�ֻ�ݿ�9���F=Q��=Ey���竽.S�=���6��=H+9=;�ۺA��щ(�e<���P��ӏn��R��AQ�<w/ս��=?����oS��W�=���<+��=0�N>�\½�v�<�����=�!��(=���=�̝�%X�)1����<\Gp=�W��F�<a����<�d>��>=Y��<!�;�%��=����*o�=�U���%{�#-�<���=�6�=��Y=C���E>?��<�U�!+�={j�jؼ�W<��Ͷ"�ώ<�Q=�� <�%���=��M�!)μ��OE�S��<�����N�=�,�'��)�=(r)>%�<�o��/�==�z==8�<�?����;<|�i���r�����^=��N���=��h�0p[����	=�ӷ޼��>���<��=*BI���I=�"���~��;��B�$>��>hۓ�X,)=��<�/��L�>_��;!�����=V'����=��a=���*��=�;����f��e�=QV�=�+�=���	��_�=��L�����=�I �e�����q������缳���ܽu=��a<պ�=�rս��i<k����Z������Db��=�=p�<��>&`5=��t=�k�<������]O���=�5����ܽ�~�y|Ƚ���=ٽ�tl<�R����0�<>[�P=*I���8>��x��/���==�]�۪�<�T�GP?=C	�<�q��e���W�{�=�s�[�ټ��85��1��=��-�N>� |��S��o�=�O=�N���@�^C��O�<؋��悽�gm5>l<��)<bi	<��D��j=(hμ˿ܽ��T>��Ͻf	=U�<����.݅=��e��'���\��O��=s�H�^jY���=���*v�=!�!>�!��[�����=���<���8�C>u��=VR��k��->k��<T�P�)�ɼh���R`<���F(3<x�= GZ<RG�<4��rA�;����'�_�h=�����	�L���lY����Ȅ�;���1�ڜ���Wp=;�c=�*��ա~��c =夀<�uؼaw�=&W���	�<���=��=�K;�ͪ�Ae����>��L=- -�k�*=a��:��<�t�<�N$�&|�=3V�=���jؾ�Od��!>�� =��=͘:=�'�<�d,=�h��
>F-��p���;�~��?�=���=��=��ͽ<m���Ȇ<��@�d�0='K ��=�e�=]W�;�p�<?Ě���<I.�|9f<1.>��ǽ�����<�꽐J{=��������}�f�r�Vs�<=�@��P>��ɼ�G���lm=�Y���7�<t&�<��Y�Ru�=��ϔ<��r��p��>�ѕ=����U�<
�z�e���DL=����P��`�=ݢ<��!_��ݛ=p��K\��U?ڽ���f]V��՞<��>�Y<��Z<�N�<C�ʼ�/=��!��B�;?��=X)���m�<�`>^��<���&S=i�轭��<f����B<2�B=��Y=�J=��"=��,i��%��=$�F=��Լ�Q�=9��ݳ��;�@#��ܓ;o<m=��=�?�=���K��9�4Z��g�<)��ʿ��O�Q�弰Ĝ�ȭ�=�R�<�Ƚ��s��Q=���G[:G�d=�:�=@h4�k��=e����¼2������=^����5t>�F׽ �>�j=@�=����1y���]s���\���ٗ>G)=�ӺP��=��<�������W�;���Z�
>&k�=ߜ:>��>�/�=��=�8=�M@�Y�=���<�)S��Vݽ�ű�*���e�=�ҹ=ߦ >�ֆ��ڽ8��<��=uط�O�/����=��=�>���%н �
�+�r+�����C�=��νD��u�6���$=n0/>��+���ݽ�o�=�`�;�Ҵ<Pˏ;͊=��9<���¢�=;�I>�q�=��=��)=�=��i<��|<���$�x�?A�=���=��ƽF���">񰂽�"R��Ü=}3�=�\<�<5YJ���r<�CJ�L��ʜ<����7*
�Ե�=�J�=��=��<���=�v���?>V}�;6̬</욽�1�=1,;@2��m:�=�@����6�0��:���=��
=��9 �>'�3=d��<W����3����R���j�<W����3���<,���.�����</V>��<S�>�ƀ���=W�6<�x<P4]�ل�<ttȻ��=iTE�s���/�/X>bd,�������<!>=R�>�O����H
>M�Z<s�弹`i<ު���2V��\:����j�x<I��=ѷ�ؠ�<K���>���`�=X�==�s�x��=侍��4�F��="ս�A�= �U�T�<=o��=�CR>�=D��=�>�������H�'>ED＇창�_(=���=����q��8�<�= >k��=z�L=���=2?�=���=�:ֽ�-s��k>����k7�<Nb2���;��̽6����<#��=A��<F	=5;�$�@�GS���	>��=�t�=������R���(�>L�O<�=���=i��<;!���=uA.����<!潽�;��E��<����R����<E���/Y��Y��^҉�-寽�K��=��<�4����r=�r=�Ƚڽ]=[�q=�+=��C>���=�F�=o����&�fH=b�%��c��4�D=��yF'>L�����=���m������d=�+�<�!����$=��ҽ��� ٍ���=y>�<X���D�(<��]=@\<�k;m�޼p��=�+��6��$�F��=f����p����=1U=��{=S�=�Z�=�Pʽ�Q<ԙ�>�	���n켔kؽ%���>j̽0_=>`��eE�kt�����*f=H����ܽi��	u��
 ���܇�����\=����v>��H����J:�|��<!���Y<��<0�=u��μc<"$<W��=��W=��h=��*���}�=�<P��*;<�Y>dԏ=�ߥ�t�<N()=��=�ż͗��o;j+�;*v�s]=����-}>�ߖ�6+���ټ����l�=��ӽ@r��0�=}M<a��=��>1
�֦�<���<��x=��d<ꎨ=��3��z�����=6~��3���� X�<��vv�$��=q�<M7�4V���ʦ��r�=K������=ƾS=�C~���<��u/ռ(Ƕ��]�=��5���}:��=����%�d�tN)�����L�=1�׼1<ܽ��=��.��f�<#���}�Tr�b0W>9u=u&���<l�=����\\�=�|	��&�=w.;y>�=��q;��3�"�="$�&���ż<.<T��<�ͻ@&B��=(�%�@�a=WW=#KG=>X�<n7*�_,J=r�彶A`=��L=`Jm���=�*�;�<�ּ�7��-XD;�Ka=<�v���;�=/���;�=��s���]�0f��
��M_�<�-g��9�=�O_=������<�}�=�/�=�@�=�J�L�=��=!p���B�=�Q��1������<�μ���=��C�L��^yɽ�` ���@=��p���(�K6���ر=˲">]�E=�s�=%�<l�h��{!��m�<�=M!���;�fI�^��=;w���r�F��=��ü�Z�=����"=\j�=F#�l.9=�B<>紏�O(1�&B���Fp�@~�=:�>�@�<���Uv��\,!����=���=��|���:����X(���>��ĽNۇ���-�Ƿ�kmŽ[�	����=����d_=���Ӽd�S>�����$�=��i�ݳ�<��>>᩼�̂���f����:o�=��x>��S>Y&R�>�ͽ�~>�Bd��U>��+��1��aĿ=R�T��@�;�����=oY�=�6>�c>=Q���g��2��\⠽��5<�j��rݕ�W��<xGb=�1<��=U�ὧ�H��ss=�@2���j��܃��X�=2�Z��=l�<|=�.��,b�����<��̽�˼y��<H�K=�|ϼ��?���[=�{ȼu��;ē;�Y�����k>2�B�"a/�\�}�5C�<Ɛ����5=n�)>7�k=�ݩ=�88<VUn�y��=��=X�ͽ��5<j�r��-��$%��G�uu�=��>��=��ý�,�<�bǽC�=���T	�Q1���Jx=8c�<�F&�eZ�=`߽[��<^�=�Z`=ַ5<ו½4�g�n3��#<e��w!=LZ����������n3M�ʛo�����<�P='|=��$�fI�=Sv\��<��3�=��<}� ��-=�����W�<�Jk��'����	��VL��=��=p�ܼ��}��.��V���>�b�y�a��=��=%�c��҄;�6O=�ٽ?C;�Tp�]sK<�!:=�{M����=���<�'�;y��"��9��0�\�3��L*<+K��4�dv8>L-�<�ֽq谽�J�=Iv�=��<)�8=:�<Gν�2>u��=��Խ#��<Ʃ =K��<ds�=���q�5>��Ľ�+��/ǅ���;�`�<�'�>0��l�\�(��˛=2t=���=�g�=XI=�Qg={���� �T��;_U�=�����=���E[��ѽ���=$��;;wk����;�:G=.K>Y��=�2�<�!w=᳼=9�j��RM>]���7��6z�K��;&b2=8�t����O��<���<K:J>��-=��^=[ؐ=��>�6=�>b�=�^�=dh>&�g�2�=�.�n�,�-`�:�7=�H�=��j=u�Z=��=n�=�v��_�!�lN3�rU�=8,�\J�)��= B%��د��X�=���=�"�+�>;n�T>��.罓�\�CU�=��3>��ؽ v}=u�0=X�=�)=04 =����ɪ��χ�F�>�z�<�B)���l�=N�=�#�<om��ɞ=F�(4h=�Ș���E��3��٭����_(�=��7=����>�S=�j��b$⽻?�=�р�_&�=U}�	�b��e�<l�<��0=y3���j�=LX�3iK<Ӕ�=���=�e>�h�=����
=fv<<+�W��>��߻<�S>UJ�F'�<tV<!+r�R�6�!-=��&=ͬ7�7Sq��Ǽ��6�YG/<�k�v��r[�=}�=< K��3½�F���r��A��=nL����:�p�=i)g=µ<H����<�����&��%�����lJc=g�[=�|9=���YX	�k�)=v7��j'/>���+<��Њ?>#ߑ<�c2>��=�C=4���F=`�=V�݆D��N��=�O��u��9�	�&{,>���:p���l�-����@�<���y�B��B��/�<�����b�<���=i3�;<#��أ:���D��ǽ�4��&>Ŭ��]�E�D<9� `]�eL��d��V��=��;��ὲ�P>��뽉�=Pv����@=��->�h�=��"=ri�=����==��=�R�;뜜=��ۼ���<�=U��D_=�G��.�=_r>	����5>�������<�=���FN�u��=tDQ=@�̼���<���<�>=*%��E௻2�r=�=�9=���<,���;W/X���=�l=�}=�
+���h=k�;=�J>�9>!_��B瓽H֝���ԸȽ�=4��=uk���J{����=�l=n�������/=��.�q=�_/=�VD��>�=�r<֝��pX�>ߜ�=�Q�_�->\��:��h��" >B�ϽЬ�&�[>���=�д<y��ul=v`��7ͽ��l>����+G=�&>d���>5��U�e>��ֽ��=c8�=*��>X�b��A]=cU�2i�<�4�=�q=@�R���&�@&��X=�ks=*m콧��=��R�i�=�g�<�ַ��&�=2S�<��=TX�=L�i�C�Ȼ�o�=��:��<9U�SM��b��a������X����(�zj@=iy6�q�<g��=vΆ�����sy߼�� =[/6=��c/=F̿�����f���=Nɽj����\��A��w�<&%����=���x=B'�+򣽉�����d9��P[=3��<��v��z�=��n<�L�<�֘=jŒ;���=ٞ�=��(���s=����R�=Ɵ��rc��r��=~�a<�f�=+��=�H%<�R	>��Z<uF�<�G��I�<�q��6V!�/��=��q<�����=>ꦼ��ý?�E<��;��=��Ļ�%�T\�<�{����=���=���^�Ѽ'SR=y3��*2�RɽpqS=-ճ�~�=3�=Ќ�;�IC����\{&=�,����=��xL�p�'=���:�9�;���=�0��U�=��<ф�<X���W��=j��"c�SE�;>i�<��Q>'����A�A����S��|�ț���}��Gֽ�-���y:c8G��T$=�I��P�=C�?>ر�ɱ>�Q�=x�˽0e���.����<<����9��<�ٔ=u�=��.=�J�K'I�ӹ��L9�<�=h���4��=ү��Q�=Tg�<��=�r;�򽽴]�=!Ƙ=�W�*E>���=K^;��=�O��hP��h��.��=V0H=��<dq8��7P���.>���︵=B=u�����~�]=T䖽�v�<L��=0P<Ol �>�N��=���=�}����=�ָ: l$=$X.>���=��<x"���1<&"��<s=Oy'>��ڽ��U���=���=��'�0��=��=+½D�D=��x>�����Ϧ��*>3YT>���������>sZ>����X��k@˽&G>ޠ� ^�R���5�=��)�V�)�;<��p��6O���=-6|>9��=��j�]�Z��8�=L��=�S=#=|Pǽ1O��g�_U5=�+�='㽚L;=>
>�E=��Y��0X��'�'����a=��ݻ��>�=Fg½M�5>���=}����G� �ׂl��������M��=��=~E���xI�[*�=
�r<�
�< Dk=�y���q�=e@�]Х��zo=�[;c�<�7�:&	7�R�c�i�：�)�������ͽlҎ:R����e�r�<.ɵ<Jh�����^F=vBͽ��};��<����/; �A�"=D>�7��V<_�o�]�;W��"�=T�=�O=���="��=ʽ_�	=��=�)�z��cy#=�V����5�q=J�=.�G=�v>��d>�m;-oM��ع=L�#������;V��}T=��p���=���;�Z�=rxu���\=�}����= B=z��<������<
A�=8��<s	=y=��=��y<h��=0�ݽ)7Y��b��Y�_D=�u7>��>���ys�<V,��[%==�]�;�H��>8>4�ƽ-g�%�U�R�,=�Z:��+ڽ�Q	>�р�M+�=�Ȕ==)�_o�;��2<�=>��3=�qŽO����=iPY=ϮS<9����<����;>�弄�=���=2���Ȗ=�!=�#��A��<��d>>�ӽ���SŽC��M�>��<���#�=i�t�� <=>R�<ip���<�r=�M=;3*=�a=m�`;����;U@�� �=����do��8=�v�=�A����<�V�=a�=#=��<t�*��VI����[��E�;>աK=l��=�� ;W�m<�)�<&ٴ��A?=�Dz�&I�<^�｣,�P�=$�����=��<[��Gթ=�@�_�=���=2�M���=Gu����c5�=e(��`U�<(�Ť��=~3�Ÿ�<9�l;��m�:<��<4P��l�=�r���M=sʺ<�#�B7�;2�>���`�� ��Ӏ���~f=�=U]ݽ��;U���?Җ=m�½1x�:����EL�\�=>��ʽu4����<��=qQ�<�Wb;A�=�\�=;[<~W�=ך��kV=5[�=9ω=.2��ŉ9=�~=�P=�/�3��<yɼF�f��(S=�ۺ=t����6�����=�O�����=4σ<���� �K�)��v\��ʅ�_�<6��!ek=']=NZ�<���=������=6X>y �g��=��䞮=�a�=�F������5Yڽ%�=�h���d�<�ӌ�n�+>ЛD=� �<��c�GC�;�6>꼕� =�=,==�[�H��=��(<f)N�Mm�<�|Ƽ�y<�~=#�}=�Q���
�<T"0�T鞽X�K<�1�=�ؐ���i}����䧇��+=d/�|Z\=n�*�������=]�<ط����A�('=�	>Dýc�����7i��M睽�K���
��!y9�h�=;,�=��=.�-�F|>��l�o>���k�<"��<7�<���)=@��=!�"��9��"�`=P[=jTẀ�>3[c�5m<��H��H>Vs>Ц��DFm�8�S=��8�A���3<Ͻ�3=O[�=Rh�=����m����.<��g<(�｜>ؼ�"ؽ������U}���.:=�����*�<V��=;>�����J�y�����/�=�p�=V��"-A���=X��:�e�=�;<����?[-�c�ֽ9�Y����=\�g<��r��=P�<M��=�m��͗��
���;�V�=�A��y�;���=\~V��\�<�R�=o�hg�� ν���>��ޠn��U�;������S����I�<$��=��<��=V�a��<=����
ȽW9�=�>
:o���P½4$����8=�;�=+M��<*�;�
>����C�k����d8=�q�=?���>���{�DC(>J�P����XO�-s�=���X�I=B��=9�v>��t5���-l�����Ag<߀��Pj���ꑼ�����
w�f��?=������=��0�wv�=�6=�\=� @���� �=��x�4�̽��->V�>>���b:��䟽)A�
7=*4���V;�W�<��=	��=�aU=���?Ѽ�=S=������<��׽�j������)�����b=T��b�<�e=E%D>s�SNQ��@�����W�Ƚ@���`=�6�S�=v�< [ؽ��`��C<�뗼_b���ɽ��<V,����Z�C�=����;{�=��e��s=�-=�1)=)C =g3�\����d=�C�<Hj���,i;��z��n�=��L�&�ѽ&P��_�<���ʁ��r��#�<��������Oy=�׼:i�=�8���������%�=��=�E�<���=��=���=��jN��Yy����=��=FF��/��T7=�;����7�ltd<#<�Ąz=�31���=kɾ�
ʿ<9߻ �=�@a�9�H�x\���1=}��Ԭ���޼Wr�=�Ď�J�������)�=?z=����׬�w@	<�0�;"��=0W���U� ��$�=��=m�P=�=ԥ0�6Y�/��=6�l;&����K����;*)9=���<��O��s=��=7���Z=��<x�,>[T<���F�TҴ=����ݐ=�>(*�=��>W��7esH��e=Q�+�,#���ʻ�놼F�/=[�̽Ŭ=щC��x�=�\2�<��<u�=� >:�N����<�D��	�7�b�>��=9oY<U�ºw�(|�=Jc���<�Dm>r*��=��m���>�H��n�<���=(,���i��A�<}X>�.���,���W�� �=���=�q?=u>g=���,�q�½.a)�!�E>��S��-�=BM�[Ͻ���=�fI�"�=m��=^6e=��7	����>�×=<�K�%�޽'O��sq5>�ͼ$D��1��=7#H����=��=96���@>��(���񼛡^<���=~�*>j��=� ���ꞽ�Nf=k����[=�e�������>\a�5x��X� ���ɼ��Z=�&鼰�=�OT���'�V<�����#�=n�ټKi>k�=巙��������і�b�=z���%�=�"���mj=W�/�>�i_�=�����4����D���ʐ=)/>�K��zѽ�rU8>2'��#R>)Cѻ*���)\A=��Ƚq�2��������=�AҽNBW=�X�<U�k;;�=�� ��d=ؔ�<%\����㽤7j=��)>iO�=�Y�<�(Z��8>����Jq����6=#R�=Q[��|rl;y� =�p���q$=n5�<�����u����<\�	��ҧ� x���n���c<��a����ٽ���=)�=c3�8�S���j����=�ɽ'!�a_5;`{=����`��
�����<��<�?����=U�����=W��'����<� >0��=0nZ>F��b�ʽ��!���-�H��=��%<?ɻsU
>d�<�Ls=��&�TNH��_a�Y`�����<͂�<�G�=�+>�x^<%��=~��=ŅV�\��<@,r:�J1�� �<�u�<�=*,-=��>��ٕ��枟<E��qx<ܽ��>T�=�K����;RǬ�2�K���;d=l�l���=��u�=5%����=x�L=S�e���8���a��+&=���9LG�)���{���5AV=�u��b�=�C�=��ּ��=,j��DGs��������=u�F=���6E��:�����7>�h���]T�2� >B��<��<ܰq<X�.��IR9-����»�Aý��=<����=]?�=���?ێ=Yw�0��=fݜ;
 R�-��7��9p,?>��[�ו�=��>_���&��=ū� �����R>�X=u�ȭ=}j1=4Z�=Kou��=a�U��|$��~=�^>�2������Eռ�Z:�q)������[�i����0��!���n>)�ӽ��R���$;���<V��A2���w=}.��0�=6?9����O��ր�(��=�� >9��=s�;V;��腱=��f=�׮�� �I�=��1��N����s�(Va�mE�;���<H���؈��
��;<\<%U���=�Sؼ�Ƚw���({=�X�=Z�=H�Ѽ� �M��<,Z��O��n��=�ݼ����[�%���ؕ<�����=�#���p�<���=h<�d�=V=�>F�A��iڽ���<L< �ӽ�϶=�Z=�ǯ���Z=�ۚ<�Uj���C��U���`�M����>�sV��=���0IW�~��=IY���N��Y�=��C�2"=����{�=+Rj�F��<,{�=P"��μ��؞���E������S��+�|��*�;b�V���������C;q=��(�pQ}��{[=�^{��y��DD��
�<��ڽ@l�=�>Mq�=:W���]<��=s��9|���U��ȥ��A�=����\=�UF�b�ƻ�7>�^>�/ｺJ���x�������_<��G�B��=�r��f>����=!WԽ-��<�tD<����h��3ۈ=���<��=���=�ļ��/��ݽ�Ì�`v���=��>U�>�8ѽ�B�'�I=
6��!�Aj�=˄=]C�=𴻻�t<3>��=	4��J��=�S>p�;�t�=��]�+�#>���=�.Q=��"=�̯=A�<���Xn�BC�<����<z=���;�y��|��<�p.��>��$'s�^�F��-	>�2�=[.�0����>"�g=K��=Z�˽��=��v�`����B����=Aa�����=qH�=1=�nZ��}�=& �=k<�p7S;8E��蜽��\��\��;?v�<tv���H*>f�r��Y�=D
�<l��;�W����<��>�=3�����;߆�NY����=U�ʽ�Y>u��=�8�<�	b=H�����s=q�l�ܹ������=��T�U�ۻ�,>�UV����m�=qM>.�(>��ü�+��s=��ӽ�}�=k�N<�j=�a��X<�L<J�;<�>�-:�[ƽ���=������V��9��=~+I9���<W��=#]Y��ν�`ռ"6b�)ǽ���=�����g�=������;{)�=��=#!�*�^�@S^��]>.d>���N��=�x�B:=6��.��=����*䢼��Q�[E=�_��|=�+�j���:>��<ib>�q��?-�<sPٽf�8>��(�w�=_J��(<��=n)����м���<���aba>6u�=�ջȍ�<85ĽSj�v�<��[�x�{=�`�<"IY��i�gѨ�	��=��=���<m�N������c��d0��>��V4=?����ۼ&]>��o������=-�=g
[=�>9}\=�x�=I����=�Hw��,�=^��<Y��=/���jF<Q3�=��=�<=�a6:>���V�滓�	�(>K0�=<=�1�=ɉռ�n	=2�Q=�Q�=v�/�L/�=O̿��Jf>��s=v >W��;T�n=��=rs޻Z+����H��Q&=덟��^x=����՞�=��(=�#�:�ٍ<'�S>���<���=���M��=�h<7;�=�	�=}�S�����NY�]��=�<�q��<���;�������~�=>=� 7�����=|9=��J<׺R�䰿�ڍ={��=��e�_ս=�x=�R&�=��=/��JD����=�Z`=t�)>�j�=A�J���q=�ް=��<��=�{�������=�*��8ӽJ�ӽ�\U�W����E��)�;���=&ع=@e�=r��=���({ӽ���=Hn�-�Խ8�8��M�=7 ���$;`</�;{ñ����L�¬�<(=�&��l8>�+>�)�=��M���!�m/�z���J>z�4=	䭽ݶ��3���V=1
b>��e=�?���y(=��>��H���*����<�ʀ��N����R�=Un�<��=E.(>���<!�==��=s�%��j=�����<>���=ʑ�<ӆ==h*=D(4=���.Ri�� ����6��=�"��K>��=�ʼ6i==$<�޼,K��j[ϼ>�Q}<�����ϼ��;� >k��� �2���`=�{�=h�=��G���:�翼�Q�=�-b<��z=8�ҽ�"���=/�x�7�<h���S�=�E�=�μ�h���$�=)ߩ<�&�=�`ٽ��=mmս`)�<[�ｅ@��R!�ﮠ=�I>���=>,,�ٽ��>=d�; N=1~�<�d�=3�x=�a=��:H���������=����̙��D5��4��;�8��t>�����g��=	��=�N����<`o�=|���d2�<����XU��`9=��=Uz�<B�2<���5��s��<N޼r�-=x����O�=�W�'4ҽS,F�R��<�V� �$;�<�R�=G�<=�OӽY�������+ڒ<:㻽�_�
]��3��0��Y.=���=��K<���7��=���_�>)S�B6��I��=x6J�&А��������(�����ۦ优ß=�^l��&��GR����@%�������׼�야�Ya=W�;Vmν>�<G�=����=�:�=�Gڽ�Zd�y�˼�/��>w$>��Q�_/X<�^���'=��H��)ļ�a�=�ޔ�y�3M���
�	p=MH��;뉽j}��W O���>`�>�6���=�
��6_�=�^���=;�cջwֽxm�;��:=Xr=�>��UC�����[oL=tj*=��Q�܏>��=A^Խa�w�������4U����<Lgh�
��=�K޽(~N�E_=��@<�ʆ=Zf�=����5����"<�h!��Ѡ�X�>�G >���س���K� ���V��L�I=y>�>������o�	���]=�C�=�ȼDM��ؾ�;]6=c�=&�\�l���<<4^=���=�=p�=�|<���=] �J�g=�zܽ�z=��=G�W�����<��;�Y�=�=��or=z�������5&�&T8<�Q���?�.yJ��L�=�vN<'��=~ ,>�^=�2�<���0�����<R��<Bi�=q��m^>�����ͼD��>�/ν�T���.=�'������G���-=�A<��)XP<V7սm�`=�|=Л�;�l��{W,=>3��=�Y���O�;�S=�f�=�Y-�I:�='� ��=ܽ���=���x�E��X=�s����gW�;�$�LV�<�>�S#<�\&9�0l����DR�=��νh`�<���<$�y=5Dм$)=�Am<x7�v1��$�l=i�L������6��L�=w��7[<0q�=����<#�=/��<*����<`N��a����V�C��̏�������y����*=<������x#�.�^<��5�U狽	�z=ׇ�j廻��>���=��=���=J
�<�\���K�b5b����<N�׽R�����=�/������v�<�S�����T4P=��=!B�=���n�;��V=�F�<�,]�i����>���<=r�=,���d��0s��Г�=/�=��K=���~�*�h�
��%Y=A��<��x9Wm>A��:�j��=2,=�׹��8̼�ߋ���2=C��=ع�<�fR��[��=��;�稽@����>�́<^C�=��=��=���<��A=^z��~ 6��w3>sA����@=.����<m
+�Dz�<�曽p� <N��=H��,\\<�%p=��[����<J�=��ƽ��r�軂=��>8��=`��<�~�="9�<��%L�=p�=�*<��d���漁� �������ȼ(6Q�#����>���b{�1Nϼ"ф����!��6�=��+<&�Q�U�=�M<.��<?/�<�=7��<r�=��.�p�F= ���f�=��ǽ����|�=T=S�
;�&>�4k=�i�<������=�a�=1�E<�����A�=뤢��#�夘�Wb �[2�=S↽�è�߄���<�=F&5=f�<=���E�����=�B�������2�����Ȇ<tN��o삽�6Y=u� ����<U�1>F���=����{=���w�<�5�;� <�bK<s�h<q+g�O�=mm��->P$�-�z�n�>�Đ<�>(<�Ս��Dp=N�j���=뱅=b�->'Dʼ�N�=�뺽����<��μp�}=q�O=h�=��̻���<b.���y9�Y�f��v�="À��3�=.嬽7Z��ߠ��0�I�;=ؿ,���Q�R��=�6�=�Nz<2��=g�m�8�=a?��xdS�H|;�y>��<:(�= �ོ�-���rp����L������ǽ by�{-���so�Y�+��$5>�{��_�μo|>=8w=<��=�	=�N�<Z'9= Z�Y��;f�(=��>nΏ;��e�x�N=C�#=�>'����:� ;����@d<׎���νZ�W=��,�`N�;m��=ʁ;<��=۹<=.K�=�7�<��̻��������<����}��^e���1�=<�*���[�N����	�=�ք<Ce��(ݽ�S=o������"��Cv�=H;���\=��=�V�;UFr=5J$<y_�q�x=Q�8`���>�G�����񹵽�|<��<�w<hVA=w"�=�뫽�I�=� _=qs�<����sy�(��#���I�N���U�)Լ�y�=˝�=u�Ͻ,�w�*܂<M���[���Z�d/½T=�lѽ(���RYǽ�O�==Y���+:��?';�����=ˉ�=������=zd=��Q=!��=ƒ�=�OJ=�►(�O�Xt�Lf�>���+)�r{��Ef�'F�=�j0�� ��~n�Ta�B��B�M=�?̽���2�;��=�!>z��<��:�>t^����I=�]�=~�>@����=_D�����o�w����<�:�=�{=���u���t�`<���<t]=l�%�����ʝ�=�:�;�S˽���i�=*F
�]��=@(q��\Y�]û��)W�n����i�A�X���>I!]��ɠ<�t;�r	o= ( =�U��I�=����=�T=�=� 8<$�ҽ���R紼�7M=D>�A�� ���ͦ<aB���s�s���j>�/=��>�#��̔��sj;�/a�J�ab#�B�>�k^�5��<�������;{�<	��=&�O����;RIʼOy�=u�<�D�����'�;/_l=�旽
O�=fԅ�Km��5��=�.U=R����R=�f�=�)�=�)����=���=��4=Q�$�cU�;^�>�ޭ��e�=�D�:'2�����<�,뼪B��TR�=�;�=��=M�=���^�=C^�:���<��];S��>�>=�~@=���QQ�W��H�K;H2��u��-�����J��<�~�<��;�n�=1�軫��=�Z="�9>�M<(^Լ�`�����+U=�l�M����c�<����g�=����D=^��=ݗ�=�N �j�e<�۽ǟ=	↼�XҼ*��&����<���=~�=�Q�E���D?� ��<���^���,�=!��<��#�i�">>�+=�t���Z�?#�=i�(�s�v�a5}�����f =��+=�Dr������=�*���3̜�bg>��;�=!?>躺}��;��	��6�U�ٽ.5ϼj_+�#F��۴.�T߰=}�T�����R�f��=�e%<�S�����)�g=��<��-����)�:�=S�[;�8b����>�ѻx��=�K@<�bE=�Ab=��N=AŽ��=�������҉=)�3��B�x꫽Bc�=���=S���[��U�=���>N�>a¬=A��=���>���=�4����=	o<Z|M�z�����>�o��m���lu��y�Ib�=��7	�=a� >2�@=�p<)IX<v;��}�蒽2`�=%/�=.�U=�KƼ+�<>:p�����K�a�!��<���=&�=�@Q�z@k�-��]���E����H=J>�$�k>�����"�#f1<\�����n��}�y=KХ=�P�x���w�;�_�=ʒ=���Vϴ���)�9�=A��ǿ(�k<ټ,���jQ_=�n�=��j=+�">�Տ=�z��p�6����;+^�=K�˽&�'�z�ý�X>�H:;�����&�������=^�e���0�\��;#e��_�=��,��_��S��6ܽ?�c<���<��=5z�;���=�ט�Y��=���"���>f�v�����ށ;�� =�[���q$���k&�hq�=���t�v=�hg=53���<B䳽��&R�����=�ɺ6٨= �����-g=?�.<�8���B=�3H��<=h1�=�:f=�R�=�ю:k���蠽D���Q������`�=Q2M�5zK<Q���/�l#����Խ���=WK�<��*=���כ��ʹ[�Ex�׍:=-'@<Y@#�3�w=���<�̢��:L����=)_��+���~��Vo�9Ⲟ;�X;���P=��+>��"��&R��%9��\����I=A��=�X������2=��Z�{Ƚ<����L��;nj�<$�W�}�L=���<���؇b�k����ZM�����_g���>�m��Z=25������~.��f�<_c%�+Wj�u�0��Ý�7R����J���+D����<�X'���C�Tu
:L�><�*�:�'>zQ�=��Ž�3��MѼB�=��Ͻ�l�t� =C�l����=�����=j�=�|�=�-Q�̍�;7��/A�=����L4�=p1�=�,<F����O�2��!�w���C�8�j�
�=*唼V����=ep=���=��������a��;��C=���;ˮ�<������O=>��:�=��=�̚=�{=�e�<�3>Gb���%=�fؽ�=���٨�� =�Lh=Q����Q��LQD<�;�;Q?��	/�C�g{<�qJ=���=/�>��=g 0��Q1��8�1W��G�	����&A<��r���6=�;`���t#��ㅽ(���dT�=��+��\ :P��lʆ=F����=�)�<��<��н+D�=��!�/d��f�= mD��%�Ru>v�O�����-2>|�
��$=6Z�=����		M<�	�p橽o�"�7]=�x����=l'(>�l�R=3@)=���",�<�=9�=C�=0[�=T}<�����@�=�/�=K����?�=U�[��L>��j=�=����=	�<��<�@�=F(�<�.�?�<�u�����!��u�"��H�;��i��V���"��=wQ�WA<6|̼���=�����C
>�Sp�n�=�`��<�Gڽ�2D�=j̔����u��;�G�=b��J� �Í׽���<^t�;�Ƚ=З_=`Z6��ռ����ˢ�<I"3�:=n�J�)+F��HS�I����4��>�`нw�;���=���<�归�>�a!�7�}�=�#=�;�Ƭ)���!=���<̉!�X/�������A=��=R�ӽQ�ҽZW�=���<W7н���=.�7��p�=�>s>���G�=�K�<	����R��O�]<�R�<[�=Ӽ=7����h$��HE=(7q���-w=��ۼ���_�Ľ���=�k��n�ȼ&u���F�Ar]<����a��q�;��[=�g=�������<G�#=䘳�)��& �s���y��_�=&(>�_D�v�<��ӽ�<��=��|=��;>?�H<{��=I8-=�D�=��7�;:�څ�ɏG=T.ڼ����w�=Q8�;�M�kJf���<:�!=B[��B���+���~=��H� �=���=J��=����q�����<Ѹ���=�>eQ�=��=t�>~ m=���>݂��5?�<�=xj�=�»�l��_�C=%?��_�=�5>�5>���H����`*��>5	�=YA����+ �=ǲ=���=$�>�>Q�;��I1={��<4�u�k��?�S<�b��5B�v��=jz��x?��@;=�S�q��=,�$=N�`;�p=1�<X���_�<����<�0�=M�3�)��=�<c<�뻽�I=�hL=�Y>=�>!��<�%&>�L�=hC>!1r����;������� �=���<kh�=Y�P�����y�=v1�=O<���=k�˼�[�<O���gD�3�z�ņc>{�"�I�h��l�=k/
<�=�Q;�J�h4��������=d>�<Rb���3����_�t�v�=�]罷����o��Gl4==/!<���=,�a;h]�ٝ�=�G��C	g<X��]�����I<O[ = ���z�]=0K�0߯<$L|�q��=�c�Ï/��Ӓ=�(��b=�����)����vW�<gm��?�<�}Q<�ͽo�<�@+=1\����>eS�=>�ϼg��&�)�:�<��<ImO=�<<p=4�=s�K�]=SA��Y�-�fP�.21����=�K���b�=�3�<��J�!��=k�<��������)���r��>�����=r�=��?��s�Q<�=m�<}���:��˼�Z���]�=���=���=�$M=��<]�=rJp�qf�=L=�=��F��=8�<>����|<��́>�������=O�=4
,>���<#�;ty��>2f��v<i	�$�<��?8��SoM�bM�:p� 2]��ɖ�1���>��<-�=Y@B�ͮ�����<ur��!,�<%�<9�4�=�B<RN=�ʽb�<t�7��֟=W1[>�7��Pd����K�;C��=iͮ<�`�6D=^=[�$�o�����X=.�������Y�D���&�=���<���L��=ժn��VǼ۫�1��=���<�4>P>�C=*�A�S���s��=����M��l]=�MH�Rj�����>�sf>�0�<i��Y���ٺ��Q߽:�<!3���Xռɳ�=��S��~� ��=�l�T�j>��)��Q��p�>����m�?=[,j;��ѽ���ɵ� �;<��Q�$��=�0Q�x=&�
�����-*>ɮ=#u�;��'������=����K<]�=��A=	��<�T��)"5<����t\��`< p��~��@l���ɼ���l"��F�=ѪA�LJ;=�\�<�=�f>BG�a7�<f�=/9��Cc�<��)>�a�}q�����<��=C�*;�G5��;�<��=D�B=y�����k��Q��쏽��w�a���]�w=@�=�
{�W/���=+�<��p;��N=o�罹żf-�=��n=�b>z7��L�Q=e��q�=�^8���3=0)=�*V����={w!=_fʼ�J��'���@=������=:=��<w���L磼�ȼ�e�=&�=���=';�=�׊��=���>�=z|B��3�=6��=��0>�\ >�>�q���괽�=����y:+=
�%=ː=h�=za>��<��������
JZ�P��&���C<[*<>Q���2�=���=�s}�B*�=��H�9����;�Ό=���vJC��"���8�=�{�=F]%>�f����<��=��U:W��=
2:��+=��b� a�=�I�=�͉<��T=?G��ޣ���=�Ș=�Q���D =Å<+�>ҩ0�}3��Hfm�I��0@�=��=I_�=�x�;�T�|i�=�}=�d9�3��=Y�z�e]*;�M�=�i�����=�w=1h����=��>���=]6�='�S=��=��fv��;2#� ��=V�<[Sc�m�=$<߽����^�=�9A=��{=2>�Խԅ��\,=Ĳ콷P>=/��*ƽ��ߍ�#�;F^�=Q^��_g4>�Q3>�?�=�Z��$4>�[�=(��=�,'��9<=}����Is=�e�=�g�<3���^�?<���=m]U=�'�S���6X�s�==IS=��e=�Z���6��< \�ZZ�=�B�=⑮=�X�=�� �z�����\N��#!�=L���'[<��3<����@�
�p`L�t��;D�0�%������L�Dz����<�>��=\�J�t���4*�=,𽟹#��<��;�M�=��?�Y�A���I��ˆ=��=����&�Ľ��}��>T����:=�}Ƚ�$�J��=�=M�=(1=��=9	�a<i��<�c<ũ=z?��v=�=a����\�=F�J���u=)Y>�*>֤�={�5<�� �v�=3��;)�����</O�=k=�6}=ռ6H=�-�=�Iӽ�+�=Ѐ�=zL�<9 ==�ã�W��vL
=���=u=#=J��5B���r>��<�)k:����@M;�̇=X���v^2� �=���<���=D��Iǔ��7�<Y��<�[�=go�=lO��6�a	�S��<�&O��<ؼ=^<����=r"�'c`=g���h`����6=��0o�����=�ƈ��&�=�Z��]!J;T��={D�=J��͒<h���<�_�<(�<��j]�=/��"\�<�%<��V<��LV��|;T��=�`h��b�<�ײ���n�钼�-b>+���)�=/1A�rcȽeA�`U=P���9?`=
�D;��=�����E�=|4L�z��=b���t�S<�(�5�=�ϙ=�/p�,���؜��x;���*m=�O8��x���w<\O=��=��!��l=S��=I�����*���<�	;��* �N���P�<_�s���u���<�`-��x=?��=W��<�s�m++=.!|�QV�N�;"Ҏ>	�����ʽ�	>�P:��b>n��=Z$ǻ��&=�~o��M��� ���<��<��E�x̽�1����=>y/���G�v�i�m��=
�N�	��) ���]D���?���&�h��<c�����\=�󎽭*��m���y��^0����;�((=�1��_��=0-�<��܁���<^>6>��|�Ϲ=_&��@�&��g��nJ�=퇼X�5�m^/=\3l=�>=�� �=�_���?������w=����̱󽰭�;��̽�潸8�=��~W>̓I=���<(��]�=�zG�!��=1F�=��q=vn>��C�h�1�j��:V��h�(�Fq>9\�ؠ1��^�=�=d���>��=��w^�u_��&Ox�R<��$y��� <'䌽�<�=�b>�k<d�����=;�K��M�8��=��=��	=�,>i���dZ�=?+�����<P�I=>qk�@����e�=n�=4����=���<Z�彻�.ǚ��ۓ�ċ<���=x�b=�oD=��>�w�=���܈�=�DV<�����B2��@B=]i=�Hr=��#<bc���!漒.>�P4��"�<�X�<Ҷ<�%���������ؽc~���`=%��<ҿi�ѡP�<�r=4U��Q޼V)?=�HN��}��*?�=g�=@#��D���^�=.o4��G�o��<�!��=�!���Q=	>">�|����=˛'<޾��r�j�!�B=u	�=���o7�
ۻ�d�=W�;��=)b�=�()=�/=�?<T�=�%l�6�>�U=���<5�;������<T�*>Q��=���<3�=��T��� =v�v=�i�=�׽>�j=���K��	���7������<���^����=g���E�=�D�=c����\>z߿�]z<b�!���=H��;�\<<��	=�/��k�=��I��=ɞ�5��=3�=�ͽ�/ ��Ә���	��q4=��=� �!�ػ�W�<�����MϽ�d=9�������=��p=���=�d����@ˑ=lG>k��=��`e=f$�=��ٽ$\��\u=�)K��;�m�o���l�=�4��=���t��׬n�o�<)�y<�;��m
�<l�ܽel޽׏�8x>���<�yG���=(n�=�����D���<ߍ�=V�<��
���s�(�5��*�=���hw0=[[I=�����W3��'�=�����]ҼU��=J/p���[=���<�4�=}���?�=���z�[o�=Ա2=�,>��ü��=?+>�#>�0�=�N�.6�;ޓ�U�>׺���J~��I��V�^=E��8Q<=�-><��F=v9�;�c�;~\�=����= q/=;�u���9�L�>��:=S}&>��F>��=sE�<t�q��_��uw�=ۭ@<�YF=��\=Ž6軺׉=��q;������<G���Ȉ������=�V7<�3K=y±�)��=:����$=�<��,x>���=w��=K��=������Í��5��$�=��j=QH�=��Y=g)�<d�=q�u�U��;{G½cz =�V=�[��� -� ���=n�4�� �=����jH>?���-�=�aʻp�%<�*>-=����Tj��6�F~��3.;c�c<� �94��An�s�?�O|>�j���x/���ɽ�q�F��~��� ���m��=�D�>��$o�=6%<SP&�$���&�=�����I�=Ю��t都)��=�ú<�=�K>>a3��Û����=KO�2�s=<�t=6,����=jc���z�=���@[=f�޼��ۻ>�[<��>��=@�s��
����Ӽ n���<>.�˽�==H�%<�p=_S��p�A�����ѝ����������2l���R=^�=4�=n�I�����QBi;6����x=��=dW�=+�?>��,=k�<�o�=��=L���AU�kc?�L�=�Y�B��=��I�;<1��X�#�z�g��=�V������=)�>���=��½"��=^
���R���>�'=��=�"Q��k_<�W<�hg��]սA�=7�=�ν��9n>G=��(���5=�s�=}>�j�<!t*�wF�
f>���<�ؤ���Z���=ڗ�=GH�f���^%�ۅ�=n�����T<���=c���CmJ����TP�`p�=�ɽ�@�=C��ڈ��o�ɽ���=���<V�=��>�
��(�\� �>�.=~X˽`Q=8�%>�=�[ʽX��=��"�4�"�D� <���=g�=E�C�dT������]��mA>�*޽��>=�<@���%(�ڌ��A�@���>=e
����̎�¿c>��=�,�=��E��SQ�T6=U(�3Ν���Q=�ǻ���<3��=�V�<:\Ǽ�+��<��-���Gt�=�����Û=��S<j<���I�=c��#���Ҿ�="���y��]�;���� �=�ѻ=o.���'��{�<\f=~=[0�<���<��o�#�C���[�d��� ,.���9<��=u�+<�=�ɴ���=;ˋ�*�	>�J�=�+�=S�=��=t>�νI����%U>�a :_��=�
5<H��=2�*>��<O�<�￼�Q�<G$�G�A=�\;��;�ͻ����L��>� ߍ���?���2�;	�>�;<�_���q�=���8�R��v�����3۽�O�m����0=�����=��Q<�-��?m��պ;�A�=��=���譄=�����5��P�">Z�=m�;�Z��ٽM�>QE�)>�9=40'��!>E ��񍼏#G=�.��`=Y���6���j=���=`";b��5�(��4�����#�<�6ּq<+M<B�=<�?�=��<�(��m��G��p0+<IK��[Z=�j��xW<1aȽq����J��2�=�:<,y�<R��<Z+ѽ���.L��q<俑<��=F-9=�4��W+�=��Z����<j�=�S��*!=�z����>�4߻�
;���<�S�;n޽��ѽ|	]=�ٽ�7w<�ݽ�T����6���<c�=%�o��+»M�R��ۼk�=�����a����Ql*=҉��v/�f�=ܛ�=�Yȼ���=↢=��z=g.'��Y �>��+��=.@�= Q�=(�=R!�<��<������;!�=H�"=�f�=�j�<�!�=���=k��,�=:��`~<Bb߻�>Hn=�=�c=�'u��v��_���<��8�'Є�K_D���=9��z㋾�����0=���;=�<�wg=a��=fR�.
r��T�/��=2���) ����H>)�{��>���<nɔ����{v��-��=��=y1��ZQ����=s�+��\
�Ah=_4=�)�;�/>h�,���ݽț�<n�Ҽ@�=>�V=f�=�ν�k�=@�^=łX�%gy=�e۽��=����<B%��t��=_����=`��1;'���=�Ӄ�K�
>�~���桽߫�bv�OT@�z�*�b7>kƭ:��z�8�<��=�۟<a8]=֢߽:=��9= \̽�y<柽i\�<�'�=�`�~1�<
��i�=�=n	�4�7�G<=�AL=��=1��<�V=qŒ=*��<W����f�;;U�<[�߽>s�̽꼵�J�\�<���=`=U�?=_�P>h&:�A�ePA=�|v��b=�
=�9�=�>A���qV�o��=��N=�o�<�$���+ټv�@��3a�PTc=�c����;k8=M�b=w�����=��ս��>k҆;ȟ�=Ӡ�����<~����:��!=�ߍ=B1�;�3�<�V��&.N=gk���=�(��Gq�<��.��N�Kd�<-�{;5;��V7=��<J�g=�:3>��1��4�<9��3$�=v���u4<ĵ�<�r��4J=�s�&>��G��p�<sFF='C２U��W*=���=�cB����;{#w��.�<��Ǽ͢�=���=�@<�h=���=.����0�#Gû�S@���=)D�<� <i=�.�=����"��=:�
>��=�\>r���6�<�8�=62�~۪=���<3�1=�xG��L[���|���=^{���u2�ٻ�=���=5]���U��,�<���=޽9O<��>}w�=��Ƽ�D�=��K�ǖ�=$Ġ�1v���+�<_�Q���=}4�<zy�=�5��:��9�;��=���;q���}5Z���l��}�ҫC��M��{5���\.���G��:�<���=���q�=�d���q��o
>��4=�AW=�!�=}���>�"K�}���𙽶��q�=��	>�L�?f��]�;��=g���-1=C+�=)�
��9�=2.�������=Xx=��g;W�C=�̢����Z	�p4E= +�=�C��q�'��>G� =��;PE-=%�<��R�=
���0F�j�=�K�<n��=�w��Ly�����Vk>��V;���;����M�=�+���X=S�a=6�ûk��*=mp�z�����=�p�=�p�=	��=�ʻ�#�h���7��Z��X�=Se3��wս�J� ��=��,=/Z<���=L3r�Wd�<
�=�i�=p�=��Q�����,=���<�M<f�=�����ݼ��<vjS=��=�5��y��=�I=9�<��<���=��=!bu�� �=f�(��ɯ=���=^���7��<=��ʼ_\��n��#�S��Z�L�f��0⼞���,>��B<!:\���O�k�2=�B�=�U��j�����<Q�L) =N���(�f<��=̿�=¬B�B9�;<-�=&hl=r�[� %�=�6�����<�y���ɝ�� v�:&i<h� >gK߼�7��:��#�X���������w����J��=�7	>�c�< >s�ϻφ<N�4=p[����5�-$`=��*®��A���=P��=G>L	�+#	=�]�#=v=�9�=خ��D��Sg$��m�=s_�=���=�V�=��=@Dd=��<��'ͽ�WH�$�&��4q=c��q�Z��1n>�h�l\�=��=9�>%ֽi���}>��Y=I���"�[=��=:Q���?=N�r��]��"�<�ױ������j��#��=�>U�:�M�>�뻼�n��#7���on�s>�X>�z� f�=%�\<a:=���0�:>� �=�?<���=֚X����=6ݽ��G��h>��;Z��<@\���
>O�)=�P >%3�==N�>��4_��6��T���a�=-5> X=�&�P�67��;�j���<�ϥ�h �<�|=�)>a
<��=q�<Rڷ���*�T8�=O#�=I��==9�==�=�d=��>����$k=+aj��=�=����
�=q:��u3d�b�=M����έ/�����8O�(=�O�j�s�,r��w����>J��=�úᆚ=c�<����&�����=Y����ּO�=�% >�x�q3�=i�<��B=���5>>��_���;#���$����l�#�=���;����Q��������=>O�g��=���<M�6=��~�j���+_2=�"��H>(d���
��꛼�yX���>�,��|�<f���<1<��-�/ܣ�	��=wc��ȼS���H�=��	��	=K%��p �=#�k�����Y��<����E���7$>_���O#����K�>�fټܽjM��!�=r߼|�Ž��+�>w=�=8i����˽��1�4�>𧗽�g���1t���>���=�Q����]=��	��4c��c�5�>o��=Z�=W\	�N�<��D;�2ڻ��<
�k�Խ��_�kz<K8>O� >+F�;7�
<.��;�I?�WM�2=;[:;��Bg��&X�ETܽ�������
RY>90F������,>��C���=��a<vWz=S>hx���>0OT=x��=L���n隽}*[���M����;�2��ĵ�<��x���[=�L�=�J?=���=�:L�HE�=��=���ٲ�;�.�^�w@w;���6R��i=�0*�~�>I>w�%N�=�Xl�ib>%��=1b=�>��.���5�<�qK<�0>_��=-D���>�������f�񼧱���<=�8�=�>�Ֆ��n��������=
]��_摽�o�=��%�ݼ�!< ���;�;��]=��=��=������<�=_��H�=Q�(<�=�,Ǽ\>#W9	Z3��Io<.��J|�=&�<>��<�\=��M<#w�=�v���ܽ�� ���$��<���[�=�>�a�=����t�;��=�IN����=ٻA=l�E����#��=�7M�oS�=��Ž���;=��<��<�P�q�k>���;|�<���=IW�<^�:��=3P��A=�˳=ۘ�4_3>_�A=ۯ�=�dֽ�S�� ��O9�e��`�=j�f=�t&���c=8�<�'t=��!��M=�施��>�4�[���\W�<���둢��;�=,{(>,�1=��C�������Ls�P�y=�⑽+=ۼ�Y׼���Zh�����>H�ͽ���=n]ǽ��<�3��U=y��<Ji�ϒ�nc}�J��� 4�=ٶ=���܅Y=*�=�����9���=���Ȧk=�f<+���AM�f'��A�;7B��l�=���<�^�z�� �=�؄<�M1��0=�.�=I�>K�o�K���my�=G6_�v��:�d�I?�=�D<���]uY�ı��U��"�1�=r��=��2=v��Y�<n��5/<�������yp������'t=�B�=CBj> ��=�1b=��D;\@g>���=,�/�ܔ��Ԙ���Jq�� T=��|�Y��֍�=�ǽ����s�<Э�=_���0]���|�Ϛ�gD��������=3�&�˽n���Ü=�$_�ND>��r���;>>�=.�(��F>���=�g>��Ͻ2����$�;����w��=R�=���=��<rA�����!^�T�
=���=��C=�P�=�<B��	>���9[:�#)<ڈ�<J{�=��Ƚ�zĽ�j<�'Z���������<��C=h�&��>�l�<M�	���<�V��=&�0�����u�>������:싽Z=��b=�e��.7=�6c=��6�'>7��<�0:����=��2�1�:<oGb<41���|q�%)y�� �=�߫�aiʽ���
=�>�=�������=Q��=���=}�?� �;�1׽\�ؼ*��=���=i���`�<x�)�56��{�;=���Ã"��lԽ��=�w">�=2==���<���޾�<0�=��m#n:�{�$e�b�>fhn=��ʻtO�`�;�{ܽރ�<�%>� �����jJ׽��>vq����[=��s��nG=%�D���m=09��2��,�5���.�תf�T�8=��(���=۱=����A��!�>�R,>�A���*>�)%<N�@�ZX=Fx��7!r<
��<,�*�T�ҽǼ��]�=1�=$G-=�=��D�ͽ�AE>==3�>J.��AF=�==�W�� &���=b��L�=d;x;a�=�׋=��нU'�<�c>��l��:��;��=M!���y=����(׽}��=����u�=wV<NN[�$�p��t����l�<���>n.=�#�=��=��9˘<�,�,n�=@�i=�l�<[f��U�� _��V�=�_�<�
;G7$=,R;YC�������=\����ڶ�=��P=���L7w=N����31��˲��Q�7B���=�]=:��=��M���	P���D?=�:��F��ɠ�G0���M��E��u:��R	�=-�Ž1c���\B��Z轋4=5�Ͻu}}��P�;�N��8^=�$��d߻�����~_>����9� I�%c�=�6�=��=��k��D)>��=�N��U�<�b�+#
�{@[;��<ٳ=w�����������d�+�K=R��<����_�=��N>'2��l>��b=<6�b�%��=T�==�����eB�C�K>MZ-�����=�&>�u
��s_=tp�<Ͻq��Go���8����!�<��;����<!����NsT=���=�n�<ձܽ�v��"f�!đ>:
�=���������<I�=o��魪�;r>�����=;$0>�1��m�=ъ�=���^�=r��~i��y��0Ӂ<>�>��=�8�I	�� >|U��x��<S���*��<����4$��wi=�w==/J�P(���>� f���<+����~���(=�{Y=�}T=2߽=cZ={'F�>���K�=���=��=�ا�=�ʼzbM=�z��kJ=��S=��k<�(=A����È<��:=�\]�p� >�+�������;V=a-v;Aô=���=�D=��T~%=�ţ=���b;Lݽ{�������?D�=���<f�l=�wF=��� ��=+ww��օ=�E�x�ļ�o��C�ýYx�U�&��� �T�������Z�:W{b=��$����=�x;�5�<��=���<MNݽ0]��mx��,�� �>&TѼo���|w��vͽ�̈́=�w=�K�	�;���p�@�8�]�D6,=ۧ��gм�=�%�=�� >��/<�u	��N<_���8V;�N[��-�=�=w��=ƺ�=B͒�-i?=Fm=J��;�(
=���=���3�H=��Z>�w���	�c6(=Y6���x��ue0=u�/=\ý�%=��D����F=��u������=O����[�n�Ž���;�P">1�A<�|>(z	=�$Q�ĔŽ�<5Г=�'�D�����3�=�j�=&1!>y��=f��<]�w�2w�=A�Խ=hZ�A��=3~���ə:�I;=c�A�q�=;����s= �R�ĸ��y �� ֽ�d�=-=�ɳ=cH�]�I;�����<�=�=�hؽ�c�����<	�D=ܷ���=G�н��<��ͽ�]ͽj�=�N���
����<ص�#���3=��/F�=|n*<㛵�D�&��>1#�;f�=Nz��g���.��=�,�<t"�{�e=g��<wu�O�X�{�X=wS�>��<=؛��|_;�x���Z��P&��T]<�R<���=���Ց�樦=P����@�<��ʼy�o���g}���ù�S������>�u�j��;<2?�e�սW�=�\������}׻˃�=Csm=
x�=�^�<
�<��� ,�,L�=|J�=8)�=�Ľ�=��V�K-�q�u<ٸże%�=t0=�1��X�ܼU�p�fr����<�5�,󬽯χ=d���8��=�)�'d����)=[0���"����<)}��ٛ齋����=�w����=I�d>N0�=N�罠V���=�b��?�=;��b!<�瀼@!'=[;`���=�K��=��>���fZ(��j���r=��=������Ǩ�&��=��=�0��/
��du<[�=��������]ƽ~p�<��=�\��A(=o�<���*����c��A	�֏��]�y���۽<����/���W.=��=�u0=|��<��,9b��aꤽ��u>9�=LU<<�p=k8������M½F��=X"$��!q=��<��B=xv�=����L��C��w�؍�=�i���M�%�պ���=�9u��=�qʽ}�˽)/�<������8�T=�O��:Қ�;�%>����^�;<��H��[����@�V=P��*��=ET)=2�=<4>9�=��Ƚ���=����h|��*��]�x<��>�3��5�U�\�=y�]�XQ!=���Ԭ{<��D7j����}&�%�h=�P=�"���~%>&m=�੽C��f8��4�;��3>�뱼�7l�#�>H�<������<J?�=CI���
=_K4<l�1�=�[D>:��������<>�*���#��q��3�G<�5t��ö<'�u<]��=Rp������-Ѽ�1<��=S{<�_i��ʽm=��$��<����<fi����b'��]s=��;���3����1=�Ë�5?l��x����=�&�Ӱ>��=�۽���=g9�=��=6��=��9=��<|��/�=�7��e.�=�X>�B���}=v
��+��;�)��iX ��T��X��m��=���=F'�=��-�:S��7<Yy��x�O<��=p�B�Q+=�r&=�H�;��6��(���O���=S�<qM�<��Լ����.�<�ak��Jg=V̆��<O=5��<�6սEj��i�i�q�����=��<r5��k�<xD��}��7��=uB��ig�=_�^=9E = ��= �ֽ	=���ݣ+��hD=�XN>��`9���t釽>g���<��ɼқ�<MuH;|0�=-�ܽ{�Y=+y><O�=+O��v��ZM��Zy=0�H<���<��:=�P=�5�<,���S�/�Ka�=�*�`�Z<��p=M�}���H=�`=@���gv�����pf��E�4�g<=t�����Ϯ=T�a=�N�<p�,=���$^�C�c<����u]����F�@ýU���J��=�"��ɯ=D"�~�I=�G��`�W����<c�j=<�=�z->4�M�I�x���h�������н��!>#�=�ݫ=)j���=�(=�u/>B�f����=S�1�&u�=.����	�=���<>a=�?ؽٛ�=V8��D/=¼ >3�޽-S� �H>�6�=��e�%C�<�>+���/'�=�/>�	G�:�5l=<�=x�<�.���
��*����=8�>���:[�2=�W�:�ֽD>��@=��;U׿�ӳ�������(�t
�=pO��^[=�s=R�ʼ#.����>��>��뽠��=�<�b={����L=�P�;z{�ws����	���x���= D�<���=B����)�z=������T�΃��X�{=���=��潐�����t���=�/��	��t���5�<-��=���;�"8=�H4���<�<��q~�D8>E�>
?���>�9=�\ĽL����`�4�M>������@��'=;����=�	$��Ǽ��>
�=�D��R|X=̓ԼC���(|ɽ!8���U�Dm'��U��������k��@R��o���=�`��}��O<�<�|���=5J�=��=N� ���>7͘�2>T_<������=e!����)<���=��K��g���> ;�=�i�=���{Db�����N{��9>*�9=I?���>0q�=�C���>�m�9����Y=GXټ��=5��=x3��Vf�ٷ�9C=��D��Ȱ<tW��휋<� �<%!���*Y��O�<l-}�@�a=鬁<)8#��ǖ�;u<���=j�n��c���-�W�9��`�=�I���������J�<c=>��)����N�Ϣd=d	%���w=;� =�$F=t0�<vӾ�[:
{�<+�<*�U�K�(=�$��ǹ=RN����B=��D�Vyj<�8��r���%��8z{�=��;,�<��=�O�=��:<bʼ�D1�>�s�&�=��w��b@�c�%>�G��f9�=w<�5�;ç\�}b�<|���<o<		����<�5��!�=&e�8��:>#�׽�r<ʉ< ��<��=u��<���;7� >Tъ��������4j���K齈�H��缱~�=���Q�8=ڮ�=9�<9f=�콃%�=�S<唠;��ѽt��V��
Pe=�!>��v�\�L�-��\B�=.��=�
�=�(j�X7�l�#�
���k�|�#��3�i��=�y��K�m���6NC��Y@��4����=�8��x�����<*-�=�&�=���=�W<�t=�<Y;X꼝m�=D�G������i��L�=Τ�;�tT��V>s>���=}y<=��=Wi6=���pn�iyҼ{���?�<^=�=@���-����D=�D�=A3G<������;e�K>�ӫ<N,�g2w=�ɩ�h�ż�;�=��U=_�C�g���j="��=�J�<l_��B�7�}���T;�|q����=�1E>�x�=��vX���fK<fzi=���0.G>l�轖jt>`<��u���V�˕�<.tW�����ǂ��,;�+ƽ#d8��>>p<�:�G�<�{���+�<>7;�c�<�"�9=�F�>�>�2��`㐼�.r���������~��T�=�g�<0�Ƽ����I��=���=ּ�5��ی�=�:*=���T�X����A����= �U�FcW�՝�=i��<G�x=�P��@�=b�b=�b�<t2<�(�<2�=��T��r`�ؑ����*����-��K`��_�=9�9��;���<��9K��=V�=��꽱	c�Et >���=��<I]�=\�N�L��7�½�/k���Y<�P'�t���<�"~=
K%=)�=R���v��o�����1>ͩ��]4��,>Ҫm=�י=���=���9g��(W�=;l�=��x���u=#�?<�r��M�ƣ <�w�=#��Q�=�㽜f>%�!�i��=��Cf����O=F�������-!���=S�]��\�=�w�p�,=�U�=�:ٽc�$��~1=��>�L=�a/�<�I�=8A<��
>�G<`r�=��=�����=�2=1�=罿��C��==������;&�Ƽ���=`be���v=�k�=��� �>���=�G�=��T;b���g:�=.H��">��<8�a>�5\=)�=#�)=�I��a�=C�t�b�j=8]�=���P�A�V���"��o��3�'�i�����=0�"<zE�<�?����=3�k=nR˽!yK�B^���_�P���[;������*<�*�;�S�<��~>w�<�\��jKʽ� ����<�PN�t��~�;���ޛa;�:�<됼�]D<mԿ={{.>6��+�s=�<=f{�=��=�y��>ș�5�w=?��j�%a2�$])>���q� >�'Q���0���m>�l>������;��=�3>dS-��O>�����=-a�=$���g��=﯃���?��Ľm�<%��=ɦD�Pq�=���=�y=϶(< ��-��� >;�ɼMӷ=��5=ø�=�RY>��<	��=T������)=I��=P!/>�$�=#@A�&=��u<b=k���-��XK��÷����3�=Qk�����
�"=d���b��=t�=�ā��X=���=w7�'A�I�s�����"�<c����<��;�9#��5��F�<��==��ܼ���=
eG=�}%�`����;>{j<j׽��<��޽�ο<Ŵ�=.���X�I�>3�<�ܪ�U���q}�=��<6�=(�=gƝ=��6��D��n������;Z=|m�䣖=�j�������r<��<8?�<CB�=ˋ�=�B��j�=4��<�*z�p����I�0��=T\����=����]#��}����<4,���!5�������B=�|�쳕�v���^Z�֞>�f<�S!�G�����������=�?�_��=F��=�SZ�W7)=4�=@:��O���t���V���p�����=��0��=��U=#(��԰=����x�;җ�=u�%<8�˽�B�=�.;vc������/4�=jֻ\�8O)=����"�>�=�M�1?��1<��9;���=�~2=��~=�Ǵ<�>�<�Q��=�S���$�<��� �,����=�芽�B�=��w��%<����T�=,}�=�3=UF�=���=a�|;P�i=��=HN���K<��#>��)��Y"����=�C�<i��=���b�K?@����Su=�v�=*������]=���=9n���e�=���<��&=a�W1T=2)�<�E���=��� ��c%�=��0��*�=g��VE�=:]/=����� �FE<���*��<I��z'����;�x'��g�����I�֎e��b=R(g��yP=���=`�<=�=� ND<��Ի�#��	��./>�� �05�9��D<l��0�=[b
>�b���<c�8V�=�^��|���[�<t�Z����^$E=�pq����=�=��>�6���T�=�nz����=��=q�>�=8�=�]��Z`���N��d�c<"��9b��FS*���=�B=�b�=�;���R�=7V���-��ё	>��=0�$�w��Z1;���=��<�Zѽ4��#��=keI�]<�<��G�u�ޛ�=��J=`��=剀�G�e=��=
��;�ѻ:�=�,�<�+���^�<��&>kv1=�;�}G���@=�������-�4�8����b�"���io��&�$�J�;���==Q��<�����̳=����XU�=�S��;�	�A�I=7��:$���tF<�0׽�=�y�=�M����=N����<�B���ȼ��L<ͣҽ�6=��o�D;�(	�=ne�Ek]�A��:w��=�<k=k�J=�H�=�]�='0V:9���\*��EM	���=d��=�UY=�6{=ƿd��В;Y
-� ��<+�z=�;K�2��<� �<���<H���>kr��y�<례<���J�#>��ѽV฽�;�Y��۽�c�=v�=�|�<�襽�½?��<���=�R�=�^�=������=y��b~>�#�=�Et�*	:�[{�=3���1->����>�=]E�=.G]=!W=�͍=��ཁ����$w�T�=��ڽl�м�a9�R��=�)d=\ݠ��=6��zF�<��5�lw����d5�=o��9٬��t(>�05�g�Ǽ���<�\<p企~�;����u���=���;2�=�>���=n�ݽ����婤>Z
��#>�4�)�=�@������)��ڼ���$>�n���]ҽ��E|�=����=L�Z�ڸ#����<n�R=f>4<�(]9..�<��f6�;���O���8�>��=`��=]X:윯�>{ʽ~�;z��=!�"���=�W�=`<]�M��<�|������lr��t(>ou�=^N�=��=(�9=ƾ���g��G�=��=�Z=��V>T��_̽d��z���c=w�==�� ��:���:F�/��>^n=��R�(^W��*=j;��##�򞽭B�=ƠQ����o0�=K��dk��n�����$�-��ӏ�w*�<�	�;�z�PPH�Bi�RMI��؀=[�3='�>�������@ߪ=7���+<V��<
R�=3	�;�1�9�Њ=��x=��<�=h�/>;�2=��Q;�=�'c=�v=�#�;oc���<�_��@�<�N�=^�E=&Ͻ���<�>}<mY����#'�=V��=�c�tS^���.��yD�9�/=D�� �=m��<��*�=K� ���F=0X>�r��	�k>¦��l=bZ�;#'׼d�<��{z�;C�T��*����<;[i��&���q�X��/P=�e��$���EȻN�3�s��n���W4>J�Z��0$>��i�m�@�������oĻ��:KTѼ���=���=�q�=�6'�j�]�Vr�&>}<R�$=�*{=��=K��;Q����	=�t<����T�=�����%�sK��+�=3-żI*�<1�C�0�<�f�=��>=΢>�L<D�!�Z�<ք��HJ�={�."���'w�(=��xfн�V�<
}�<`�=�<��۽��,�)�s�i~F=���#���.�=��>*�C����=�Ml=[^�����gǹ<h�=��I=�(��ڌ9;�p=��i�r�=����c'>љ��"'"=/$<݊��Jz���G�=8�X��`	==ޏ�S7�<IX0>h�ӽ۪>yE=޶�=�f<=�>�\�^�:Uൽ�c����=R��=�׾��T���.���^=w9ͽO3Y=�Žt�=����5��$?��2;Y�½���9I=ar&���>;���	Ӱ���"��"��T兾�pռ+��<y�Z�k<���1:�E<"�i=��ּ!5Ľw������<h/-=(�=��J���z�i�����e�>����V�,�=�A�<Oý}H�<v�ٽ	�<y�E��=%��=�`�=�T�=VCM<X;�=%�=��L=�ޥ�!�ռ�C=�7�<��;7�dÐ�J�"=�l�=29?�P�O�8�=�S�<l���-y�=������=���I�]���<����z�"�=�_r����� =;�Q�Z���p�=��&=r��=�)���>�B�Gڀ=
"{=�	�pu�=�����:<��,>�𽯵�S*�F�a<��*>��N>D�<�	���������=g���(l<�u�=v>�
r�=՘� �{=� ���+�5�:�����w�� <�{�g�?� >��|=�7���즽���='��4�>�t�<�>��?��A���;=L��<�����=S-=<���=OX���S7� z�<���=5������QyG�L>�}���ҭ<qB½vu�� �ý��r=-6�v�5�=�g�=�m&;���?�p;fD2�������<rVl�0>p�RZ���ܲ<?�=�y�=�20��
�=g|ٽ��Q�i��=cg=�X�;Т�=���O=U�=�*�'p,=��;I�E���6���!���ڼ��0�� ��=����x6��y��<�`�=��=�A�D��<��(=*>��">��k=��>����4����7������&$��p2���ǽc=�=���<��H�K��=�K=��L<lv1=�q�;�>�}|����=�:�=�{=̘==�yG>ppk�P(�<mu
�gI-=��=l��i������� \����<t��TJO=�ы����:�ȽI�}=$g�<{��=�J=�Dq�;����=b�t��0�=|V$;�X��M��=�N6=�(#�[�>�<�{+=|�><�0ͽ$6��:�<��=8N�����)ӽi�8<�5�=�#>/"��$g�=�:�k��=���WXD������5:f�=k) �$�==�����V5=[f>�V0>G�<v�=y�<b�?=���K�R?�=�e�={�<ʕ׼��=�3�='��P�x<�d����w�Ƚ:��=�U��"v���#=v�7> g�ΰj=_0>�9��F^=N��<�9=�|=lY��ʑ�R0��K�
�R>x�=���9��<5�'>�W�<��<=��=�B2=#L�=8��=P�|�y=5�<��d����=)��=\��=�<�;�k_<>헽�8޽rl�=���P$K�_���2��<�F޼i�f=���<T�	>����2� =��G���=׭�� !�=w�>B���I���S�����<��۽_T콖l�<��=���=�>)>�߽W*�<��<�5:���q�Dn�	��=� 2�^D�;~Oc=�;�=��|�(��={Z���4;=gN=9l�=1@�=U�!����<q]�=@`�=!*i>)LR>,���Ѽ�v>��ꉼ�ɞ��1��F=��C���<�N�=�=P+�SK�<$PY��fW>ߊD�wǓ<,Ɛ=*ҫ=�>�<[c=	��2���}=�X�ʒνb5�=J��<�YJ=4�<��Q<�w�; �/<RG��{��6��=���<Mn�3Qb=���&�<3}>�c̼�l�`�=Hks=u�=c2���`=���=Mx��#:>��综3�<~���W"���p��7འWZ=r3��nB=&�i��ș���;�9 �}��=�a��ݘ�=��ռϧ.�Q���=]1<�fռN�3�NV><>��5�=���=��ļn��=��f��b>?뤽U���#���^F>%ב���=N>"�~�!>XT�齸:��=s]�= l���=�r�<F}��4��m>����������SW�=��=��<�Kٽk������=u[����>�-�=E�=j�>RS�<�>���=ԕ�<� V��4t=�m�<vRD��==��=�\�=��	>@P��wf�?o<�B���a�a���^����/��{^���d=��P�>�����o���=?��V�;���<�`<����Z~���>������; ��":���Ih>]!=C�=v8 >z|ߺ���\�=�ȑ��@e�E�ƽ���s������[�;�@>gx�=)����V<4�=[}��`��]�3<���\�������8�<"]�Ld����=�":� �r;y��E��.��ǲ�t<-?>/~��Y�%�,��<�s<W/�<�Z�=+o�<�n�;Ծ�=����ǚy����;ݏĽ�z�=n�<|�I��.�=me<�g7�=E�<���=$wN���=�ս��=Ĳl�#fh=�,J�s�M>Od���w�^-�=6��ʧ�����1�=��ǽ��\��ܵ��%�Ҝ�=ax��2f���(=��N���='b=JL�=Q�ͼ��%����d�������"�jǩ=m��=[���q�����8��=���nP����o=./��mg!<bG(�r�]�+>²I>��;�����>���B�<j5ؼw��=��$��f�=bS���Ļ<ݢz�y;=�=�B�����k�|<0�<��-�n< =#m>�]e�=��>��b<��=��=��<K�9=�J�=Ӣͼ���v=
�ͽ�T	=8G�=�qi�	=-s�30Խ����J���������=���6X=@�x=H>=����n���=�Q�=�=C�
>Uֽ��>G S�d:̼N��yB=,ӗ���H{x=�L������j�=���F$�<C�o=aB=t>�=
��<[t��ٽ:�����;�g2�k�(��3�=o�o=�e�-�������O˼�o>hh�g��4�>��~=���=���XX><�ͻq��=��?>��=��@6<H<=�pt=^N�=����z��`��;��=�Wq= Q�=�ݙ=Y=�����L��K��=Dɻ�=zUE��%5<.d_=A�*�J9�<F(ѽjJ$=�>T>ۈ�;��=�i>:��=��车N¼i���=��H���2��a�=.�O���<�s=���<��N>&#�=Ve)>F��轶j�=��7>��)�j�ŽɊ���M*=�X5�G���o������=�D@�I�D=���/=:��=��=���*m=x�м�ȫ<����!��% �[>V<+=1�{<@�Խ���v��=���z<�o��;Vj�=�<Q<���C�νƦ��[�͙��C���lLL=��>�u�ة
�B9���8�Q�=$��4��"��<ӎY�F�<�|�3��kV�<�x�=��=�`���Aܼn�	;�]�=⣼Z|�=|�=d����`��S?�=�Q3�"�=��P==��=�~=�)��=�B�=�| �v7=S�=�����h=���*�=D&½�S�=��/=]�<6+�;MF<@}t�_�L=˷�=œ���ʼD�="'S=K�<��2�0>�=0�����<�� ���\����9���S�=Q�J�T�(�p�g=�*�<�M�oC�=ГӼ��Z�=d(�:�}�=X%нl�Ͻ�A�=H
�<�^�����1:ս��^뒽���:��!<*C>�GX���3<�*F�&���I��q�=��F�����a@�=�>bT�����y�l=)b�=`�=���=�(�����<��y=��Լ�����QA<��=�f��n�=�!�=y��=h�=!v:�gXF�Ne ���˽��;��~=H$��!U���=T�t���/�:&n<m�=�����=�@�=���f�B��Ȟ�T?��}�����<H����n��>��4��:��<yo<.��=�)�=
et��3���k��0����=���n<دѼ��s=��F=�P�=��>���<�^��o?�<�!���A=�:e;���=��E=�	h<�S����\=Ω>5㧽���RA=jQ<� >Rb��r6�^Z��D�p!���*<��0��̼	�����@�h�s:`۞�P�^>��>��Y��O?<��>�
>�lP���<�0�;�wy�I�������෻�K|����<H�=�/�=@N�=�g
�V��<���֚��7���>�I��n'��=?�V%>��=�䉽�U��.���B;�=���>��������?�򪽈@_��9C�X�ƽ�ꤽ{���H�<���M�B��^�=zA��`Q=%QD�DJ�<+~r�|���o��B��@���>n�<�s;�{��8d������A9=3��=Ok����=�b[�94;4�=c�I����۹d`?���>��<Y�;����_�=t-�=�*׽��u��=$=0�=�}�<�X��Z��=������=��ǽ��N>'�����?d���iq>���D"\�Y6+=3K����8=���<<�=�Vk�=>��0�/=��㙽�:=M���s޻hM]�
餽Oo=
S
�	� =8U�����<�*F��󼢸4�	!�=S��<m#�=~�[��4�<�JO�A[� r=��=ӹG>3n*�E8���m�=X��=(�b�h����C�,�>p`��L��=�bo�1��)H�<,��C<��ּ^R@��vX>	�=W������=2�=W0ʽ/I�={�=Q񹼢%�=a����,=��=��Y=��(����<��%>`�4=�ğ<-,ؼЧλ�Y�a2=9�Γ�j����=n@=�>c��4�d"j=�����`�=I�Q�Po=P �=ӽ����u.����=�4==�W<;�˼Nb=���b7�%���0>8Ȓ=e+Z������s=c��<s�=]��=��=l��9_{����>yl�=�=8�!=�ƨ�n���h�/�1�K�������@<��@��(������X(�=� �=v����;��'���饼�7D�8b�<~��<o�=<>Ӈ=ɍ�-ؾ�J�x�>�w�/�G>#4���>1��j_	>����򆽩@T��[6�=Dk=�Y<�~B=2��=7}P�S� �LZϽ�?T<�u�<M`=��=�(e=��<<,�<�t/>�j��<3?��@�=Y�{=�ƽ�T�;ٝ��FY=M�ռ��Ľn��<�������y��Z��<���=���=�r�T��=�����xλ� ƽ�|ʺ��������.�=�z�A�=S=/���V ���r=b=˽~x<=6Gۼ�tڼ��>������ ��A=|�3=�d�=��<��=��+=8ޗ=d���w=J�.�����yN�=�)��5�<r�R=��k<d%ҽo�̽���=Muh=?	,�qp���=`w��u��>��=?E7����&PM�~��<��ü8ང��`F�;P����������L�w=LH=��`��6A�=�)�<��û㾽(y�<�3>���vA=�9�<0(�<�os�f��=co�<��e���)�2=,��Y�,>�������:q�#7�:*ܻ��ݽ����؝=p� =nop=���=D��<�ս�R��G�=����w(=���:sd<���=Su��<=8�����*ͼ&p��(>=�KM��(�=��u���e���Ԥ1>��q�L�<
�:U[�=F&==�M< ��=EŌ��_B=@Jչ���<)��<'����Q�R��;>��<u'üc:�����9�ݻ��T�����n.�<��.=�^->�T�<�ͻ�����߼\���B)�������=�����"�捃�cnZ���,��4��ӝ���Խ���=~�`JL����<�&��@[����=��h��L=
�v�Mһ򧯽��=� >�E���f��#U�W��x�̼[�&=�o�SD����=��>��P=k��=��.�~�6�N.�+[�<�j�=�!�< Y�=&$��d��R�=�ȩ�\�T�W|���۽��P�ۋ��zȽ��>Fԁ�c�;�^�󺤽��u��p �xL�;��<eh��4����&<�H�=��-=���=��6����<u�c�O�S=�=`=��=m��;"��<p�=~ϲ=�wֻN�溜@��7]Ǽ�+���v/�u���
м�����;����^��{z>�.���=�	���Ki� �@��j��g��N+=!�%���=�!ƽG;-;���<�������=È=�^ٽ>��ռo>�_�l��~�ֽY��=�2�<�tb��(,�������}��<�^?��6�;���=l+лe�=�>*�<.��=���<�\�=� �<��`�jH�=�=[;b=b� ���,=-��={4s��н��Q=�M=�<=�e=5�����핓������`=�<˼��3<AH[����Y=���<U͉���U��=>��>����ʼU�߬�=Dn�յ����Х�<��E>�f=XV�a9���z< ��=n�=�X��e�ƽ��v�S����=T��é%=J�Q�0��;�+н�[
� ����<��X=�G�=Dͫ<�[�ګ{;���罙�[=D��=��I<��=&>:}��[s���>��=j��<�$�AA���z��a��׵�<ђ>�W&{�e#-���<�S��xJD��>< �<5�=���P�����$瑽�[�=�;���.W�=� ����p�S�->�$�<U"k=��鼔J�<,W�s�|=�V>/򊼂��=�-(>f�>,ɽ/��`, >$�,��wҼ��V�>{>7��:?<E����-%��*�=�$�<*�v�2+�=S��=F�뽗n��=��<E�Ľڅ�=EvQ>�b�=�h=˛u=�>�+��a
=eҽq�;���p >�>��hO>-6�F1q����<�\�=����{���6���轋�~;N9�=�T���/>�<f�E<��P=,��=��̽<�>�B+=D���V
��++��?1�x�����=��=�%�=��˽��ýN_����	=�K��dɽ+��Q�Խn���
��/1>n�1���=t�(=x=]��=Ջ�����jp=@�u;�^�=e����> 3 <E*��k=�7�e�W�`6���K>wϽ/'=��P���役�8Q�1�-=�����@۽:��=m��E�<eF;�?�������J��<"��>>C���W୽�I�<�o�=8[�=+;�<����òN��٠=�f��y�;��������$����<�/>	�=�Z�=Ze �h��=f}(>м��P�<��l�_�r=j�q;�T.�,��=�6��T��;�'�z�=c�*�CM�i7b�I��f��=��;/ýW����<Y�ຓEļ\P�q/�=�ܽ�z�9�#=DY���;>�u$:�2���<y����0�;t�߻Y���7㽞��=�t������X2o=a��<Q�g=�踽���=��=�o���L<���� T��+
<�j�;��"�oY�=��=�bj�;k�<�ڻ�s�� *<L�ӽe�=v�'<�Qļ�i:=^�}�(h<X�"=x�<P`��̲�<����������z=�U�/�<AeI�-W>qI><p?�L���j����;=l�=bi�=�l��K|��AS���(�c*�el0=��˽h�����=���<y�(� �`���P�= r5>jW޽	�H=�=����>��a��;�����=d��ē���5M=��$���p=���!��<��:IH�:��c��)�����4��x����=J���b���s<�m�=㏃<�C�=�e���Ŭ;v�=�z�Ͻ4�P=��e��p�<,1=���׼D=��x��=�<x���95��eZ���=�Z��R6�����ӓ�<䠽��D����.�< J=�=K�=;Ԑ=f����<gͤ=�� �Q��<bD�� �v=V�2=�2�=�=�� �����$>l�/�P���Y^�#=s!>����&t�<�h��w�P�_�P�w��V1<V]'>��<�	��܈<3�<�=���?��^	=��=|<���3g=�g<�%3=Q'��|�=9����j����<Xn�=�/��;�=��f=)� >��<�>�G��}=��N��=?�:=n��<�?�=g�>��{��x콴wQ=jm=�N�����&`d�>Ma��X��v-8���}<��<�>�5<e�\>�gL>�KC=�֒��=��;�w��PM�j�߻��6��+�����%϶��`�<�k ���<들<����� ����=k����|<��>_�<�ĽY=��t=��$��u=y��L�=��<z{=`�$>�U=	�񽻊d�J�R��A�����O���ޚ=��5P<��P�=��j���dx<5a�=<9q=��J=f��;;����=ax�<X��=��Ӽ��=�w=�뀽ܥ+>�d<�oT=���=��x<˓�<_嘽���9<�<�b�!>T>{#e<W7!<��T>��s�
>��j=������<Df����<6=%e�|B�O�<��v���I(=j�>���<�d�/i=(=�\����D�<�'L�5I?���=v
=Jߙ=~Ө=���=d�.=ޠD=��=�m�=G{�<$t;��a<�Dۻ��?��%���
���>��#� ��=x6�=�n���@-�y�Ƽ欄=Z�üE����=RJ�>�2��=��==t���>��W�/o�<Y���� =�F��r<�^�<�q��ꆽ�������=���=?5�=�J6�A2�=��o<*��?�D>���<Գ(=���<UC!=#�)>%ƽ�h<�$�=ɽ�?�!=�jY�	~=�+v=nUZ��^��W�=�hr��+���-�7\�4�;���(�߼�<ڼr��X��=C=�L��z�G�����=�!>^�1��	�=�]����U=(�=��ǼQ:��0�= *�;�>���DR���A����=�ʽ��{=���=\�B��:񽍲ڼ��e�=W=C=��=�� �O>���<g�7��=�5����61>?��ő�%j��/<-糽�]���{Z�}o�<$&=P�!=�m�x�����m=�\���;+���G<_�=)����ϻ �<�sw=<1�a�S>�3��~R佯>5�s��6�;�Ǽ��|��Z�=c���P���� =�>>�.���]����=˥�=�I�=8ϼ=L�q���C<"@<<�[:��r���]�<�ļ�(U�p�<XH����=�d;�Ȧ���ռ�����н��D�WڼT��=�=G�T=� >JD>>1|=��>�g�=쁼��>�>�*��=|=��;�/>$���Ă=B�Žk�|=(���и��Mo=)�=���=bf`;�)��'D|��=ڽ�qq;_�=�&=��=�1`+��A�������	���V�=��=O��=�3�t�<��x=����Ŷ���@�[}3=z<T<�ޤ�����ݏ�=UW�=�TѼ�q�<�l���>S�>�ǁ���Ǽ�ʽJ��;�)e=�ٕ<$�<��>ax�*Ž�V�<�<<��mH�=����X���	���W����������.=��i��[׼�j�<�:q�vR!<��A�+���oPV>ظ�=�]=��4<�z�=���;#����@�*=��o� �W���B<�n齳f�#�!<U!-=��0=q�w=F�<�$����<���=���<u�y��̖�V�ij>���p;>�n��G5:0��<���<��=��)=U�s=��3�1<�'=_Am�:��<�J�;2P��8T����=<�n�<�+#<�8}�/5\���:=gy�<�Bx�!���h��=y��<����->��]=��O=��;r�ֽ
Z���]=]p�=��F����=?H�<�ż:��#�gew��0��+���=I=���B>ª����r�����5=eN���.���=�_�է��=X�<VO��H5��v���n�t���=e��&g��G���`��8����=R�������_ =~����񈽟/ý��S�=w��&W~���l=2SY��|=>Ӆ���=�a�=�p�=���=땙�k���s�����=$�g>�A@��s罼��=��M=Y"�=��=�?��G:>�"ӽ�'����=��\��|c��/��=e|���<m��=ƽ^M�<�ԍ=���'1���H�J&�<���<� >��6�S����>�V���k��v�3��@>�2���a�x��<k[�=��=C]��	��>��=����C^+={����ؽ�q��E�=8���%��<���<�=fS/=|/=��E<��V��������<���=�n����w>�G=Za=���=��E��>"j�<�G<���l���h=���=2�< [�=Fp�=l����;�����<�S9=�=��B=��#�xk׽�7:�6컪〻C:V=�R���7��SA��v߼�%�$��=��ʼ�C��}�=�b=W�ƽ�me�gB_�+�n=��=�!=tT�<fV�=*c���TC���=��?�

���i����T&����V���];�<1��<-޽:�f=�zf�^#9�R뵼ͩB=Ҽ�<�� ;�ѓ��YF� ��=�K����2�nz>���/����==�3!=�6���x��pc��"/B�����e���=#^����뼞�=!�޼����<�,���f=_A�=�s��A����>z~���'=仹=�N�=BM_<�T>��B�	V��ӽ >TQ�=,;	�(=R ��\�=��=��R������=r�K�>����4I�45�>O}>D|p���=|t��o,�tϽ�n�=6�#�� �;0[r�a�꼢=�s�p��=��>�����<���I��2t߽�<G  �bI��uC]���׽�F<<���x���>~3�=�Q�=��
���j�ͷ@�,T��#s>�/<��˽�R��R�R��<n��<��=Bw<��8=F�ʽ�U�<�Y��_�&���夨�$�v=�c����E>=�m��g��;gU��&��:���9I�强�0=w�:�~Օ=�;e&�<�Ѽ\2I=d�X;݌��܌��e��W�HT�=v�]�=��<y�f<��e<�Í�;G���LQ=��R<z�=ߨ%�$h�=�U�����)*�=��2=q�=5��=QP7=S���qt㽣��=ŸܽQH=Ȳ�=G|=P�=��H<�1h<Z�,=S)��0)=R{��7P=��=���c���m�u=�2�<Q=�;#�����9�����v�Qz6=���<�`�=��6�u�E١=%}w=�۴<���<[oG=g��=�=�Di=��=6儽�0���n<Y�M=��ª�=��+�'��n�<��n�l6+>DC�;w���F��=B[�O�I�;�<�+>F�߽�獽�����Ak�B�=槚����=5�������P���<��=��/�1�3>w �=��L��w��0���=gl$>��ǽ6�=
�c���,=ꑽ�<�=�n�=&�:~��=[f�=]�ӻ��=G�=*�j���=:�X=Ø�G�4;Ho[=��4=ZhB����=B���X��<�	����*=W9�=�/<���=N���L뎽Q(�_=30=��3=��=����������@E �[.��9����C>G�P=��]=� �=αc=Y�R=�p�v��=c)�=wT�<��ܽg�{=��g�b�D=r4=����ա��%�Ӻ%;=�d
>��k�{z��Չ򽡓�=31���J��I���PQ=U�V=�e�ٻN>�<���<�9���>�J=��ٽD��<M�<�ʽV*>�|�G��=�&X����=u�����Gc�B���׼���=AoH��YF�8�<�=���\<h)!=�mm=|��=ZlĽ$�=���i[,������Z��[>F׽>�����=j}�=�>e����m��<ݛ>]��x}\���TⱽtG�=�N��n>�����\>���=�f��.�=F�1��#����'��i�;n��;��q��P��z���~>Hr$��J�=�F�����=���Z�ֽ�P�=�~�<�L�U�5�B��=;=w;�=L����<��:��>���=�3�T� ����=0#�=�w6��~=�w�:Q���w�+Yi�A�=1��<�Th��56�"R=��>�²=NL�����h�<ӥ���;{!�=Z��=
=5��m��=Ӿj=���>��:g�=���9=@�%�C����y_�Y!,<>���+�>N��=���=�ê�)Ո��^�<��$=��ս�]����n>=;���-��;n���=k��>A�<6<��7�=8�Y�j���i�����･ۮ�q��4�l���=UVŽo���Ww�;�S=�����M�<SlB=WA+�>�o=��;��/n>),����H�}4���>��M_���}<x��;֐�<q`:=�uM=���ʬ黙��x>��4��Z�7=�U�<�A�=��3�I���d�=a����JO.<$��ם�� U�<���^�Fs= �=�v0�C=�����e��w+>�>�=hŰ<:F������ȽU�;��-���=ҁ�/���Y��C�=q�q�$�;<[�'=�>�1�=����k��;�0ɽ<r�=���<ȅ��עy�tO=>^��|މ���R=�b4=�W��9�͉=��$><`#��P���b�<L=Bi��S�=�Q<�<&mƽ}�9���<#��ؘ>�y�����<X7�<�}�=�
�=e�~�k�=O�=��=�<8|<�s���)�=�8>t2��|	��E���v�2D ��x�=c��"�>��w=��5=)�= i�=��X��_���=U��=���ሀ���<h[=b�>�Z������<R�,�.Tv�Ѵ=^He=��=���<�p�p�ν񺊽�Q�=��Z�
�>�B�Xʒ<�O���)X��G>><�;���c'�=u���K+ǽ�糽K���|���=`>��9�=�k?���P=�3���|���-8�4$=�5�^Gq=�ֽ�Q�<~�3�g�~=�+>?k���H>���h�3=A!���Ϫ���>��ʽ;'��=��=��>��	���˽�y>
��=�j=����=�K;1>�%�=&�=Q��&��~��A21>�U�;f�=I��<Dĸ�
�I��o�<�ʉ��^|��,����=�Ő��ƺ,��<.��=,N��k��;�C�==��S���N�� �6���>D~�<n�=��h��=�
߽�:��	�ýݓ���l�=�؃<���=䟻=��׽�@3�����ʔ��������ܽg	�q�:���=#��=2�]=�đ=3���GD�=�L���%��� ���i�11>�I׼��x<�v���:�<s ����нv���L.�/@=|M�:��ں��.�ͼ>�Ƨ?�yl�<�ѣ;G���eN:w����<���� ��a��T�8��d�����=L���
�=fQ��� �9j��'(>��@�G��ʏ�`9����%=A��<$���}4=g��=K{ڼ���=ǉ����=�V�=2��<��=��=-�Ƚ���Sf�(3�=ӏ�kr!�D�v=�!Y>�ҧ=!��Ms�$�뽟�4���'�	]��)<ڻ�<�s��]���%��=-�=�^�=���<D`+�#�;�<�=n�==���=����#B=2�Z�Z�g����=g���o�Y6ǽ������	�)�=EО=D�=^�d=�n=j�?<|�Ӽ>�6���Q�m��=���=���fn�=E������=�b��mJ�=մ=EZ�=�\i=MHϽ����^�&?�j�Z=SѾ��>nbϽ'�="ὖZ�;��н|�мHT½t����`E=�/��,�>�X��E��#9���O>qګ�$���Qv ����;�W��qB���"���E>TN6;�����D3=��`�6=�G�<�9���o�<��>>�\�=�v��wq=�@=�ę=�ZV=��~��i��)�>�+3:#M�;t8� E���ͽz7"��r"=��B���k��=w�k=��<�ǽ��V���_���<^�
<�^�0�=�6�P��=h+�~}�=s�=l�y=y#=R�v=�"���m�W�m� ���p'=>"��<�݋����:2�=;>�;>}��=������=u&ݼ�X<�2� =�,�=yj%�z2M=�(��� =�E�=R˫=��=G9d��B�=N����=�%	<c�u�K�ٽ\m=kI�<ga>4��=�J<�Q����.�(���>���=�,���=��E=��E���̼F*�=5�b;��'�Y�V;-��s�>'"�<�=��@87��=� ;Ѿ=�l2� ��*�4>��#>��̼����<=F��[�f::��#]�=R^���`<Q��<�>q;��=9VM<�=6�e==�Mqٽw��=�rf���<��=� ����;�ʘ	�������4=�~�Xߝ��<�	=ݡ7����}�7=���=b�X=p�����<iK;1�*�g����F�=y�-=��Y�Kq����<c�=rO�<Bk�9:�M�	<�FO=Ν�=����;��>���=�M�:5���V0�<���=��8=�ym��^>��=�|�����#=���=�rV;f�s�I��=HE�=6�}��b��η�*b���n�BՃ��������;���<��>1Yp=L*�=G	�<��5>٢����[��4=�л�n;>>��=�p
�S��=%����y�#��=�=?��=�!��<��E=����D��sf|��v=q��x���6�����H�o�+<�����V=���UK�=I
�=�ʼ�����V�lz�<X�<�[�xp���'�=�NJ=��_x=�c��($>�/p>��:��H�<�S��lơ�3,��U!뻓V������f��<K�����=D*�re6=�=�r��ր>��
�oOu<n/���;$�.=��0�%=�=�>��s��ϼ�@�%��=�p:�*�=p2���6��Y�c=-֭=��½V�z�^�*<F_9>���ǣ�=�|�=���S"��E������Uo;�iM��g�=u�e�|�v����=H_����NE>O��s59�2!J���=���5����=����q�<�%�:R�J>�r�;W�ĺt�:t��=�,���n= ��=Ϧ�����W ^=��R��9=��=����O��yڽr۽u����+<fC��Uu(=�m�=8�b=�H����������^����N�(��#�=V��=�/�=�Ѻ��`"�5W���\���F>��<�O�WS�=�.�xV�&3 ���g������&������zC=? ǽ��<#_�;�{�=��b=�Ԑ�Y��=*/��xZ=��ܽ�_�=��<BG�<�[�<�,�=;��=gm�=�ĩ��#�=�<�T(=A=�A��l����ݽ�2�������>n��<-��=�{�=o5>�SǽLR⽰�^� Y =�A���z�=� �{3���b�)|=8��=4�T�fÛ�QĻ(V�����!ཱི8�<�E���V=��8�AP���j�~�>\��7�y���g=p����%�=h;�\��=�wr�+���I�c=-����=u�
��+0���D��6ռN��=�<�$ظ��$>I���y��f�z=z�p<����;��<�Q<?1~�Z[�-DK�VC�=!~�A�*>�_���3<�mQf���>+�;�"�s�;f����<
�̽���=��o��f��MMX�S!=�F=�I<�[�=��򽯒��(��>F0����D��=��K�W?��¥=,i�=� �{r�<f=��}���.�;�!$=��<>��D�������=�4�Q��<�|�Zj=gh8;i5=��k���G�=�-ʽ�4�<l�m=R꼬8=4����}={�(={Y�=*��= �&��q|��ڼOM�ş��>�\Q�r�#>,��=�h>Qʔ����=qX�=���<c_
�b����DY=��=NK�<!�<Ŗ�;z�i��b�<S�'��(�V]7�Q�i=]��7�ý�x:>�q��u_ͼ��%��Yx<���9Q���x��N	�=+�<�DC=7�>e��?�ҽG�=�� =e��������s��h�<���=~lV<+ >J�����)�K���e�b�-�=���Ü̽���=T��<R]���A=^_��ޫ�<a>��B�����M�����/���S��=u;X���;��tĎ=���r�G��B�<}k��7�Ƚ��:�=�τ�@d<��=�e>M)�<�Y�<�x�=.f�T_�=ɽ�=y'2>Z�����;���9�H=w�սtE�;���;{�L^�<!�����=��`;bg�=j�=TG�ʬ��硽��18����=�s�=�w�;�z�=0�5�};�놽~+Ƚ��y��>�>_�I=��>���o�=�'T=�I�,o<�Py=�!x<*=���@:<�>�)��o�5�$�H^�=-i����P;����i+��O�<�%J=�P��@�;"��=���=�˽
�=�m1����<�R=4U->��ҽ�p�~��=z;0 ޽�(>3��=��E=��=��������Q=f�q��~��iڹ=sh���j#<t��<p�a���/=!μ��>��=ۛ�=������;I7"�4��<s��=�W��h�=I!m��\�;5~=��B>�M�X
�=�� >R=<j)>�B�=s�=cn=gȢ=�绻�C ��,8��
�<�E��+h<Az�=&���3�<=5�`7�=8{>��=2=���S=������T��Vg������=겺��,b=��;���<���=��<z!�����=�7�_UP;h�/��>7<q�r���B\P:0�p�Ҹ<�>���撣=�����=�Z=�L��p(>u�˻[\J�Q�漑 j>?�Ľ����[��#�Ž"{=���=ڗ��&=[�H�K�$>�:=ƭ>ԅ ����=������3���W���=1Z����м��T=b_O��>@=/yG>c}�=�D���*����G̼�I�.s���;�<G[>� 	���X� u=_5:�R�����>���6h����=��мǋ����E<����c��=�SP=AY�8��;�~�= ŽyC��W��\>�˼�=4߼�n�����=,���:��='<��e<��G=���;��=`��<� =���#)������ &��ż��<�<�� ��}������M�=糆�2��=>�<v�<����<��/=<�:"=<<�;&^<��W��1>�<>�q�=�T�=zâ�Y8��K�=>�h�<�,<zS�Ќ�=�̼3H�=���_1V=�f��fv�<(ST��Y=���=��)�8�&;���M��=W�=:�P�O�.>A�=��@���>�"|=i0�]��<�c�;p�g=}E�\��=A��='tɺP[�<?}�<���=�)=  �;�՘=��9��<�ڜ<�a�:]�_�KK�=XK����=��;�f�q?��33���kڟ�A3�=�:���G<�1��'ڽ�S�=�Yn=�����/�=��ν�yf>�Ҕ��A8=�p=0��Z(G�hM��
�<'n�;��r��od=O����ʳ��aX>I�Q��Q%;���H=&̼�v ��ݼ�:�;#	�� ��L_��L <__�=;����=���<��P�|*=O/�=쳅=�^=i�-��17�s�D����=4$�<r��==��<=P���;2=z42�D`<�A�=������V�1��=���=Vv�#��<d]��z>���<���-;U�G@v<�`��|)��y�u�Q�<w~=+���ꖀ=L�׽�L�=�&���F��
�=�����_Ž�p��?���;9�m=�p(�*`ڽ�=���<���=7�;Uf�=!)뼜w$�t��=� l�#����=&I$<������=�r=u?����O=p�Y>D�e>P�)>��=�a��tS�L��lL�O��
ȡ=H�<`��=��<�H%���)���<�6^�8�m��.�=�AϼE6���3��hȽXٚ��>�8��=�=,�Խ����qW���<��<�Ѥ���=���e��=A����8`���<����=�%�"��<�ꣽyÜ�1q�=77 ���<�]>��B= H���oN���=��@���=�%�u;�=m4)�;-=jZ���<�x�����;*�h����R�����<<w��܊o�w�(=Fzt��0@��t���d�>�=>N_ݽ�ﭽ=<8�E=<^�o��X�:OR<��=R��<V�"=ۋ�<`I��h =��(���<�Ľ:�=�Y=�zc>� ��5����<��=�f��""<���37���L�ໍ=��=	�M=�ﯽ�=��=��2��;=�~S=3f�=k?Ͻ\Θ=���=n��3�:��=t�&=�X�� �8<�����:]=]�)��=dD=!GȽ�~��p�=L�P�0<���:*惽���@�s��x�=%�f>�%=z��=��A�:l6>@V��}�<m�>>$EV=�7�<�T���H�;1`5=�C�<�k
>9��=U��fv��E����<�z=ѝ2=	��<@
�=�M����=�D=2LG�G�^��q�E��<�`t=@�<:|���>>D^�b(u;��6�~�S=󁰽XkW��}ֽ� >$&���=�p�<�#=䘅<�я�Ⱥ��w@���Y���5�0�k��^h=iO�i�����]��Wi�V�ؽf	�=}�p=l�+�.�=��/�ح�=��D=�(�=�����PG��*�=�e�a�;��<�뼇�q��m��L�[=�}>l���F>z�н��
��Q�l�c��=R����i�N�e����$�#>II)=��	=B6�����?"���'�?7��v�=�O>t���6�=��;O����x�w~�=�_q��M?=���=�J�=F� �)���y�=�ع�Lf_>�����}�i����`�b�E��A�=��=� �>��=�FY=��=�L=Ͽ=�2>P�:�==��ͼ���<{�>������%�� =W��=0S<=�]����=�w��	`�&��w&�<��>傸��JG�k3�=�i��Ӂ=S8�<f7~��,<�g�=�Y�<��<?=�=�㽀�ȉ��l�=s�<�$��x^&���Թ��4>���U��<���4���ૼ]f���/��lۓ����;���<�?۽��A>}3��\;�:�n�=ei��h=CE�<�&y=Rsa�f��
�=�����`<'N�=���xj�=]{<=��>|Sʽr�=��W=~��<�x�=u��<`��<Y3�<�>��9��%�c��]���C,��l�<�t,=]��<*�����=�����{�bɽ��;���<�\&��0�&�=�V=��m߻h�=%%�=��݈6�;v2=�*��x��ť;S����d;�0�=r*�<�s;���]�6�RĦ=�ȓ������<���)<j��<�Y�:��<�ڗ���=����4=0'���WQ�j�V��۶�ԭ�Í�>�C�53T��C=Ε=�h8=��<b�=�B��?2E��PR�V�
�y�H;�~S�=�m�,��ֶ;����M�=�����ɻ5z�=7/�09��~2��BN���b�=+��!y=��<L����u>�S��"��O�;�ض=�=@��Y�j=�~�<������~�I��om�;�6=��>�d}=���8�"=�]:�ؿ��[�=�o?�0���;����<{=��d;<��=�z�=���s��S�$�:��=d�z=��">ڌ�=$7ͽY�>�!d ���=V��=�j@;gM�;��n��[ >��=��]��_>=N���y�ƽ9�>=�V*���<���y�_<�1���<��t�BK������ܽ�������Vl%�I��i���mS����W>�d�W<�>(&M=��-=�2R�����6&�^N�<M�P����<��d����=*̑=� �<���[���r����<)8y�\	�=L��Χ�<� �gE>81G=��!�	�><8�S����=h��<I@8�r�I�qiG>�-�<�w�=��V��>���<����*>��ڸw=�/ż��+�������.�'�<�9[=v:��H= ���i=����;<-�=x#�=k�'<R3��P!>���$i=���<E�+��h�=m������n��|d/���>3�>>J�W��)�<0�t<(E�]V[=����{�<��<4�<��;��G�p��(�A���<,��=����>�O������
;�@�j�ǻ�Q�=Mǫ=�.�=��	����=m��=��
>t�=��=kf�=�=��=I�<���м��C�p��<������<i���H�9S��G��=3�=p��<��;}d=���������:̶v<�Ͻ�0q�(>�b��;A�;���=�><ٱ���U#�����+�'	D;#�=�\�;��j=3����=:��=}W˽�ս5�=7�;=T�����<((��{w=O�=���<�9�)[=�f��� =�4������l��2�n��Oc��+���L=��⼺ő=���;~>�#>{-ƽ�<�����=`�<�Z�;���<� >�ݽIƧ;[^�=m��<���=��=��N�rٝ�6��=Q��=���Eg�=U77=�h+>R;a��=�Y�=�'=�D�=���=Z+4<�]��:K4=挝<r�����<�md=�)ɽ^���&�<����о�]������<�S:��x�ӎ><}�>�b:>_�s��M=�R�<�ǁ��S�<r5x<^B�1m�=��h<��j=k��=⾒;���=��>��=ܝQ>�[���D�=*�H����ޠ�<1GA����u��=�x-���>�H���7���5=R�<=M�=DŽ��=���<����G'����$g�*)�<_ >Ӳ�� ������Z�i=a�=6O=��\;��!>�S��9���¼331�X'=�{b=ZWڽ�*I=�Ѐ=R����N��;ݽ6+>��[�+�==�DP=w���r�d=�䛽v0�<$:�}>�､�>��k�>��=��c�Ȣ�;.��=[c���p��u䯽s7=wˈ�[!��u��<ꀭ=�b��+�W�9�;�Ns<���=�k.=�^o������;��=^G5�2E$>jq{�/�̼�ϔ=+|Q=��<�.�=.��CfR=Ͽ>�<1c=}��=���e���UQ2�
�>���2^=���<���n�L5`�`&��ˉ<k3�=�ad��>��U=�NN����;P���4�=߭�=��t=�!>���=�X>�脽E����9,=�h�=�"v�5�=s�=��=��>	��=� <j3���"�<7`�<V�$=�3Ƚx���$��tƽ,1O={~=��:����=<��<M%�fa���9ɽw�=�M��E�;Gi�=�����?��c=-j=��R�o�>w@�=Hf<=��<�VM<�	>6P=ϝ�=�xy=���=��U��ޕ����=jv�<#>��;$����7��0�1�t�b;&�-���~=v�=�k6���{�÷�=����R�Զ]<5�r�֙h����=��O�q�=����N���;O�K���E�s��S���2��Q�<bPҽ=k�H�9����=��=c�c=jb��M���ъ=�ڼ6�=��w��)�<%�<M�$�0�_=Q�<ՑN�Sz��>�=�=��=%�u=��7���{�3��)̐=0&�;Y�=��q���$������Q�U���|����;7�ܽ����7�֘:Oߺ�E>�O����"M�|wҽs��=[�ѽ{q�����=�������;�Kؽ��9�>�e=�&=���	Q$=���M��H���H}�=;�=I�	>�Z�=�?�=Mg�N�=��߽��;��ű=b�b�$�A�=�>��r��5)�4W�'�;�:���a�2EH���>�����!��/p=��,���9��NüV�ݽ�����eý����x�:�-�<o�x<� ��|M���B>$�_I�<����:�<%��=���.B=�,|�Z7 ����� Y�y���
~U:;��>��>�����=�)��*�<���=�:�ih=�1���\�)9>� "�O�D;D��=�F5=�^��lhŽ��1����'�½^��<�cc�4���9'1= >�*����=�G�<�B;噽�y"=�>�:r�����BFH�tX�=�7�=FK.�/�4���<������=�۽C�r��-l=:�ҽ�
>g�R=�>��_=[*�=d&3���='�,�>p��:���<+6�<}�"���>�����J(<H}�����%D�ҷ�=ԅz���Z=ϊ-�&_ڼ�g�<fo�l�=� m=�=�m����o���e�=��S����^K�=��<!$��� <�Ħ=���=���=��k�z�9=rv#�x�
��<��*��=���!���T>o��8�l=?���-���:����8=����<r�<��ٽ h&��ӽ��n����<+�=����H{�=#�C=)�Y<�&
<�C�p��=���="�|�wU4>涖=�Cs<�M���>wx�=�C=�](��x�=W�ٽ�X�=k�p�w��=������>,՟<]8ɼ.���l_=��{�<��ν�[=Ѧ*��Ǘ=�<��Z�=��ڽ��½J�=��i=�޼��Ľ�P�<˘�=E���4�=�7'>��=�q�=r�.����bg'�} ���=���;64�=<=���fj���雽��{��ܑ<-�v=:Z�:B֒9jz�����~��)O=��=Q�.<?>�j��+�?�J�Z��4o=��>V�f�2<x�D���=W�㼅�H���置���)\���>>�ʒ��>�J������ ��Z W=�;�����=���:����.�w���P=��=J\=TB]��̼�4�<�6�;����Ծ���v�\�>=��U��R=9�3��kN=�5����2=�O�=�Ͻ?d�=y��<��&>����k@>AV����s=L��=,�<TnZ>j�k=�F>��[<�Y��"�L�qڎ<+8E>۬�=��<w��c<!�v���@=� <8��<��1� y<=^�;���]� �d�x�4�=rCD��>=V�J<1�#�f9�<j+@>�#�"Y���I���(>=ˌ��X4��l���<4��=�A��3=�=�Z<'4=S>T��=<�p?=���=�\=->Ev���(�0o=���=#�=�޻>����=��@=���=�:��m!���+=c����I7����x��� c#�˧�?��=|y�D��`"�R�{�������S��k�= ��=�<@<Al�=��>���=��ɼ�H���I��3mܽ���<�<:f���~O���k���&��쪼A��A��&6=���������
(=M��=LHg��s��J	���>� =�G=�w�=�.<=�����(=s�=��
�8��H>�>\n��c�=�q\�5��=��<,X�[�x=�>�=e5�=�>q=��f�%>~�ӽR�<���<H��=�5/=�2w���=�^=M�^�G�O��r��Pm<�=u�;�d��,i@���н�dr=V\����<�r���=���<'���D\	�~�<�w;�#$=,�">ٺ <�+m����<�Ҿ��}Խ6a�=��q���=�� >	<f��K�=�L��>>�ص����=I��=�a
=r�<�炽Y*:=Z�=��"����x4�<!?�����=���<6�2�7q���@��OJ9<Xu=~��=ߋ�>a���Z׼"�ؽ�Q=KW������/����K�Z��<ɢ����="r=�>C!�����>Zi=�#=�~ۼp0ҼN����=��y=��l+>�6����w�N��=�}�����->H�W�យ=<��<+��m�׽媼.=҅�V΢=c��=,�I�JW��$��>��=U��2׼��g=���= ��<Q|4> b��6�l��=�!ѽ8��=#�>�!>�}=
m,�����I/1>1ky;��l�nͭ� ��=<���bܽ$>#Y����=7��=�h=h��<�߇ �uV�="���RrQ=�ŻI� p�<���=���=�%�<��;��=ֽT=kYh<��=��=f1=� ��g��]�,�[�!��TV=b3��˘=m[+>EAQ�77�h���w�Ž�:K��h�=/�<�a+��V�����<E��=n�=M��=tS���'�����=+��җ7�����@���t�H䷼O�W��|���rS=���g�1=��=���׊*���;��=�������򧬽� M��M�<v�ý~2��"Bƻi>k=�{Q=Zwk��I�@��(o!=!!V�91=�	�;Tx���=�:�=��I��)�<����M�(��iP�a"��k�>��=�fH=�w�=R�۽+���7m<� �s=�7�J��=K�$���4=�3,>V��pP�<2���<q��<�܇=�k=Xߑ�RZ�<����$�����<+�?����=��M���b=���<o��<�0 ����=�	��i�=�̊� ��<�9�{憽�f�=�_��[ȼ4�սdO/;�l'=�|:�\>�W�;�Y�=���պ�����=*:a=<'7�wYm�G"�%U�=j�C�1>�s/=�h�=�M�=V�^9�aQ�͎=���=�yؼ7�=�/x�y}%=����~��eo�<h't���V��O����1��>�<p��6�:��<z"=�妼�q�,�!>C���&�սJ��E�<Qi��o2�J��=T�N��P<3��&S�=�?R=�$=r�d=�W��/�S��$�=��
><e�=��<���={��=d�<<�sf<�V��q�<��D�8��=NW��*ߢ=A�m�51�=h=)F�;O�"=�K�d���_l�wE�=;Q�;O��<M�$=}J�=nj�=��J���<��޽k�$=b�=�2<��=�r����A���=1&���=>ʨ<_
��'潜	����6�\���p,{��͖=4����a>b�x=�/>��=,>��S�H����o�=ɀ������⦽9�¼���=��=ӻ���>�d�*��]1�ex�=�^�<ّ����;�@�=�<<�;*��%���}��'��*�=E�����<��h<�B���M�V�=&��<x'�lJ�����vC�QO��b��=�H
>_ř<��<�\�;ZM��p����Io�=@F���=eY��� ~;@�">I{������k��<E��=�6���;ݻ}�>�e�f�(>�R>sI=3Ɉ���`�b�����Ժb&ݽ�槽�E�y�<�tB;ű�_2����t����=@&����<2B{=r�=�Y����=���<�#Ƚgv���
	���=��	��ݰ=Л�=�P����	=���h��	%6<mo��9��;��O`�zI����=�׻D������n�켘�y=��i��=J�M<=��@V�Vi��K�F��}8=��H�=W�>�=����H��=�j��G.�lg�=]����s��뛚���=�� =���Z:=�P\��(�=�����KC��;k)>E%ü����{ü�Ж�AŽKl> ?μ�>�=ɱ�<ۡA:	�νTၻ]��<0�<�仦��<�I�{��|�f�+�	=@٧����&9��1���f�=�
���c�< >şٽ0 >��Y=�=��<׬��2,<V��
�M�:�E=�h�=c)�=��7=����%-���Ƅ=�8����<|�E�_��<�)=��>o��}5�(��:Xy`<�_��~=s[ >J����<\]���X���[/�"�3�-G=����}�=���<F��uȕ�)
�sP��; �l=h�>���<g��<�	w=j����ȡ=V��<'Z�����=��>C$=�l����=�-	�rD�<JS ��]#�/�~<a�:q+l���~=��=o�>�+�=r w�L�#=Qt����=Z3v��u>����i�<�w�<U��<DoQ��A<{�<X��=hs���=���= ��Ij<NӖ:�޽�e�"=/� >��X;���=qR��HF\=Q�>�G�=vJ�Ԯb=h >6�����1<y��ܼ�<����V{l;��2��=�B;=��ν~]����H=_�����w<[�Ἴ{r<bԽ<��%���=��A>� <bv<��D=���=֧=��!�R��=��=i��=�#���j��p�O�I�Ii�<N�׼p;6@���N=��=.9�=2�t;GÇ=�h��qY=�-=s&���^�����Qx��*��=�U=���TO=Ҋ{��{�Rt�=O�ս#*A��<_��=&���7H{�e>2=y���i���W=�f	=����P.���[��G��G����-��!�b>P�@����V=X��<H)>4�,=T==88��Ŭ=!�j=]�6����;����J&޻D�=�E���2��{+�䨆�i1>�)=�O�<�L�<H�g����3=C"�;����
)�7��=�c׼�sżDս�v�<��M=�ʼd= mt�����[�~�u�	Y��征=�{<h�=����$�=+=\�<����Ȋ>�A����:��=����f=��F��1�ʢ�<�fƽQ��=	�B=�����<�C�=S헽�*=�'�m�Y=���\�= >/��=���z$,�~==,)��;�=N׽�婽��<����0N�	3<����iuP��g=&��:i\/='�ǽ=/���N=i5= w�����7>�cy= �=�o��x���>JP	>q��� VE��m�=W=�~ڻE�`���밞=~*<��N;<f���=����x/Z��й�/ŧ��t�B��=- �=�M�3��=�ۭ<Q?��Қf��i�2���wL�<�a ����=��G�bV�=���)�Ƽ��W=O��=]�m�5!Ľ7�=�K%��&�:�yX���d=T��<�;���`��\b��2Ľ�tu�+.� @=�k�=���=�g>>�{����Y�]=��<*�ؼ얓�P��
�����[�Jd�*�o=z��<Ig�g";���=t*�=c=
{�$Ƽ=(�>�S�?�5ku<���=�a�����<@ܽ������鼰'<�<*;`��=Y��VL�=����� ��<}����[�.����U=|�.>���p ?��$�ѵ𼭐�<J����=�۶=��=�󉽭q�r�����=
ՠ=?��`L<	�(���z�-wؼ�+)�l�<�Rؽ�R��X@$�;F�R�ּ�(U=��ҽt���m>���������t=���=��<�"̽��<���r�;�����P������[���Ƅ=c�ƽU= �=R�H=^�q�Nм=gs����'=-��=l:�<�<�;�5:;��8�%�;Tý(E��� �����9%>c���=S�1��$��������=�\=TJ[=��z=�!r<��=)����>oנ;���<�9>�b��g$=�A����<srʽ�߆����� �<
Ќ=�q�=ݝ>��=WԼϾڼ뼽�O&����<1�8=���<�)1�~f��$�=�Yۼ�v<-k�<�A����=�Zo>\��Y�=`��=�m}>���<Rf���	'�{:>�p�<�Ͷ��{����=S�<J抽qt�<Yc��9�>d�<�T�=�\�n��y
м>����A����;��a�<��)<������=���=�x=ϟi=�ʽc�R��;f�=W{�rT����=ŧ�=��=�Ү����=�>�=�<r�=���=r'�����=�����i��'�=7�ƽ�S=�zb<is�=�<罌�˺$:<-���Aɽ(��_=?Yx<�������=���=��櫽�,��ى��R���2\�<� �=�w�=+��=���<M��N��I���[> �ܽ�;'>g{R��OJ��E >�!�=Q3.�����½l�>�5>H�����>�O��'�>��%�iG��f�<Ϸ=w����-�<B)��Wt=!�!=�Bi��|�r�=_�V=$*�����&�H��=Ħ�=��>�z��K� <���=i�Q=iς=b`���=�}�:U�㽊��=F��<:&e<�34��*8=���<�ME<��<�,>�6<�|�=�,[�/���9`<^�������[�<h���L�ݽg����ϼ�,�;틽.w��?/
;�J6]=�cP���<��E=��>�R�<��l�]�!>�q ��H������"��Ҹ<���=�+�<�W(=(��C�=�����1=���B?��E޴=R|���ͽX��="��<��2����=�����7��x�<ZӼ�� =T������Ǵ�zpp;f܊=)L�<�m�j�>�Z.=���<���Sŕ<$Ƚ����e�	���ܽ��=��
�V��@�;=���=�!�+N=�=J2��U���㽻3p�3T�=�8e���۽zi�<�
�
����;���|,=��2=�1�߅<((������a�|<�%�=[bh�-�>`���n�=���=�ξ������2��=�x=׉|=)^a�v�8�:��<�*�CI�; b��L���Ǽ	ā=��=f� >�������=xa���;޸ � �=��u�(+>X��𿢽��q<�/��xМ=Wv3�_ѽsg�=�='=��*=�D�>�6=�FԽ�hX�@�ҽ��&�>�!_>K�=�.=��¼�sJ��n=�ѣ��ӫ��_~=��v���<�c	��`��\�=�o�7+	��t�M�+�z��8�<j��0>�<|�f{A>ip��Z,>9H_<�L��r�<�1=|_�=SZB=��9|��=4�=<���i#=5�Լ����Rj�W����#���$:>�5�( �=K�v���=@��^=�R�=�H��-���%�=w)v��Y�慾&��K�o��>���=Z�d��R���*��g�>��7>oH�<�-�<��T�:�=c}ý�0�aǩ����V*��@v��@=�'��4B��=�@G�KT�<J��=�����B�;��<���=I�U<�S��e���~�=���:�h�=
�o;��˽�'��{�Խƴ'=1bF=`����k��4�>�=o��=����~*=�k�0��=� �=�����t<�g=6xO��>>��=2󕼕O���z<>�v�>#9��޽>�v@�6q��E]�;���r����@�#��<ؼ��������	��<=��Y
#>�V�<Ǯǽ������ҽ��׼��
��+�����ݟ;夙;�ռ��:=z�=#OY��v=f��=��=��d����<��<���=���;:�:���= ��<D�M�~h�<;�T�r�=�ߖ��0>\�ڽ
�L����;�~��sC�=�zS���)=<8>�ڼH��<��=�G�<F�=�����@�=6<q=)��=��=�}	��v�=�����+5>l�<·G=�b<?�U�0	X��MY��Z=KЎ=��>+==�84��U.�&��=R�u<�n�<�}!<׷=�m��"?@��=�ý�r�<X?n��ּ��?���<	pﻑ� <ۏ;=�I��w�D���r=`�:	i=zbS���r=�=��R;��&�=HC��� >���<b���z����<>�>C�p=�g���d���>A���c���TҰ=0~���J>Zɽ�z�<�hݽ����y^�<�,��cp=�J���>�&�=�╽M�=���=6��o%2=�{=�D�<W��=�=V:���F>�$�=�����v=|�=y����!�==����սs�_=Ym=�\��?��=R��8
��ߺ����=cX2������|~�jo�=��=~�<�
����:�Gd��N3>��>!����/>�
���)��V��0ؼf�=R��nؽ��=O�A*���?	>D�2<Ъ���0��_��󃽨07���;= 8�;n�{=Lݲ�o=��=<�=�	?��.�۔�=�=�|�=Z��~�q��R����b=�;R��=�Ts:"��9w��n�=VC�,��=p��<h%@�[t�=�s�=w��<�x��Z�E<?;z=0k�<��<�/��k==�����=����3�T=�c��-�W0��>�Um�;���=��<�˼�;��{rP����=^��;K���f=���=����2��3=�Q�5�$;�q2�r�����==S�=0��=���=�X=���?l�=�h�=E����޽�Ȳ��1;,P�J�>�q��7ï��ˬ=��׽5m�<(�S����W��-'�	=@۽4��=��]=I1n�{�G����=Бc�g�e��̮�,�ļ.�zbf<u��~Ҝ��@�=�A�=:� �9�H�'�<��V��)->c����~=���������Y<t2)�b����U���Ǽ�LI;��W>�佸 �7!5��S�}=���J����
����'C<*��=��E��>�(=�^�����/�����>����=�� >wHw=�
�=Bc%�aWɽ17�=G�=�m >[������>p���I�=�8>s4��Lh�	��5�J%�=��@���O>.����">q��=��>d{�����?Y<�S��򃧽��&�/���g�=jY�=}���*�]<)�G�Wp�=Y,ʼ�h񽵍>ӭ/�5�=B�Ƚ�)>�<	n�<B�M;%��<��=&�!��'�:kF���������x�-�==v�=�)��9Y�=�x�<��)=���;��<��˽v,4�E��>�����?��0�x��(C��>�
D�;=U��<����&��_C�<(J�<{8�<�W�9g|½XnW=F���L9�<��U��4����=��;>�e�u=6����ν��׽=��w�F�S�=|�<i�/q>Y�=��C=1*�={6�=`˼w�F�'@���޽!�/����=̖�=��	=b�� ����\�=��=���<�0�=��=2<�=P�X��<!=Nƽ���%�<[>O������=��>>�3�S!��%�4=�≼g-�	�1������3�;� �o�=��ս���������-=�[ͽʂv<;������D�=�r��c���==�Z���Mm�M*��i4�;FF��4�=���QM�����$�3��AF<�����<���<F����<S�Z==��=�ۃ��!,=��v�&x�;��<mj6=7�"=K\=�]ֽ���z���@=��b����<���;=%�(m���'=�#=W���~�t=8>�Iʻ�AS�4Z4=��Q=A�;�P��>��\���W�i1=z,=�!D�Gt�O��=�m\=�W�<�a=�Ꞛ=�1��i���5����=�n.=%�ս�=�L�=�9���̴��u���U=�.+���ҽo�����O=���=Y��<��g�_Ҋ=+K�=钼�_�<jֵ������1�N�缝�Ľ��2�,z���� �q��<���<���=
P>
>�������=Uq<�ټ��==!��:����O��?#����<�(�9�r�~w��=��?�� ��(��]Z��ӻ�
=�Y�<����sg9>Z	�<~�%�Ͱ��@�ʽr���n�=)W�/�D���N<Q9��g�=�Ւ�l�;=�&�A�<�Z����= � �lv�=��<J9�8�">�G=���=�ȹ��"���=V*=M�&=a`}=�7=���=��U�tVQ=���-I�=�= N��iI�����=R��=�J�=�����R�<Vޭ�Ս-=lF�=�e�<#���/S=*��=�B��qF�_�D=l)O�i�r���x���~=��p�Ō�=�H�=��L��)<A���#�~�i=���<�a�=�ʘ=�1D>���;��<%E�=њ��a���)=�n/=���<U �=�����=�p�=�Fs=�(�<f�=�]>*(��O�<?&�=���wf>�O�<�rR����<��);��Ϧ��}���k=x���]� >J�4<��>��(=@����	�7�,�� >�F��V��;yѸ<m��<}�#z̽�.>�%<A��mǽsغ���;�pJ<�v�jiZ��꺏�=�x?��P\=�=ք�<�c�<o<��=�4�<)t�:]==���£ �^�;�����������1=��d�LLܽf)�=wg2;����o��G��S�=Oٹ�����p��z!>�5A��[0=�����>iK꼷U»#A��̎�%�u�������;�3�=� ���ր=�0<���<�oν#�=��g�����{�<��̎<���<C�`=�4Խ�Y��,D�=����1��<��:Ԕ��M8����+�P��=@Rt�����l@R=D"����;5fg�������h>�M���(=�:��g ��� >볔�e�<6�c�p�ݼ\����o�=�=p\̼Qso=v�=��=���98���. �<6��=CuӼ0���"@������_;����.=:st=� �=�R>n�H��&�D�}=_6}=�'�ق�ƌ=�}:�k���Ҋ��gy�-�6<U��=J�J;> +���Z�	B=��{����<ps=�u`�=[�q�j���<��<��=�b^�Mh��Tr$��H<'��\��=�U�I7��U1�d> � >�;��D<��4=�Ox=xjɽ���<*,��a�X>��=<¬<�3=.R�=��T�ߋ�����K=<�Y=�T�����<g3>��>�[�;$0��"�PS�=q� >�нlzT��\ɼ61I='�J<��������b���=���M�н�M>FtD�)�U���o=�ۖ=�F`�v��=�!��Y�C;��>�}���<�ͩ<uU�=��"8��!Y��N�=��3>
>5�}Z#>�Y�= ���|����Q�=Iu=���=���;v��>�M����5������$��H�=;�<����^%>�l��[��j��Z�f=���Nf<7@#��D=̅J=z�l>|�=��9=�L��RSս�[㼛c
����1 ���=^R�=�h��M����O�r4۽VǼ�D�=���=4�=�<=k|�eSl�(��=ҽ��BN��p=���;�b���j�uT�<:T�=����-f̽|��=�����;�8>0s=�=џ̻��=�҄��z<��~=��r<�Uѽ#3!=a3Լh��;��=?w[�ec��{O��?3��.���=�W�=��Z<��ȹ�<���BF��m�<��ּ�b7=e���}����9:^�2�=8o���z��x�I��ʛ�=��;=�==#��=�=��$���W=sF�=)x�)S��bd��W�?'���T=t6���L�=�Ma=d6y=���=vi���H�=�p½���=��|=���=���<��J�l�����iz>1�<�6�=|��9��=�h��A��S�;�H=�%�ث�<~+=���|���p=D4 ���=b�Q=���=l�ܼ2�=�11=y12=E�;b��h���m	>���=���=�����o=w��>i��Vؽd���Kͼ���<~���m9<se��E'�=841=���=�)ҼxI�<��=g����O,>I���޽'���V�E�9�7�i�R=؝B=� �o����&,�&�L�Jh�=>5���7<=�b�=��-=�ԽtV�=|��=1<1�#>�m��������Z���>H��<?�"�9���g�=D��<�_=+��: G=��V<�z����RĽ�V
����5��=�Y���=��f=g��=/:�,�ʼ)���]�nѼi�Խ�9����1��{�=L�#=��6��u��#�:<=�/�Ϳ1�I��=`1�=��<�15_���f��l�<K��뼽��b=�U�=�<���H=� �=�
�I�ۼȬܽq0߼ʡ'=7�$�5k�=�_<��f=F-��*�r��>����l�4=�#=���=$�z=e���)��='�FEG�ܚ�M�=0>�zq=C��j=�>��bZ=��8>lt����L=�A	����=�~l�S<�o=@�̼�e�=�1r��==j�=�3Y=d�=��v=;h�<�#�=��2��j��y�=+��=?z=����/,��H >�޼�/>#�5=�l���"�/��<^�W�;���\l�=	��`>�6��=��"=>X�=7�=�X>e�b=B�i����= #�ݸ���� ����=D	*�!$\�&U���s<H'�=˵�����=�ļ?Ǫ<�н<��=����j`�=X�!<2�E�嫄=6.�=�}S��`�=6�=�\=M�ƽ�Э�Ҩ���R�<�=�6�����������<��k�U�������=�`�=�o�i��%T��mN9=�$�oL�=���R{���j(������6�}"�=����F�=��˽�>�rs<Q����Q�>o�b��ؼKj��6��=��_��Ks��h���̹�꽏=�]�=�(q�1��|�=�ڥ=&���U�=댷����4�=EV�=����M�j�@��e9��;���ʽ]����_��n��<T�0���&���=T�<�,!�s��=I�a��	A=+��=��=G�+����:�;����^�c��>�"�=֊=s=w=�9����=B=5��=.b8�Ҽ?�4ҁ�S���,�?�=�6.��m��RL�.kA>b��<*Y=	׉�h��)��<��f������E��i�F����9ڽ��}� ��Z�=9�=BƳ<�/}:؛ҽ�?漣��m�D;t2ؽ��<�!A=' >^��Kὓ �<��'���w<>��=��|U'=��ٽ��<0U�:���<T=�RI=}J{�V�a����`z����>σ�=��~��!b�����"��.��6D����=c�W���M>i�<��J>W�>�?)<鬖�%uK�>9���i)=�	{=	IG��G����=�ň=)�8>�r����ƽ,�.��ü�>���;kU�}]�ǘ%��I=�,�=�\[��<�<�o�<���G����>p�=a�t=��;��r;{}�=;~'<_�j���=V�=��s��LUh<��=��=M�=6��=���=Dm�<>51=��>��0=D����н�Լ��=*~��!Z_�ڦ�����H��:���<�� ������=�ϒ��O½hN�=}�x=�=��S�����=�@��P�����<J2=�x=3�h= �e=�?�=�ւ��R=��O��|�=2V~�1��2�=�k*<r�<G?	=`��=(��=%rŽ׼4<ׅ<m��j�=��@<�r<�`�=��8>�qϽpâ=�X�>9B<�S�<CxA�T��=f���'0<�;�=u��=�E�{��m��=�#<���<��}=huG=k��=qI�=h��=����=��d�<Æ��)[���e�<�څ=���=ەY=$/>�s >@83�!:+=���<�:�V���g2�<Q��(ǽ�&!>s�����<"֯=6X���	���<"nܽ,�=E����웼�=����=B=G\L�L�=Wd��,�Ҽ�Ủ\R>��<��=~)0<��;S�R=��ｼ7�t_-�������>xD�<�6�<H��=��%>��t�KLU=*/=��j=���=�m<mk����w=MX��"���={�<��=ukW=��ǽ��ۼL��co�����C���nS�1e=y1�=f~>l�<L��=��%=^�׽�pd������;��ƽ�����#=���I%=��K=4��=l��ZQ;���0>��н�T�=��[����<YR\<=�
���8>2�.>osĻmF����=g@�~�$��'�*=������<�1=<z�� �^c�;�[ɻ7��<�,G��=[S�=�->*'�==lG>s�H>B� >��|�@<5�d=��L��%��l��Z�]���@Y�;f��0�=���:m�����*"t����v��=�`�;�=���ZV��Ƽ]7J==üi!0>� �=��<'�(<��w=���)z�T�$=~`�9?Da=3Zc��$���=����tԘ��ķ��hϽ?��<�p���½n��=Z����l�=[�5���Լ9�`=��(=�=�;X �=l�=MZ��|V�<皠�.X�<U�=���=29�=f	���+����D�M�(���=Ǜ�� ς���ڽ2Ih�5��Y�>�wg������=i��È�/�/�r���4!>���<R�z=dC�=3�}=y�z=_L�)�o=��]=kj��yټa�h=���=M��Q,%����`�Fֻ|�=�̼��@*>�G��]����8��.�2�и�=W=�"�=r{��G�=�5b�?��i�<O�=�2�=��V�]�Z�R+�<�o�=�9�������A�<��/���h�vp];;0�<o�R=l���'D=�w�=�<;����%��=,+�ij^>{�=
���45�O���Eƽ�R_�~p=`u=���Z׆����<G�+���Y=5���*��U��=������>:ॽ��8=��=�k&��CU����=�6�L������i��Ө�=�i���<��-�ՊC=��ļ¬�;�>|�O=N��i��x�w=b����A=.�>� >�`G�7��#��=�Ad�l�н&�=*�8>C<l�2=����^�=,�񻶾��k�=��U<����ã�
��=)Z;:��|���B>�]�<�8w>��==Z����;���=���<�ʎ���/=&N�=���O��<i'T>�ýEL>r�f=5u =����mR=��̼��=={�=�S>D�;R����G�<�ń��4��l�� 1<�5�=�v(=*f �{��q��H�(=^.�<m��=B�-�<�s���Tx�u.�;&K=p�*���O=��<�!�=& H���<�>���ﻁn��a�=���:h�g���6=�zI�"lм��Z��j8;���=c|<��>��<e�A>A��=W~�=���=���=�U����|�=�=7݀>@�	=ߊx=���:{ʅ=My�<V�=��N#">�2�=7ߴ<��m=�$��D����U=�`z<��=�A/�\U��l�`=ek4�ͨ�<�b[>	2�=�~Ž�����=t���v,�=0l��{�o��f>��=��p>�tֽ�ty��6= g>(�<����h��_�'�|�xz:=�!��I��=�=�� �:d�1%=`�_�n:=R���+]�:D�G��G��a�4:��<�a�,��=yΰ;zБ���!�<��=|��=i�=�6��7Q���=_�y=��<b�1=\�Z��_�<o�%=Ue�=�ֽ	U{�F/">r��=#^�Z4�=z�;���=he�=�ɽ%5>��y:�c��=��=sc��A>��_<'м �<�Z���8�=�5
<4�G�傒��j!=i)=��D=��ۼI���4�)�\=��$��Y^��>#���=cU���=T%���=bE��v�����R�=)��=�gE�p=
�;�r�='��g`�=TW�<�;>/���ue)=�=�Ա=L��<�r��q�=>hs��6=QN>��սh?=q�L=p���p��=�0D�g_<���=��-��|�=��<�3�=��������c9u��H���]���/�=�f�=��:�G=������0���#�>���>���;��#�e�+=��==a��=�p�=���A#>oC۽�
�=-b������h����8=Pҽuk�<K��m���᧽��=�d�=-?�=>k��>�;�B)=7i��Ke�y�V�˛�c|H>��<�W`���.>��=�6 =�>\=:���b��
�=@���н'����Ҵ=��d�!
>*6�=�IY=ҟ�$�m��J��C<�5���@>�7p�}r=���<L>��ԸS=�`N�*��;"z5;�p����=*2=*Z1>�V�=�2�=so� O���>��=Q$�=��S>�M�y::=�>�9->�#2��"�>w�c�w� �j���~�G%������3�����<8������<X	�<}_�F��ҷѼ������S�!�=dϼ����-�x����=��e=R
=����|��U��<���'�g<J>���9�:=H��o�<:]�<΍]=T�e��E=��;�˶<�ɾ<E]k=@s��N�B#f=CL��\� ���<+�̽���=�}�<Q����@�����=�]��l�ʽ�c@��?�� �ڼ��>��71��f�y��;��e<�U�=*���y���N�����<�u�=��=w�n=9���f?��?T�<��U�,�4�8]=��μ�j�� k��^����2�4Җ���G���;�<��=Fr�=Pl�=c�;��<����n=���=�k�İ)�#8	����ЧZ�5�<���*|G�p��\�нaB�:���=��5��P���i�<�ӆ=�`�pr@��L���lؽr
P��n���T��@��=�[���,��9��-���Z<�~�=�݂���=��	�b;ٽ�Q=h^����� 3>Ŕ:=��潡h!���<^Q�4��<ϝ'���3=���=�?���0һ�� ={s��@��<��&��1[�goԼF�=99�=��->���>�Z����>_z�������M>ɖ���<����=>y=�������o�=p>Ҽ�=�ʽ&	>���Y��x���{U=^��=�C��,>�[�=S?�<�*��R��)U��w>H=/@r>9�:>�_3�"��d��<n{�<�Q�=r(��=`�<�<5hT�V�4=@>7�۽�2@<X�=xvT=5��T��aR�:cj�ڂ��`�J<��:=�4|��+0=<D�R���O�a�o=��=s&�=�H�=�^���4�~�}>k�\=M�o�F= =��;>��=�%�.��Lؓ�!��̳.�)�9=l��=ּ��]=Y{��m?o=~����c��H�;[�{�n��=_��I���<����@>H��=��>A�-�x>ݩ�=�5�E���.��Y�>��I=����\�B���Z{���Q�:=�%=�<'雽ˀ=������+I��r����=��<=�Y=�:��ϼ��J�P �<� ��N<k�Q���[<�˽�������<)I����=��I���<�3	��ς�~G��z�5��=���x�J��!��h@�����ٮ�=���0i��=B�νR�v>XҖ�/~�=R]�?�7�;N἖"��X0=�k�;��m�OS�<�4��n�E�^�L��h�����7�=AL�6Jc�Z�H=0٠=�Y=sx=1ֆ�$�<���<��3=��;��=l�>���=2�ý|���>ʹ=e��8V��=,T>��>��9��R=r��=��5�;�$<Zʜ�SC�)O=�N�=PX=�!�=���<"�=R�6�p5�b3���	>W��; Ǯ=�D��Qx8>�9T��Z�<,���uӽ'5=�9>NP��Ϋ�I�����<d�^=*�½lz6���;�����Q���_⽜,R���=F2�����=)@�=��<�f>�t=�oy=�!#�޻(�؀=����,e�=+��<�2�<�n�=�o�!��=t,�
�׼��f(���z�=p˵=���<W��=�_�����b���?�='����6�5��~�?�ʻ���p�=�G#���%���>Y:�=iү=N�K=%�>����p���U4��(���O��+"⽣6=��j���&>�==�>�ʌ��!=<��<��;ԭ�<��ĺ�_i=�$^=Ri�� ����<lf���>�]�<��<T��
�!�Ƈ�7%!>"k����oA�<�;|3�HKi��h�=�#+=�� ��=:-)����=�9;��G>�v�:�	�-C�u�6�s��<I�c=\�l��Z%���=A!=%��<$s�q#�=Ö�=2y����ϼI�U<��=t�	�N9>��>��B�=������R7>?�>f��=�v��X> mI�U�{�7n������x=ƽ=d�A��ֻ�9j���=�XY���<��7�5=����E����9�lg=4f�b���c�97�G=�z�<+z��n�<u~O��@=���<IP@;�ҽ>��<25^=N	�=�[�=�Mm=���`�=E1H�r��Q��9S=��K��$�=}R�<�F�=^�׽G昽[m>��>�W6���1��	��Ռ�<�4=ŢS=��˼tĸ����g��8��=�2=j���g�M�V=1�~=��ҽ��#���=���:�y�<���K�ٜȽ=�XĻ�h��	�=��ҽ[@�= ��d�����=�̱�X�|=�l��g�c�]��G�^�fk:�D���n�V�<�;=�(�Mڒ=��G�e���u�=��=ަ��̽��~���:;h4=_��=��<��<L����Ѹ=��6����=�P�kU�=;9׼l�yN�;؃A<=!߼A�=������]>D�=�~�<}�]=>/+�� C�ۣ�<,�=x&(:|�|񌽢y�=^�=����D��߹P��,�0�0=�(J=�}����=+��=ITk�ڳ�=4c��K��p����X<�)��=>?ػ����<ٓ�<ǥ���|�<_��=<?��E���o=��
=�m.>��I|i���˼w�q���;U%ʽ�\�<�$=�1�=[��=�Q;CA�=������K�Re!>���%W��\�r�4=>̻=����Μ >H�=��(�٘�=�B
;���=Ꟃ��\Ҽ��<�:>5��NL�<��?<���=�N�=�)�=/�}<��7=��<��=�ݫ;v�?<i�>�G=-�J=v�s�L49��c!�j�==O��T��#	>-C�=)@�t?�=qg�<L�>���=/}H���>{n�����<8$ҽ���ɗ�=S������=�.�=G�=�}W={�.=n4�<�n�=��_���=��7>_��=�=�=Y?�'G�=8�==/�=�h1=r�(��#!����<�<��"ܽ�J�)�:�WΙ��R�<�@�=� ���<��W�g�A��=���;G}.�$��"z��&����c=�T��.���<�.<���=c�>��g��5�=��=��<�����%̽�.���Ӌ=b���by�=�� =��=gWq=2�)��M���<�6#>�=��u<?����a�=�T�=@�	��F����<�B�<ZV�;��8���}=(F����&<J>�=�l�=�y���3�y��=M=>�b�&��=|���u�$�b"�-©�V�Dɚ�����������D�."@�@u���;�F���K1��:.�I
>=�~Q<a��=�1=�Ҽ-.=>���̼�O������b�=��=��s=��Q�
����=�?�m�M=�Zw�E]�1�ǝ�D�x:�a+�6��;c�;"o[>�=���<�*��ՙ#��f=������+<�q��Z��B2�-i����o�����z#����<,�:εv�s����T=&Vx���t=�����W<g8��]"���釽�!�ߪ=q"����<
�O�ȅ<�^=<F�>f�<���(�<��Z����=٨��~^�<CA����=z��[w<��g����=�!�=|�"�=+=9=	�O�V���G7=p���������=��H=�N�=w��=@]�=n���O���k=�}�=Yr����=���=8@���}<=F>%�=d�=���=�j$=ki�n��eZ�=��=$־�\Ps��<✽/-����=��N�ܾϽ ��^1I=��;$H=�5��bg�=tj'=8���1���,��=��r=\]�<�>]�;��꼟�=�'O����\�?>�x��;(�W
�<blz�^6=�,�%��<�i�=e�2�8�=�u��$
?<�1A�퉴;TǦ=�Q�n��<��r�\Ǌ�E���S�����<z+ >fs���+�=Ң�=�����G�F�=���|�F>���/g��ʆ=pK������x��=�P�w\�=��ٽ��}=��$=�ػ�}��o>Tlؽ����y���*�=
��%��=$��ݦ�=�������=MFe�zNi=5=4�)=��=y(�N.�=�F>m=� �;�j<ș<���=y��=+7�=�\��&{;�$=��F=���`*��ʄ��<o��6�¼��e=L�=��<2�d<=6���[����<�;�k=����=�#�;2}_=�-�w�����=fi=0�C=v���e���@F�0�=�s�=8s�2���Cq9�{s|�Q�H=�v����=`�a=�TS��*����jj�=k>���2=A7���=���+1*�B��<�R��Y缞�7����=/;�<L�f=��=m8�=�����<+�:��>>�y½�˒=Ih<��;s��W�=������T:�4\��V���<t<h�s��5�=0�����'��l<=b3>����J��{�+>��<2P����=�RǽXl0=Lj�=�I�=�,��+ʁ<IW���B׽�6>�eļ/�'=Pj�7�>=���<ń=c�
�H�ѻ�}���;��V��r ;�r�̱Ͻd����,�;����Y�s��,��i>Wc\��Ǽ���>�S^=9<=�=^��/��F��=���=o�-��v���.u��wx��\M�I��<.=o�A=ܚ1�)Ӽ�n=|��=��n~��N�ٽ{>̊��h�/a�=�ܑ�I����W�=�i�=�Q�<���=���=D<�������A��Y�ﯞ��3*��u#=� �=O[�=4���-�νÖa�Ã8��<��<�=�ό��tE��'=c >�E�<B���<��=�w̽/�=�{�;BВ����=���;��,���<~�8=$���qս��><4����q=d� ��r>�,=�F�=�0������B����ࣽ�x2=��<�H��Y��=��<�M�<q�<dOȽ���=���=�Ͱ=�v>�i�a���F�<ѓI���c=���==D=��4�v��ʷ5=lw��^r�=rHd=�?2��!>�=A=�ST����=EӶ=�(=S4=�@���ow=�h�<��=���<e������R��=�:=<���=ه���w�G�b=��=n2�=���<���=��;���=M4T��rڼxO�;�"�<m)Լ�&�:#kA=�7������|�<��=��=l3�=b�=��=y���@=U0����>��g����<�D=$����@��q=��F=��>=�����%ݑ<0V\<�׀=;�>�p =����O2�=�)��#�=X��<Sd	���Խ`=��g�5��5������ʼc��<_���|�<h�����4>���=Cu=�ս�����=}8��*�����ɉ�=B����j��l=�=ǗW=Ҳ>��<6<�,��&D�=�=<�R;w<�<��)��q�=�ɒ�����9����� �;�>�=�Ƚ��8�0��=-c"����=��<.ō=u�ü'ݷ=� #��V]����8KC��1t�Ff];�f������<���;oP�����=�� 
�<<C��ǉ�<��X���]=��;�X^�q��=��ýy��� �R���cǼ��=��������-=@лչ=����S~����<�tĻ�8=��X>T�G>� ٽO��=�
A�H<�<�ݵ;��R=D���6��<'𳻎)��;��</������<P���k�ƺ�Í��7����=0?�)?����^y>��)���5��@�=5o�z�< { =�dR�d �K2���5>N;��HH����=�u�=wM���%;�š!=�r�=�~=h��=�?=�\��N�i=����ݽ�C�=�3����.����[<���=�R�=�I���'��,ƽ��w�~З�/��=1>��s�&2����(��=]{>��6�)N/�O <e�%>\%1�e;�I���j���cI��>�Y���pg�66V���t����=N�;��f�KZ%<	�5<��=�d�=���%x�����u��=��u=�t�=��ڼ6^V������=Mz�=��&=Z�A<�<A���dO=4��<5c�=Qt��r�=`���9�ż,m�<�>�=�2�=gh���O��4��m�m�U��)��x >��4����S*���YZ;�u��;����=�<>8l���$ּ��=�g[<�!>�K��t�=�34���=��P�gp��h}=S�t�hCZ�j8�<� ԼB�a;��<[��������施�9��?Ӽ�V3=���<$�<n�*��������'�����֣ۼv��=~|ż�� ����<rl:H=�e�<�x�<��s=��g��:�=1ѥ<5�=l����=φ=�#4<�0�=�=^�K��<�_I��N�=d�w=���=/�>릎����������t�)�u�K�؊�=��<�K�;a>�=��@<���X�����ڽ��E�����MÒ���?��ל�CE�=�s$��}�Z��<~��K?>n��=JT��>��2���Ү�=7�U=��W� �=�w4=�.���!�<�Z��u�$=�d������-E<p�;��$>Fߝ=պB=���-�=W+��E�;=24	���o��<�<�R8�Ee�
�C>Q�;j��݀="bU;��<��O��N�������9:��V
g<|����=;�=���+�'�%�X���ռH<G;��d����=AQ�=3
B=�A��� �=���ڿ̻6}���X��̻�j=@�/�꥽�֗��-(>���DH���W�=��=Qt��X����s��3O���o��w,=��K=KT�=x����&��ڏ���`;U)E����\ҽ9�3=���<����x�=?T�=&��H��d�μ)�����J��H����=D�2���^=��4���3=� ����=X��۲2= �d��d=4� >������)���=��|��r7���<��<�U&>�uѽK�c�ym�#�=��z=�=v�>{�=WIȽ{^����B�>9���Y��T�=�W��4�=���9�<��J=��6��S��.	�<$i^=§��#=r�l,����O_��0��=���=>P=1���x=�9<�F����&�<���R�<�=�=���<.�=c%�=ې۽�����G�_(�;�=3;M�FU����� =H���s�����B>�e\�=b͖<Y�=��=N���=�伩4��|=p����` 9���=gw�7���� �=���Z�7�|���AZ%=����,��=Ȑ��z�<�F"<�vн�̽5�#;=a/�ψν�9>3��<�� �L���9���0Ļ*a��ks�=9���6H�<&/�oS;&T>�c<	 ��K{���0�����*��ʲ=#� >xc���=>�W]�7�R፼�Hf�Ё���у=gI��?F�<\=e�;Q�л>�;���K�0>``��4D(=3D>���<��׽�T����&��C�=�>?��<5��+'>�Н����=���=|��<���=Er=�ǟ��˽��=Cm��=ݽ=�!=���;���<ǻ�9'��������`�������O��p��(�rt����:�
=��ż��׽+ =k�<��e� / <x�ǽ��y�pw��x�=��=F�@�i)=���W?=�=�T��=��|����<�K�=�aǽ&BK�u�9�������#�A>�P����=�C�=�=J=�L��Ώ >�l	>�I=lb��B=w=�aq=a�g���>��>Jy=�L#<��n<�����#=�78����|^���=�N�=�Q\=�F�=I�����X@!������8���=�=��-m=��U�=�&X�^j3�t葽]9��	|����O[<�ؽ@7�<@]>�i���ض�ɛ�\��=��= B�<ڗ�&ƾ���T<�����w=�0
�+7
����A��<,|�<&�¼̤�x�=�d� ��v̲=!�>V����W>�l>�Y=6wz>�鄽͠���8>KP&���������"�=O|�=�֬�+1=l
<=�\�v��=f�üSh�=�탾��Ľ�Z@��O�8)Y=U�\�O�����=��</
�;,�R���<SD	>��/=ʚ@=��c�M��<B�=��<=F3h=�J�:T�ֽF��<�y��M���Mr��w�=���=k�ݼ�č=����s��L��S���<��#>��׼\ r;����{�4��7�=X=к�<��O=�k@��]��+�^ ->��=-��<�V�q�=`�<��߽黳��T�L�к�0�=�w�<H��PW���B��f�S���뗖<����!���J�<���ݙ��L�(�Uݜ=�Ҽ;�>�]�=�^�����U*�H��W;=�>�<UR����f�P�t=��={��7�����=4���O=��]=�v@��L=a�<)��\ϛ=��4�,^,��i����������N;#�����H����7>ݝL�)���������Ũ2<�����><���(<�<�L=��f<�--��P��L|��i�=hk=�P=M(���+=�������?|�;a�μ	�=N:ý �	��x=���=���o=3��h�=�·:�;�
�=T=�&�9��=���s�>�RC=t��;�O����=�=�#�"�������=����)�=���=�t=y�������B�=)��=��I=%1��S�=k/�=8X`��k>�b���϶;U����ͼ��㼒�!=>�=��̽���=ҥd=_�]<�y�5�g=��6>���=��ƽ �=����<��8C����=�h=��,=�f�=�C1=Dk�<	>�<iz�=���^(�=�8��`�<ꉧ����o�=�������:��l��f= ���
��bJ�=X��C���\->6K�=�Q�Z"X>�v�;Hrs=���<�7=��]C>���=M��;�޵=9��=���<:r=��<��B�,[%<��
�(񲻥�[=%L�<��9����T�ʝ�=/�)���T=�%���\=�ɽ����^V���$=Ik%����=`�<n1��Y/�'T<Ժ��T�[=�0��8�n�b�T�!����5��b˽�Խ�H�ͬ��`#:=�T8�KO;=��b�D�����<�����}��쯟��=7=ܕ=��=�vý�Fy�~��p�*=Y���)����<�N;�ڢ<�޹���ǽɻ=bȢ=VK�<�^�=%ݏ��Ԃ<C�{=@t-���w=�y�=Df�6�Y�<1<=~�����=m�����,��`^�]f���8=�w�=I��=I�����=ě'>4�$�Pl���y�����<��#<�.¼�Q�=��n=D�Ͻi7��m>�}��ᤚ�o$�=+�;1#:�VaѼTsƽJK�=&�==|��态=H�<$0��F;=����A�=�8��qt��qhm=]��<�N==j"ڽ'h�_.�=�s<F���y���$;Nr(;!F����=��D<eYӽE��<0��=�m�l�=�5����l=�>�=���=�"�=�0z�8��<�
_=�4a�q����"n=D���I�=��$��,�;�m���E*=h��=͎ڽ���<F>��$�=ne�����=|hڼ]�C;�!"� %@�舼c���!��#�=���=�P=�=��/��8�=�潦ԛ=�*�=�>�<T�3������|=ު�<�C6>x��=�u��g�,�ƽt�&;Q��F �<�5�=���%�?<�X���|>�#;���	��a���;"��H�;�u�=��=X3�=v�"=L�=���VB���S=ll�VFA� �B>��Q=j�;ԑ
��,=�	h��Ў=R'���	�=��=����#��ƞ�=���?>����&ҽ�Iw��K����K�����k�B�>y�=Y�=~\=U�G��㜺��=J�=���<L\����"=H���h�=�>�f��#�<cx:����\==��ާ��_�=v�</�@=��'���	���=�i��Ѿ<�ҽM<<�B=�HP<���ʼN��=E�^�*&�s�p���n���Ͻ~N<�u�SY�<Z >�桽*">����P�����=xo=��#>�-��\�=}[=>>�=�n=�m=��<��=E�h=�=��=<)�=����/�=�X����7=Hٽ�p��<~N����=�5,=Ǚ�� �<{��<�'�֧+��^K<��`�y|=�ژ=�㾽����T�XkZ��f��Ӝ >�=���=vx�[N�=&�=��=Ŧ�=�:0m(�Z��=`�;C�=
��=_K�<=�ٽ�>o�ֽ�?>��*=Ώ���{�;�:μ��0=��=JԱ��e+�.�$=�Q'�z���/)�co��4hC������ӽ�X�=?as<��c=ӗ=s��<e����ȼ�Q���F�<A=�
B�׳�<�H>4�����i�x=�a.=NS�=�)��[���ֽP�Y<�������=_�<w�R<��=VEJ=���.��8t>�x�8GX�q�f<f��<W� =�ߟ=b�=���=�.�`�=�]=3���Cɽ��>��O��0=��м�>@Ȏ�3F�Լ�5��=#��<�U���8�-_�n��JS>�	�T���>�p�<A��|k�"x=M[;�`�=RL{=�-��"�=�ќ<�[�Y�'>�ۓ=f5���5>'!�<hFA��@�=��D5X�o:�08��U���;��eZ��T9>�=2�F=W�<�����6>�X�=��=��v<m��TgX<t�=M�
�Q¸��N!>��A>ｧDV</�ý��x��}*�=�->)��=T��=�Æ����<��6�Ub�;�ط=���<�f����q�ۻߋ<�F�����=y�f��'E>Y�
��<�ro�:4�=�L�?�7�l[ǽB�>�@���9�=`���uCe>�>Q�K�=1y�=#9���<Ɇ>>KB�Q�"=q��h�=۴Y<����\��~I⽛�>1{G>�0"�"�d=V�˼�x�=���<qXy�ѯӽ�N	��)Ҽ�n�<+ѧ=:PP� ���ę=`-�=/� �<*?&��A��i�>�v��/C�=^7��* >���=@M�<$j�=���ㄡ=���7�;F/+=�v�=]I��Jj�<'^ջ���=�ȼ_n��(�=}Kż��=5��=�Z���G���<�>�^�d��<��$ҽ�m����9=l��;���=�rn=j>>=��s=�aʽ����w� �+�j=;��=p��=<.{=>�=�$<h,�W&>���lGM:���u"���q�Q�ཛ����= �=G|�I��HZ��ٙM=��$=�Ș:����=����m>���v�:��Q0��6GC�(뻼�lL�S����!�<���g�W伎�G=��C=�FE��=� @��@�=�U�X��Cw=�臽u���0V��}����޼�>��<m,�=���=��G=��N��yF<H�=��U=PJ�]S�<�d*�*�+�_���
��B�ɻ���=z;׽��4����=f���	��;p�U�d��B�<t�>�n�J��VL=
R�=D!����<U���=��g���\�X=��=B2����=���=T�j=���Uo��ŝ<�Q�=�,<���=����,�K/^�S4<}���n��V�=m���^&�!'>��b�<O�=Dmʽ���h��=�������B�<f4=�cx�ߤT���~=є_�F����&��>�P�c�ўO��ؐ<�d>!<<�h�#M������),=�}�@g.< ���f)>g��<#V��m-��%�=�"�<)=0�<������:�C�=iB�=~�E<w>\m=sC�=Lf����'>9mɻ��m=ㄮ=e�D��#��Ӭ=/`�=VI>�a�ă���vۺ�\"=c�_=����|�����=Uw��g��<�6ļ�A?=Q�;M�*�q���=%�e����-�Ľ�	=�9���'��
�=#�%��6��]�����ƽ�T��7I��t~�?R�;2��<��c<���=8^�9����fˉ<����Q���A>Ӳ>kv�;k�Լ�uڻ����M�<�P��e��=�8ּ���=�%=�9D�S�d>�j��p�� ��B&>A(<��s���g��û=NC�=�^:O��*Q��eQ��S�\;�6~=���<F	f=Ӻ�<͇���,F=^��=�X�<���=�$>Nk�:�Ѽ�B�=_�뽙[=�(�=أ=Jνv[;�
	>�6<wz�<��ԽW�����=cX<h�>��=Ѭ���p0��n��.=��ŀ=�J�=�#�񷘽��׼E�ͼ���q��=է~=�|�IX��焽���=~���]ϽC�=VD�<71/�4�>�ȇ��8Ƚ�"b�N罄���h8��7|
�B�=�\#=-��1m=��L��{���}��fd�WH�<��><;�Žۊ�=�Lx��L���D1<dv콯�Y�ߐW=,r߽)jԼ��>�ֽ`�l=~�=M�f=��˽�,���
��
�<̴C=ˮn���A��~�>,S��@�V|ὖ� �93>˂t<�'���;r؉�b��=���;_��\&����<N��;�L���<��m���r�?���¼	�>3���q��=�>w=$c>9: ��{�=dF�=ib >��B���5=)���X;�f��m��=}��<S��\(����=#)>�� <AW&=�Մ����=���=�Ǉ�?})�G�߽_Z��{�=��
=q���5��=��=£�<3=��,9=f<��>��<��
=w��~���k��j�={ٗ���=�Z�<��k����J�<=��=�س=��R<���=|�=���=�`�:$��md�@p<ٖ=�w�<���<�	�<��W=j7��a�=�!���3v�$>�.��=��=�->��<�^!<��	���={$�������=��=��'>��	�C��=�SK>��˽�䙽�Y>�c�<���n2^��#F�E	���bG>W&	=wZ=�f#b�l�=�{�<��꼻��=`�,=/�=�����łJ��K=�>>�rɽ�X���W�=��ɼn�UKz��:�;a�۽%=�!-�}/ѽ:I"�D=��>=�A"8��=���<��;>�>e"��4�=l~��*��1$!>>-�;f��<�&�<d)�=���?n;o�I<j]<��
>w.��|C������=��7<��oa0=#�= ��=�t��q5�=`�=4��|���N���I���	8��s�=�A�����=\���Ez�=eT�GŻ�Hh��_=ɶ>�<�<�� ���=����޷�=����>{+I>9�=nu�<�*��0<��X���5�=<�=q�<��R{5=��%�⚽�[�=���̓�����=IU�;b;�=M����0f>��OǸ��>�
��qc>ћ+>Z
���&��,(>�=8L =[�=�y����t<�1>L��=;�~=e��G	�=�3.���)<�$E< fB���>V�ϻ2,>��=г߼��νCh�U���23=л�=�&�����=��������E����򽢰:o�=�
�=��%���m'>]Nf��=k¶��u1���޼��:=;t�;�;K;�ǽ&js=Ӓ(��U�ܻ��0(�=�O���ُ�_��<�F�k�>���<>A�=���=E�{��n�N��=: �^��<?T�����=��߼.�B��������9$lw=�a�<���<�;�=J;&�x�=�}�=��Y<�@q=��>�"�=Xէ;�7:x�=��%��K=��ļ1��=&��<)��==���%>떗��b=���=l�=X?�=g=�6>9�#>yk��0���=>һ����:Ӧ<���w����=P�$��L<+�'=�0�<���<
�=9������u�=Q�-=��=�庇=�����T����<Ĉ�=��<�w>�m�=fZM�-�R�R�=	�";9~"�^�s�Ju�=��?=�S<�#Y���<���<%%�#���������=�Z�=��m=wk�s�=�f$�
���Nл��5�4 =9�'>wiF�
wI<�8���=�X�=���;1dӺ����е
����ڥ�<4z����=�NP>x.�AR�:��;`;�U���Q��=[���ȵ*��DϼՋ����=}̖=�2=9��=����%���=��=�tλ�*%=�μ��;<���=��E�m�ͼZA}�§.�8��=��ʽ+N=t/��G_=�|Խ�!=�3���S����Eڱ�B^ֽ�G����O���>��.=?1�=�{�=�<N� ��!8>�>#�<������)�<8G<��	�=�Һ�I#=�Ԡ�&+'���<�a$�{?�[uo=��꽤8;�rE.��%=�ި�O���h+�77�=QU�;�f�x����0�oCY�p*
=&C��'���4��U�n=s�����%>h���-�<��a<������S/��3O�< �J�a� ����z���ob=F�����6��T>��˻u�>���[.=:�Hʋ�R�=��=3�����q=���u}q<Ck�='tx�����Ԏ�=����0fk=g�2=�T�����UL����=��v�~����QL�S�b=�7����F<èi:
q>���=�^��@�gU6<ZX�=�G):'���\��<y�"=�Tӽ_�l�V	�<�L��D���=�y�A�G�2=b=�s�<��晻�슼��;�=�Ƌ;&�r�����b=��D=t>|9>�+��`�'�qc �˘P�D��l`e=TK��*��=�W���~=J��@e�="�=���v5�H�g=ȭ�=�������<�����=`�A=���Kx=U^����=�RQ�����D�>�XD=����-�=N��;=zg�7r�=��7=X�Whd;М׻��K��':=��/�����=�@<q[��/>=�ZU>ǿ̼E�=8����`;�0)������ ��ռ��<W��k�v=8�W=WB=�;X��3,����<��==����b�q��)0�����Hi��z���A����4=v��<,eɹ�*����U>І�<R�>�w�=,?�=H[��� >�@1���U=���={�>�d+=L!����C=���<6꼍"�D#>��¼�c�No�-Е=u��-�>�@}�W� �^�c<��F=#��,�8��;Xھ���d���޽\sý�۽� t;�dl=c���c����ƽ���,�>j:�<�7>��; �{=�)=��=j��;;��=O�1=�]>|�;Xn��>И��򒷽N�ͼ ��@%E�6�=������,�=͠=E��=������I=i�<
�����;N����ˡ<�ý�(>Ɗ�y�<�!E=����U�"�j�=�<���;�4o���9<�C���LR;BW=��C��=��=쫉=��)wU<�Ff=�i�<����*�;˨�<���=w���o��5"M=C��Qw���c��5���">X�=Ɩ�=X�5>�����
>3��-���Ț�=���</{9=��޻C��-/�����:���<�i;�[�=�G$�_�=�<L�<�;8��}<�����߼j�J�s��;���=�C�=eψ�x�2:�[a=�Ll���<�����=�\>���W�<�=��<��FC�k�Ľ=���5<>�5�U�;���#�=��"�?��=R��=��$=AC�=ǰ�%�;�>�����;s�/��I����@�@tT���Z�{Ā=Y<S\��;g>��<Y�p<���=����'����*��佻?�f<�<t�>>"��0*>�^���<z}�8��;��x=�y��[h:^��=�lC]�5
l=#�#=�)�<:��<���=;�e=t ���gV=�̌=�W�
{0��B���<��ͽ�2�=$�K��zf���f=Oqx����>uG���=}�N<���<��=�Q������t��3ҷ=H<>#RM�������MG��}<�it�퐍� >�
��*S���㽗I�ҍ<$�=�*���8=���T�Pý<�~�V�Խ�B�� ��2�:;�<=0�����!:7Hj]�[�I=��ʼ��b�#�;@7����󕽫ǽܬ
���溗_�=4��fJ�x�-=�!9=�5���&�ybV�:��<d8ϼE$�<���=>��;�.�
t��}���u�<C��=џ(��oݻl�=Y)c=pt���i�"=��=�nd��x�<+t��Sr<�o&�?��)q�@9>����?o��5x�;���Mj�;H�=|8�=�����Ȣ=a�[���ܻs�v9>�퍺�$��4�>���>'�;�Ӝ�,꺺թ�<���=�ˣ=�%�;�����u����V���=�p�D�:�j�B�==�<�YY��mH=N3=@b)>>B�/r=�	*��F�<�һC۷�Qf�<n�!�Y6>��
=ݽ#@���*�<�<ػ����.�=���=>�=I�<�&0�&	�=F�����Ŀm��ǥ�*�=u����9={_>��=�J�=�ҽ,�5��>��u�;����P�=ajN��ǿ=WA1=�Ls�yyZ�Q�l��A[>� >X�=v�u9p��o�>�q6��;
>��<u�'�"�<
��<� ��j���=�6�=��p	>n�<X��;�'��[t�<p_�V5�=c�<��߼�@>w2k<KvL��C=[�3�>q��ȶ�>:��<���=C��=`��=�C�=Y�9<�t�z���3=?�1�W<�[��;M<ճ�n���
*/��s<���>O1;w췽~k>�a=v9<)F�pN�;��R�"����v�!�j���}z�=�R�<�<��'j��0�=Ƀ�=d�=���>덽�M�=��=T")�f� >7��; �q���w;�4�	�����x=D�B=����ɬ�<�a�;��}�I�J>``&�=U%�hmJ������;;���/��~�2�6�A:�rν)�r=�Z(��}�+�ٽ�=pP�=�Uy��,`�n, ���5�b)�\9=\��;�)�}H�=�l�=�!=tt�<�q�<�>�e�=��<�>�����X��S{�<Q�W<ĩV���#<���<��O;G2=#�m�7�2�=��`=p�>U�=Θ'���=�|��޼�c�=�m�<׾�<W�˼[�O>M�Ѡ_=;Z�= �
�z=�l4� Ļ�8���ݽȵm=	�>g)�4���3;���>�).=�̧�"��=��Q�<+��=�I=qt\=���;��,=�<�=�� -!�ז=;�	���E�@��]��6=@���t���c�=�'A=�k�=�x=mC�<%��<�i�;C/�	R}=��⽞\��#꼉}��1��sB,=t��=OR����<P��d�\=���_��="S=�"���a��u�=Y��e���-,��P@=R|>��=	,��="���������=�<�<=3jƽ�E�b���/�Y㾼!���~=�X�=^W�;0)����;�'<��f=�v'��L=��=R�6�%�J�ͼ�=Z�����'���=��=[o�<�<C��=MwF�G��=���� �x�[^���C�\.��9��< ��ѽջ[*.=H?�<��=C"I='�<C�ۻ?�ν�<�<X��<�����F=��u�w/�<EB����.�c=5~B>a���=��I2�=U��=� ������B=��=Vx5=o�X�%��=�>} �=���3���5=1�����<'I;B��<����H��=���=�C�<u!��u54����ʉo=��۽x�=�[��9�=��ߺ鎆�I��=�s>���=S�<��#�=.9��~ܼ<��<�ɽ�>n����k�=L�v;��5��Z�<���<V�O�>Ӻ�T>�Ξ�A���@>\	x=L~�;��	�	ӽ�=-�Ǽj�ܽƜ�������_=Ӿ�=����s�ʼJ@q�\��;3陼g�<ĺ���j=ۀܼM���#��=�m=��_=���=ˏ���&=�1�s�0��CܻF�#=��)��A��0��ho��s'���=�r��bp!��Ӳ�T�<�3��ȼ~���dj=�ŭ<$,N<�W㽁��<�C��z�6�g 1=��ǽ�ӵ=O:�=�}��r�=E]��ۙ�;U�M�O��<��d�m�^����=��+>��	=+<	��-L{�AJ���"��T�~X*������ ½�B�=���=>�=��7=bX�=��˽|��:"�*���h��{�<ؓ�dQ�=��<��<��=��=�=��������_=C��=i\*=�m=gW�IȽ���=uɊ<��<?����^���f<hf`<䓽6so��>�<�����=
�=����х�x�=)�<=A��O8��O$�oS��Z���v�c�;iJ0>����I�='"�J��=���e\�=�>\?�<�Ӽ�|;��G��s0��w1�F����7���=z�C�cHP���>!�����=�뼝@>7�%��f�=Ɔ��m9���O=� =F��=�S���S�*�
>{>ּ��u<{�����=���=`f���ZS��&ʽ�;=����~�&�>�^I=5>��=o�(���<X�
=(1��`=���=�㵽؛1=-)>�{�=K'L=���<�>plL��>�>�A������=��3<N��a=�9L��ރ=A!F>�B�=�EC>b9���;��e��ݴ����>�4>7Y¼Pk�=t���To=F����ˁ=0"	�L%<ۢJ����=��/</:�;m��R=�ͽW��=S��<��=�Ϗ�Uj=t�=�6r=K�=t<ܽ�"=���Pn=�l1=vB�<�kA=Z��<><�w�+��=`E8<�]ɼ�3#�|'��^��=Z=�sa�/�=�:n;�&�=�`0=�N�ߙ@<S��p>`���U=n1�u����]t=k ~����=$K=z��=�����ţ�
:��j�=�ʟ=���=����Ԇ���ꆯ����=�l=�����S�� ����/= �*=�*Ѽ]�n��s�=��>NN�=�	�����^=��=�p$����#���A�H��=y|˼f�*�:?��O4�=a�=�	<�Ϡ�]�O;�!d=T��=a@t��f���˽1Ȝ�dX=��=�9���ú�<(=@Ƌ<	�)>-��=e*����B<� �=�ף<������E��]�<N�p�{OR�v�=k��,�&��4�<�S=��>���
��=�ϸ<K&��p+�_'B=���=���m'U=}��EGN�w$5�b���=��`�-s�=�G��ؽ0�=��E=�v�=u�=P[�ַ�<Gv<�"?>���=$"���=p����!��J�p<��=h>�᤻���;P�R��л�J��^�����	���ݡ��_|��E,<�N=�E>�F
;���=J�<_��=�|���̽PR�;P}콄뼽����C��1�5L�����8�G��<}ɼJ���>�^< �����=���h�ż�AK�-������=.Y��\��R���;x=�M+<	Z�V*ڽGx5��R���iҼ���;��F=_t�<g���L�;Ƽa������>��=>�[=��/=�A���"�;�j��K̓<�S����x�O	=˟x=sg���E��|ν�i*=Tx]���<�P7���=�ż!9޽�:=�<���;��=`CD<|j�=���3�>[Y=�Os�=�=���9 �=���<��=�ȏ<k�p=�V9��8ǻ"֦���=k��=_��<R=�υ=mz6��Ǽ���>�j;yކ<:"�� �¼�c�<BL��S[t��Y=ho?�:�+�]4�ڝ�:�4ȽR�6�)�����=KѾ�=�	>%B>t����=�����<� >>�/=���Ӑ�h�=�}3�#�=jG">��>�� E>�"�=eu�[�<g����Ӳ<��>�p>:��=em)<녘=U��x�(��pE>Tl�<�������=s=	��<J�=�>3���ݔr<��C=6�=!�=<�::�K�P==&Xg���ռ_7���l�&k�{&;rn==�����ዣ��#>�`����O<��/��U-�G����h�<YU���=�,��v>�@S��'=�;1���e�=�8*=L�I�7<��i�?��7G���#<��,��;�=��H�j�1�/x����<����z\�<�f��"�=>��4�q��7	c�dK>�:��I'��Q��e3�^��i���ں�I��R�=3�7�h�h� k>D��=
,1�lg=A�=�q<l}�=F}#��)�=���9�=9ӽ��O>z�����U=��뽶"+��NK������|�=`�h<rԉ=��	<�p=�m��7��@�>���Υ�v��y��=��g=� �~��^T=P�'�E�軝}���0�=�~	��>�=�U�.�=_��m>e�A�dս�h��R>�-<�l���	��v>	�N=-�!=LR)�d�ʸ4��=갴=~����z��=�ER<�C�<�:=*`�=���=��h����2�ͼ';=)<�}e���}���#>��V���2/ǽ��>L�.>��=`��<�)R=�8� 1�>^K����<?O����>Zb��;>$=��=�F�^Q=:��=��C�==:�=���=��x��B�<<�!>>��1}�=�C�=�� ����=w�=g�p�#B=�I����ӻ�}T>�;=����;�+��#���e=��_�nZ�;͉'=� ��F���3>u�����=q*E:�´\��<�u�<K�+���&��<�1��3�%>�1�=2���Pύ=q��=�"��N����{=^[F<���<�I��w���,>,E>܍��h�I�p������="!>v7u�����=&�(>�f������@X=�@8>�R�<Yཅ�f�W��=C�!��[�<
7=ό�="�:<Cfμ�����7�/��=S�v"�=�e���=��>2��=�N��+���i���x��@1�<���<:��=Z�>F�=E�н��<����m�<�μ6� ��@�e�|<�@�;�'��5�h��:��<��<�x��������O��g�Uh�=����9>=�}Q���
��w�yڃ����=��<{��<R�=����p-�Y�=�(��~Ο����k���#`�䊴���ƽ����8�<��n��3�<�g伆����켺x�<}Ľ�� =g'-���$��#Ƚ;߃=��=����	_��U�/<�M�����<3����/]���$>a#>��=�o>ڋ}=�!���R�������Q��Q��=�=D
=�nQ��bۼ��ｹ�+Y=�NI��<Z0��`>�f�<#I�|���ӽS<
��=��=�Z��t7�=M�=�=�C�<3{��V�;I:�U4D�W-<�=����ɵ��#�=O�<� �^�{=1�.=������g='W�=����:Y���W�q�˽�Hb=�$|���p�w��M�؅�|�>��8��;���M<Bt3<~�滛i�=��#=�C��on���8�l�p�t�c����=s5�đN��|�v�B�V�=5��j>������\>�JG��X==����C��a�����'����#�=z�=+���e��}��<�翽��/<������歽?R�L���z�T�82>;c꼓1�S8������kY�;uC�9P>[�<Xl�=�?�(��=9N���'=>Rp<�g�9�i<8����ӽ��<�i�b�Y��W�=�D� s�=u)�=ٯ<��<��=�Ж��э<��<<3�潍c�|`�=�=�x꽜��<1b&�+�>����ʧ����=M�!=������X�>�u`�2�7�M^	����^P> <�T�<�0��{!�<Q#$>v��]���n�ܽ�=�9=ڲ>� �lD�=fO���=�;�=*��<ϛ�<���r�=5��=���;�{�<⃚=_3׼��kMٽ���<�@)��-�=�=��j>h*�=@<�7K��<&�=�ߐ�K�=h���0�u( ���⽙ꮽ#�J=	��;����ļ�9>]Iͼ�׍�%��l>�I�L�p�ۊ>�1�;|�мKΧ���=0(7>��`;�o=�4=�-��/���D�ڽ�Uڼ�}���	���_�.�=]�ż���k����=׈!=NU���
���<�!��=����8���2=HM���������
��)�=�3��B�}�Sx������6p�д><C�<u73<��g�d"�<���M�5=���=)[,=
[�;N⽜����?{�_W`�%�Ь�<0\B�u�=p��r�ļ�Z>��=d�ͽjӻ��>��:�x�< ������N��D�;�~d<p3T=�GL���>Z��=^V8�Ty��r����=��Y��t��N�>GJ���'���>��=5�/=66;>�=�?�rg��M�=�ü�~��ýQ��)T=/��n:�=
�Mֽ��=��>X؟�v���я=�� ��=��<�l\���=���<aQ�I�=o>-�M�}5���j�=�}>G��;��~=d�=�n�=����<��TӼ/e�<��0�=�p�=;��x��=!T��3�?�a��=�=Ѿ��{�����=+�X��N��-C˽��>�
�=�b�=*E{��=弟v�=����s>xk�=.��E)	>�[q���E��=v�<�����>1��{nh���u�6 �;I�>��=S@��Ȑ�=�潉�<n�=�q�=Oh����O=���7�=X��3[��� =���z,�Wܝ=K���}��<�=���=�t��ĥ�=���=ce0���ü~��;�� <#��<MiA<�n�+�<�%�=B�<F�<�[�=u����ES>[h��m�uE$>)	��<���pv�O�<�K�<-�<U<���=�I��V*=���;���<���@U��>�#=@�f���9�=�#�#*���2=���r��=�<�0|=[v�=X�&�����_���@�)>��a=O�ż>��=˵̽'n>�} <�Đ�P
7=��b<XꎼU2>�A�=������>1S#>ƞ�$����>����9^C=����w�=3s�/"������v��< 4����h<�HC����<5j��J��H�=�ܽ���=Zu@��=\�=,��=O�e�&>�נ=���=�uA��=|׽&�<��=Y`=Ƭ=��s=���V/���=';�=	�N<>Q<��� �����ż��-=��<ʶ>~��<O������R��=w�M�L�<^X.�ӶL=/��&� C�gT���o����=*����<���<�a�=?tk=�Z�<� =NW��N����s=&&�=���:�t=ݚ̼3)�=�·=��;<�l���&����=��ü�$�=.>�;�8��M�=��=cT=��=r��=��<��<�Zӽg��L^"�!B@=���J[=����w9=L��=2=�=�Cӽ��:=7��=�><�=�-y=tu=�B�}��^�<&.�����=$�Ľ�ώ&�?=�̈́�F�ں�&�?]����9�Ak��������½�t�=�R>�Z<�m=��i�o'K=�$f��7	�J_�=�}�=�������;̩���Vս4�C��봽%��=t��<�s��9�]�O���7��/u��V>�4G���o�u~/�fWȽ�A����<���x���ؽ��=H�����=���hM�=]���e$�q%�=9��<j�=Q��=A �"=�ݩ�M㫼�N=`�e�>�3��=��`�C�J=b`h�or�=��~=�"���zy=Ε�<����!�=`G��p>
D�Vȳ<��ʼ�J��	�<���=er�<U��;���=ᒦ���=.��:�d>x�yH�����7��\X>�����ɘ<��>x2[=^���Uj���)��T��>%��:,��ɗ=[�n�K��=ޜ㽲q�:[����K��gI=�EǽZ� >�Ԛ��=}o���e=+���۸�=iz���g,=D�e==v=zgż��'��������=�_U>�r�����X.>�u-<�?�=+�>u������v��<v~=�;��NeS���Z3���-�=�t�<�0���S=�Yp<<��=�8�eA;��z���=pY�r4ʽ<[�<�Va=��=a� >"H�=w����N=�ල�=1����{��֟�=�7=9b���}r=Q*L<����CL�;�y���M��I�=�	��_���H����={'�b-��b1�<ƽ*��i߽��
>�n�����!=����J^�d_��X1ݽ��c��|�Xb�="�h=X�=���)��=z��=�� ���<�J>��h=<v���_=P|��E>�_>&z�=BUv=�c=��Z�q⛼�=���<:��=�B��s=���=�V�=��ټo�<a,�;����mz9�U$=�Լ=�U�,>������=���=����%�"��Kq���=��==� ������=v�^=��=l�?�M�y����=�LS�t�j;�
&� ����*Mռ��W�M�[=��~��O5'�a2�=ͭ��>�����ϩ='0�������<=`������=����ȵ=A����e=�|�=�ؽv!˽��9�|A��m:��r�5��q�X�B�X�ǽ ����K�����{��;�T>4�<�Cp���r=R�g>
�-��#M�/�L=5C>��=ILc��k,>��ͽ(���Kt=Hz<򤤼�ʷ��됽V0���}=��&�?=1�K��_����R<ʦ���<>���C����^O���7�z�=y���0�=�o9�`��<CL}=�Pu����'R2=&ܴ�*��=�&�Q��<0�9>HL = ���ٮ=ʠt�����j����!�NbF���>��I<$��<+�K=X�P�"�p�6&e>/�<��:U�ýĵ���<��i��������q���d+=Ȥ��W�=��=4�+=�&=B�A>�&�=�	Ѽ�ֽ$E��
# =.������<읽
hƽJ���������= ������/��"�=�:�=��>9�H=()B<���.� ;�b�=�ؚ���ڼ�"˼��㼒�̻� ���#�z�·>H��<����t�<s�t��X7>����U:�Nx>=��=�C^=0"'>L���:j=~M��/�U�����=��=�>ސ�<�*�;[=��ǐ=���x���1rL��-&�*�>wr�<��;Yn@==U�J=ή.�<I�y�k=���6tͻ�� >8�%>4_�� �=@c�<+ޭ�s�;�>�&=1�D=*jf��
>��Ľ��=��_�o24=�C;��">�C->y�0=F�j=���<����'�0�=��üYH�QǺ=�ce=�v��������i�Ξ|���4&'���<gt�=C�=���=�#:��:`{u�i�ν�`�����=�=�=01��*=Xu�;����(=�|�<7,<)�3����=���=D���"��}�t�M
������=��[��<�"�<��*=�ӹ=k�9=��=���<�K�<A\�����?忽��#=-�Ƽ��<��5=�� ���x<�9e>.�=�]>���2�Z��
ܽ���=����J�N�>�T����@���<���TK��1��H��ܲ<���2ci�L�C=֤D��S�=�	ڽhI�Rd>q蓽�۾��s=�	B>����C���=H>�ȵ��ۍ=%1=3�=��<-�6=!奼�pغ��>���=\���T>.�<a?��0�=L���n���R'�\�컿aļj�=��=lK`=~���>��d=u���.���O�=��<��=��l�f�u��r;[����H=d�����=@:]<�������.i=�첼��B�Hx�=�8�$lW�]�l���K=���Px��k�>�3=)�����.="�=P�a<�������5&>
��E(�<T���T�=�=���=�� >V�[�����=h��<�BT�f�M:bL=}<ݼ!s6��j�<�)>zCi��;<�)�=�x=5�h��=�S=���=l��=��~3e�WSܽˮ��󔿽IĞ;f�=�e=�w���=��1���&>w�����g�;�lѽR���d�-<Yy>�{�;`��<�G�<N= c)���r=A�X=������NΒ<BN<
tD�;b�׬�<w�:	�<�˽�D�=x�6=��t�=��=ː�<�����`��t6=��<%�3���S��Oc��	����<��?�L���JU>�⽽A܋��3�<�Ӓ�Sh���^=����h�=��n�<C/>	����=|l��d6��ҝ<�<�=��}�J��<2�u;���=������x=��R��}=r�����<[
<>\��ٜ/>����%��b��=_���""Ž@�>��F�xmW=������Q���g�6ZZ����Y�g��<p���X&=9�=��;KS�=���"@=�N%=ƅ���,�<�H�=��>����<�����T�H5>̤�{=-㕽��Ľ/<5f��0�=j>�= 2ýnx>�q�������¸<l�u��:v=��J=��I�Ѳ5>}퟽A5>#�� fM=+_��<�=���Sݣ=�>b��u,�L4�����#��ą����;\�<��<}Z=�4<��p�h��<l+��a����B�`<��˼��B����:�ܮ׽&��<�^`�!�ȼ��2���#��x�'o��,�=P�M=l�!������x>�0�q��������=�է�BCx�����O�F=�Vz��%C�pV@>��ּ������=W,�$5������=�B�<f�>ߖ@>��ۼ,���v�����:�k=�ѻ�rR��>t�G��_�������u*=@��Nn<WO�;�#>�u�=Y��<��=���޴>m���>��=����?џ�}�輄P���=tU=��=������_��Mi��oѽF]��ϖ��n����d=^����=��q:���HL���ݽG�<�>>$�;,�S�2o�=x,>�!��$=/���=���=ᕶ=�;�<��ۼ��ڽ�Ӱ:Hm<F�w=���=H�;�_�=h Z�?��:�ڄ��������<Xs�rp�==�/=�	\�Z�2�鳶:~\=XLν��x�]h!�f�>�����dr�GVO�*p=�ֱ��NQ��V��T=�~����_�O�V=�/+�F�W�$�����!���p70<��<���<N->��'=*��Q �����Vސ��;��m�;��=�;d�ul�:%a�$K��Oo���p��Յ��ځ=�彭����7���5�}��C�D=��F=D
��@��=����ڽ�.�=1c�<ӻ=dܬ��*����=u6>���<y<�MJ�q�=̫H�-Tܼ+�L�����`=>��mH =�ћ�°��to<�u�=�Z���S='��;g��<�D�=�4=�&=Ni=����Y$��J>@�)=�+> �L=�g�9��<��<ТŽ��/=�">�X��!;=��ս��=r���׽�ۘ>��r=���=�Jż �M=qj߻�=urc=������=�����"��A-�+z�	pͽՈ���s�=����q���l�<>���������dR��u$��>�V=��=z�`�E=�6��ߖ�<���=�֣��B>�$�=�y!=���9.���V<�l��@;�eͽ��l=����I>����=@�=�>=������< \�i�����%n̽U䐽@���白6�=��<#�(���=<-9]=v}�=��X�=X��=��L=�/$=t������<��=gJ4<�->�3��b<<�<��軄�=@ 0=����]���>U�=4h�<�7�=&�)=l�=�6�>G��Z�<��g�p�+�8�&��+ɻҭ��y{+�QWH��
��]�=}�=��ܽT��C�z�ˁ���i�<Ʋ(���=��$=4���
S=��<�>>�#����Q<�;J�I��F�>�z==�N���D��~>�Բ��i(=O��=2F�=1U=P�h��2=eg"��,�;��*>	n9���[���t������'�=v<�v+>窩��h������:u�C�\�.<�=�/�<�j���3��?�=��ֻ�u�<V=��>��=�tu=j
W�/�v=�C�*��:�Լ�[ =z�F=E�����=����7p��C�2��ˡ׼����^���!:�!ý�Ϧ;R�=�t��`��=�e�;���;V	���<f_������S��JR<�	Yx=���=q��,�=���=�J�8΅���=��A="x>�� >�Z��:=������7D=i����<C� =�m�=�z>���<�,(��P�<@����s�U��=�g�<"��=˔�G�޽1�����,Q<c�<��M>-�v�?m?�ˏ��q�=¢�½�������=ܽ�=q�<�a+�����6 =��<�r=�ǽ?�=9Z/���q�?>-�b=�M=����Z�����=S1��ͺ=O��%�<�r/�X=��U��@�<
]��Ŋ=��<\�;H?=�}��/���=�:8��-r��f�<,��lI��8��U~�=c�ҽ���=�!:=�u��޼���=eTl�g��&�KJB���U=r ���>�@�<ib���=���"��=~=1ʽl���8'���4��v�v=_��<���0��;�t����=�w�yd�<q����3=�H�<���<Ȣ˻� d;9>�=g��i*��C���q`=�h�=S�]�O*�=�
��]H=��=H��?yT>C���ܷϼP��=�Ԗ�P��:>��'� ���=�7&�մ=����怽����`@�j:+=��ƻ�ƾ��=	%�=�Q�;Ժ���d�Б=������[�<�X�=�k�=6ݜ�"��;4-3=j">�����G��=y\;��+<3�>�нo =f����B��a����.=��|����=��;j+�=\:�=�m�<��^�g�s=Qض=e=�Gv�h�T=(g2��Ȍ�sR}=N��<!�$t���=�6�=�z	>lS*���J���7�[�=zo��.�=T�<�|��=�H���=9��r�7=_���J�c<L��@���<9=�5{==6�x�<�b�<�����>�Z܆=��=�h����=C��=�&�	ˉ�5?�>�<��˼B�l=����"=Z:�v�<$����N�Sc<mJ�=�>&ؔ<�$:BK��B\���6=i�½���_>�<�`����#�� >M�
�b}�=���<X�<��=G��<�%�=�K�<�<e�Ԏy��+F=܋�=�/����Xp�5Ţ���K�M�m<nSh=�h��4����>yظ:N[[�Ï����j��/�=of�<o�=�c�K��|\Ƚ1�;W�;c��=�*�=��s��<�^<�i�e�=���<�����νZs�=<�'�I�
=�������=J�>L����S��z$=\�=e�'�OlC�,KQ=�&��ִ�h�>�����,����=�6>��=NՌ=��+>��@>�=r�a��=��4=�8��Q��$ey���S��j�����ʡ�D�;N=g�8��n����=I�d�8"��V<­������zz�<nG�Q?��-�?�!�E|�=�z�6�=0?��'��f���BĽ	>��+=B��=�����ē�~~�=�z�=w@5���=��u�Z�=g�=(fF��n
�ͽ����L^�Y��<�`|�'|F<b|��$P�:�T�?����< 5�F�˽z�:d���.��E��=��ѽk�ƽ�K�5�	>`8j�	/���@��oA�8��W�=] �=?ɏ��0J��B�%z�ݷ�=�_��w�<��L<���c5��l�Q��@4��bG�zN�=���=W�>Q�+<���=�ϽplX=>��CJR={W�<&�ֽ|�����J=ޝR<u�B=CU">�'�=��=�gV��TI<�ͽUj�����=;�����=��=����?�=FW"�Cu�����Bܦ<��;o��<���=n�м�U�<�n�� �<��u��!+>	��G��<���akm:�_s;+G��[)��L����=��<)^�;��=�����<j��=�w=I#μ/W�:r�,�v`�����<V���W��ꥠ9p��<p�y�ނ����9==u�*R>Rz��nt�<8�2=���=��'����=��*�Ȍ����d=C"3�J�'����H�<�[ǽ���=�Ԗ=��=La�x��=�>75������"�=�S�<�w��3E�����;�0>��>͆�ݼͼ좨�����eD�­���꼍`�:?���=n�̺��=��=�D0>0�B=(�=[^%=�z?�����H��>���:ݣ<�ܔ=�V���GH���'�W�?���]�	�z��m��¡����;��=�1��tO�<x��=߸I<��=��S�=��=G>�ލ=u/��M�;t�c=�8�=X�X<05���ڽ3�<G�A���=�6�=�h=~��<�6=���=�=&=iS��;e���Y�=��Z=�I,>��w=� ���<�\@��`�=+	=���Ի=��=[8=��=i���	��}|6=�W=�v�����=PG>M44�MȽm��=�_F�|���V�2��O���;�J��a�;m|[=m�F��퉽54+>$0�=�i�<��"����=�>�ၞ=�	�G%<��>+�x=hhK�``=C���,�=�*������բ�W􏾁^A��ꥼ�s��`Q=dN�=߿f=��M�B�9�>�3�9ڐ����=Ƀ�(�6>�<��X���2~=U:��:�r�V�x����o��y�;���Y~��ݥ@=:��f�=��=Y��<��N>�䦽/��<Z+�<���=;��=���]�<!Q>T���0ŽE�E��z
����=t?�<gH>��*���,�\#��Y9ٽfo�|8����3����F?���=���=���<O3D>i>��a>�p=�x��!g�<K�A�[�T�Ԭ=�"̼�н-�����j=&�ֽ���=U^�<D�<O�Qɳ=�蠼��-�S���)9<&(�9ۣZ��0�PN!<��v=��"�:�+<+��<2�<�Z���̴<����Y���=#�=4,罼���g�=�>/=U�p<`���=0�Ǽ
��<�=�r�=W�<�+�=e��=�K�:%�=9�����<�~��&�<��T��5�;��=���=&�ܽ��l���!=��=R�B����= ����)=�����S���a�<�)��}>�Z�O>Ls��Ӂ<w3�� ƽ�-�<$g����U=�F�9k���J��!��=�%=���;DHʽ��<��=�P�����=N�=�梻���<�Β���h;+`A>�O����t>��<oJp;mν��,b�:��⽾�<_'=e�9=�j�<��=�����,=�*>�8=����%1����;p�>��=-AA�, ����N���=��=p=��ս�==��
�媐;�!���2=_��M<>����R�A=Lg ���#��Ί<E���ӫ�`j�������(��Ѹ<���=c(�=�f;	���=X%r���*�~<���q���jƽ\�!>C���߬p=��½���;`?%=��=�J�����=��E����=Շ$>~����e=L�V��ཙJ= :����"=�&�=�o(���=�$���ؼE��=��=���=��'�!��=&�.��7�:)&ƽ��$>��c<˨=����)�8�6'������ѽG��4�=�+�=�y:�ɕq�z⍾���;F��W�<�,��`�z=�^,>�Ī��d�=�ֲ=��h��*!=�OV=�C���<��';ܹ<2~ú��d���C=	d����{=a�<�}P��I+<�">��=���=AO<T�4=�+��,+a��� �8�=ͼ���[�Q=&�0�k���`�7�<1�=��@��ڹ�8�=��5��W�FE<!Q�hJq;��>f(������-~=��=?�~�5d�;W+���R�������=[x��5d{<�\<���;+Rμ�-=��	�O!=����uI�<�|�b��=��<��C��\=$UB<j��=@��=Y�@�=/���� ��f���)���$>zWg�i�*=!冽1�=��>Ca�=�=�x�<viG��追�m����>��<[����=�d���<<���s�B��m=Kq���p=�U��d�>|����3��#Ͻ^�t��	�<[P�<�>���V�<g�Ի�*< O�=��I��#�<ҨJ=��>�.!�g�r�ӓ�=���;e�J<��=�O���P8>����jzJ��3���]�=�e<N�z���=�P>I
g=<�i=�'��שF��
��v��%nN�dƅ<��l�eY��%�>�ō��F	>���=��=��B�RN����x=ՉU�}>;����!m�0ǎ=ͱ<�IQ=�[�F��=�,߼��_���T=ޭ�<�]5���G<`�{=�ܒ<te?=����a:=�GF����=ܰ�=�[���o��4�=B�_N4�:ȇ���a�3���[����=e�b<*�1<���=��y���=k�����<��<�����b���]<�+=Ҫp�B�ƽָ�`<���>J�;���=��=LQ�<�C���%g�1=��	=+8�=�<���=�����y��wZ�f��ĸ����\�Ȳ������p�:��<���=5车w��ZȻ��R<%/=0te>1)>l/�/�`�#s=ӻ=a��<v��Q�;/<��@<��Խ�[�ԇ�=���=S2�;�#g�z&�L��=��=��=�]v������6t*=O�=P������A2�=E�=Rb=�5�=n=�:�j�=E�B����l��<��ͼ�{4=���=5x�=�<B[�=X������#�սԋ<���=�7˽M]�;��<2��๽ 9_>�3�m�1'�j?�<C�����=aIZ��-�=b��k=w�ڼ7X���W�<�|o=�R=��=4�=`�=��=��X���<>�2�=�_ý���afW�7����u�:wӒ<ECu=
�>WɊ=C5�ls�=~�=<P�<�S�=y��<f�<�H�<L�o=M�8=�J�b��=�1����=�N=o+�=?B<=�#n����<���6�=t��;]˽�f�=FNz<a�+���5��~"=t�	=:�_=�Ž�h;F՝��Yo���<�s�=k�=mN�=fO�<(���?����ͼLW����5>%������Z�>-����;޳B;�E�=y۟�~=��#�z��=xn�ଡ଼=�Y��2Tν���;��׽�aE�h��&����5���>���=ym�=�1�=��D���=Sl3<���<��=��o�7�=T��=v��=Y��;�:�=����ｻ���,vq=��
�?C=�:��c�>�^�=2�3���=�7���*>�C>�h�=C�=I��=M�Խ�6�=;�V���~��<�i=��Zi��� >fn�;�W�<���= F>__�)q5�>�<��/G1>�ѽ7X)���;�3A����=�N=&A=�>�=�����<�,�¬�<�U����J_Q>�]=�M
���޽a ���	��K=�=,�=5,:�?�9>L�S=�m�=Q�w��X�<��2>�<�����I�:tN=l>��A;��$<v�r�`?�=���=n���V@�=�������g��=JV+>!��MЕ��X����b">���k��Cy=a�Y=�/�=��'��%���<��<$���l�=�/�ڨ�:����G��pp�ժ���F�1�W�^F�<�NW� ��=-�P<7��;$qr<)@�=��D�<����O�<��=vg�z�>��5���(�N:;=
��\�=�E@���T�������<+��=����a>�=�E�_=o��NGh>���<�%��>6l�+�=UL�=��ѽ��\�]x�<ta>I��;A�>��Fd�=)��<�@>K�m���i=�6��Y5l;X0=�=�=�!�=f�X��="M�=O@�ó��T�>�_Iʽ��5=}�Z=���=|�G;�ݦ=������<��=�La��Գ����=(�罇<<܏�=ֻ���>���>/>>�5<�A���E�x'�<u,S>�f <"��J�3>��e��\��Ts���4>��=�M,�Ƴ�A�=K/�<��5�&��ĈĽ���=�=	��Z=*�3���>A�Լfܤ�Y�����GT��<���=�=1>;�y�a���=W����J���=��̼���<��m�<��>f����=r��4
=�b�c݈>Zi����V�������ý�hZ�ҡ�<F�=/NA�}�=�`+<8��=|@Ž��%�j��=�!=T>ʽP�9=��=�*�}6���Av<,
�5�����<������<g�=d�{:�����P��«�n�7=h��:�<��޽w�!��T�#. =�����)~��u�;(���2;����+��=f'�;���u�D<2{�<��Y={�?=~�U=���<Z���;hY�8�h�1���j=�=��<�P�=�oB�<����<�9�
�<;'�6ݲ<��|���������
�=/v"�?lH����<	TE�����e<$ʺ�DB���6�=�'�,J��-s�g��ֽ��Ž�35>4[@�z;���#���8=)2>��M��2Q�ds��t���n½q��=�Ԉ;�Q?=���ܪ�����=k����m<^�4��=�=J�5�K���
>Gj�=^�W�=�r�*�6��Y��D����h��c�=%R*���0>�Rl=`A�<X8�=�9�=��Z=?�=���dK=�V
��99��(%���n��`��%�������T�=ކ��k�=%�>��=	�<gH;����Dt�=����w
6�P�j�R	&=]R�=�ؼ�	=a�O;�mѽxyܽՔ)=� �=ν�W�<��l<���h*-<���=Kj�[�p=$�)�熪�R��=I�E=�`��_h��8����< �Y=�����{=[�>�1��<I�=�#＃靽:2"���ҳ<�ٽt	<E��3!��0o��л@{=��ʽ��Ľ�{=Nǽ�V�����u=��=I�ֽd�ҽ��=-�2�	ʒ=�=��L��<Z�O����=�n�aҚ='�>.�+>��ԽfC2���;���^Xs=��=.��:>aU>���=)@=�w���<<�ȽX+��|�vv��;�|O<&���{>��������d�,�p�j�=/J�;&��=��>��[=g�s�I-=�=�.J��k=�D$��֥=��T=�/=�
�_1��e����y�\᥺�*�=#�7=Dh >"	Z��9t=V�V�-����B=WA >{ȴ=O�>��2�'�,��|>�=N���<�k���'�� '=����ߛ�=��=��+��޽�<�/r��k+=bma=�5�<�D=lا�YĚ<@d�=��}=�bL::�
>���=k�< 
�=nU�m!<Jv�<r�?��t�<!�6�s뼿R��J���v=������Y=�]��=9>:�O�a��=}�*=�)�=~�>}���&ݽ(�+>A>G]>6�&=<��-�`=��/��Q��6>�T">��=1P�;U�~=qr�<��=��:��e>�b�=�V���5��^�=І��f��=�%"�L!<S��='�>҈c�,���2=�G ���:L&M������-~=^���R �^4>���=����B�7�.�h;F=$���m�=�혽k�������������*���.=I�w=��<ڤw="E3�;����=;�U�|O�;7,!=�w ����<��:�������>i��s���ֽ�<g=����+
���;��h��jt=^��.��<*�="s��}U�=�t�<���"�FQ=�n�=R�>�Ҩ����*=.�}��n	>l���mlz����=Gkv=F����O��0�Ƚ�ݨ��:>m���Z�=Y�#��l�"i۽f��+w�=�8��&�ؽV�=�Ȑ��i=���=(����Ǉ��H>��=9�<��=
M=�'#� �=CW<��q�L�������<>Z�=y<�6�����=�z�2S����p�=��;�
�]}���(�='鴽���=��N�����	1=�*�J�;=&�=wx�����=��;� �������=jFa<���ܰ=g.3��F�����ƻ����Q��;2Њ=�^;>�BE�`Dֻ��.�j<a�̽����{���[=�ٽy�'�̞L=�,y=:�=�1�|�=�F̽�Ҥ;{�O=;4m��%=��U��ƽì�=?dR=���=��S��=_?��V�=0V=q�=�$�=�W�9RH�=�i�=y"=�����\ۼ#���>�!=E=8=12���S=R������۱;D�=ai���=&�F%�<.���bB�����"��=��ҽ8o@<�j=��j�J�v=����<v/-=jb�;~RA>)]��#����=e����6<R#ǽ=���e��=�[���M>�.�D�=��=!D�=s�>�q1����=�� �^=ʣ�<��˽�-�=i�>�7�;���<���<P��=� ɽ�t=��"�0�G� >�<1��=�v=����j��;�=
c=�W=������]��=께=�*��;�Q�ۘ��7��<�+(>�� ����=Id9>�Pļ��a=y���BJ=�J��j%7=~4(>�a{�S��� !-��bg��@�=���=��<�ny<ҩ�<��:�#%>1�ڼ�/v=B��=7�r=2�����=_=j�L��� �ڞK��<�<-�'��=��>=w�=:^P�@�<=1��'T����X;�!"���4�&ix=x�=q�%��"	>�\����>
(�y�2<=��A'̽�Qu=�^�������=y��\>Ü�z��$A=���;��&<.i<���>Ϝ%>L*н�q�=�駽)��<G���漼��=�j\=��;=� �ڧ�=mnl=vL��	<=@K=�܀=��������L,��.�bU����<�㯽�`�v�Ž4�={P���Yɰ=w�;�΂��Q�O�Q=v��<4Kż�T�=�S½k��;T�=m+��--�0��<�k�<��=QK�0Uɽ`�>س�:�%�x��=)��;�rl�Q��=��ǽ�<k"�ǀ3��=���½�2�KY=2]���G�ý2r<��=�S��6<����1=Xz�����;��F;oC{;���=坽Y��<h�<��)=���=x۽�͠�=��/�<*�W�
�=�e�=�݌�s]�=-�o���ּջ�<# �<�1!��J�)�=���V���f�O��VL���6�<�3�;7�������W4��9��0��e;ΩٽJ>�$��&�n������S����x��<��=j6��9²=��@��.�=N��<�7�I�a=�R<>2>;��<[m3=��A=iV�<n�#�G�����q�ё�=�AS;P���%��	��<^{��צ�����(���@W=�%�=#μp��;�~m�@Ӽ��
�@��=��=FP@=��Q>>�h���=o�=��>�ڙ<j6f��<�.��=�*����O�;���<hd�<�+�:lC��2�� 3=����Խ��¼1��KI=f-2=El�=�rһ��)�fu��T"�����=�sT��;�<��>UP�;��U�Q��_U=
+)=o9=�B�������&�s�s�h=3D�<����n�M������[�����=)��}�M=�籽_V`=��*=���=RǕ�˰�=ړh���{�=̼<���A��,!�����E=*܏�if+���<h��=z�<�Dҽ�*{��tS�����=�G�=7h�t�>4p�<Zȥ�@�r�f錽ۂ;[L8=�R�}s�=\7-=5=���Lp�=*��<	Y
>r#�<߫!=g;M<I䠽�W:>�̼z�^=Z�+=��=9X�=�vӼ36>R'��aܽW����M�=b[�<	\�=�c1��k�Ŭ+��CM��R!>11$>��<�h�XL=F�=�r�=O��=�K��o=A6 >=L�=�� <ƙ���=�ɯ=�ߊ=���=M��=6�x�����ֽ1��=�l<>{(����>�oG6�?�7=�0�<?P?=�9>TH�=�>�$̃�Z�Z=�S �5c>��=�p<�P�<^-�=dLϽ��O=4�⽑,>�;���d�Ε�=?�;­�=k�>x�R>tE��Ϗ���=���;-=M�a;��<�P�=t2��V�<Ԣ�<���=Y�T=�娽/s�>�><m+>p̽����$��=�wf<f�ǼCF>�gY>��r=�)(��ߓ<�����=�W���y=R�r<3:�;=~��WW=X�C=x��<��=�D����;<M�=,ι�7A�<B���<Z��;�a?�$��=�xQ=���=�[��l�=1�ż�"�;S!����=�e����<�	=��[�����S���_�=�4�\�6�5z=ܟ���=v��9��)��ӽ`i��p�CC�8����q>U`�=���=�6���`�*�b�@ऽ��_���f=}=�=���=7	��Mc=U�.>zݭ=�t=��༼��q�0>��=�#=� �ǹ��AM:��1�	>���rT
��7>�,����R��Lq��0>�D�gm�� >���=�5=<�^�>./i>+�=J�����b>�_̼�n�<RM~�X`��|���HG <���>yP=(l�<���=��
�h>���=��̼�]$�W�r<@K�=�O��[=�,�u�������w>w<Z�,=72��=sR�< ��M�3��i��<p>��X�\�;�W��_���G=Q�=6-�,!��8�F�A(�e��y�-��.K=@gZ�Y�Y�!�<9�M=#[�
5�%
��br<y<�{\׼
���%y=�7=;��?�<nA���g�;,u�����u~����N�*6|�DDS�w��=5X�=�ɻ�>�=�["<:�=���=�	>�D>Ɲ��d��u�<��=��>b�^���I=�v��n�;]�=�Y��5��I���Jm=��b=��*�������K�''�iz��d\��W=�ܽ�p�=��/;��=�7	��S6��5�v����<<����C�=�3
>���Ma6�5<���<D�<��	��h���8��<oz;�Y��t㽯����ȁ���7=�^r=\��=h]��CRE=��=ڍ=�C�B�"��3=n�;_�=N 	�ƌ�<����w��=�,�<!і<�B[�Dm=�㟽 x:��OI�N�M<͢�<��={�ɼw[���``���x�'de��V�{�#>9"��F2/<���� =���[=^>��ýY���ie=��:���;�>�ڣ��ʼ7��Nz��ڽv��=�~[���z=���~��=��c<��(>%>�Պ><����=Xb��F�=pn=�b�� d���&>��<�:��:�m`���e޽\�>�<���%=6�<�Hٽ��M�<#�W$½��=��=f!̽*��<���<��2��<Y:�x�=�%H�fA�2�%<.Ic���#=� ���ɤ�5��= ����B>�q�=�!>=����@p��5-��|˻�$ּ���=�p���zZ�*��=ut�<�ӈ;66I�zǖ=�C�=@�<W\&=����ȓ<�=5��=��Ѽj� ��ɺ� ^��0�<n﫼x��;¶�=t)>�}�g�9��2B�4�ڽD:�=A8D��F��Ŀ=���[f<;�'���{�倸<3�4��q�<�hr��i�����=�Q�hcٽ�m�3�н�PC<�E�=��� 5�<&<t�=+�>��7��=j6�y-����=���R#����=�����_�=����9<��e���.6>R�=��=����Gk���p޻_+]��ڂ9V�.<��ؽ���<|(����=M-=�M,�����y�<�Z:=��:����Q�S<Bd�����=�g
=e��=����ڻ�?�|�X<��C�<�߉<�e��=g�B=*�� ��<���=�Z=�i�=�._='i�9l�=$�½����$=*��:�+�>KWR=��g���<����ý#��=c=�UP<���|�����=�zH��;N�=`j�=*�=�<�R���"��ơ6=X�<�������=9N<Y��<*b�<��Z��<�r>I`F��p*=�޽t�Z=�v�=zkj=�������]�@;i����)=y��=?ⶽ+�2=�a;�:����=�A�=��{<�g=ԞP<��<K��=�r=J�<Zt.�	����Xν?G%�x.���ǟ;dx�=A�2��ż�1��l�=j͑=��;ȪV�h�=���=ê�=d#�=`���d�=/ܐ��S������������=�~��|f�}����Z����4�Z�X����>!`����4>�0�����<
cG�k�#���>���<��5=�i=�n�&�=����E=j�=��z=C���l�;�<�@�<|�d=$|޽���=K9�=(���$�e����}��x7��q=� +����;�1��u���OK�A J��q����)=�=$=<���2��5��=wP�=�_ּ�V������>�_�<��<����K�ƙ@�K�{�\���d�=*�i=�T�~?ҽO���Υ��7����������=VI���q�Sj>����(ȵ<������r�=�,�<p���­�/o,=Y]�<���� &>�%=®p��Ӌ�7/�=4�>bu!�12G=}F���3>�Ǽ�!�O1�=��=Gm�����=��!=u�<����D"�=ʯŽ�bE�>�<z��)=)���%Sk��=���B��F��<��ڽ���� �0X>�%X�V%,>���<k]3���f<";��<M(�<t[�����=����7���d=����}�w=�=�B�=gz=��;F�2	�<�(T�Q �=@�-<�Ń���>�T���̼=�=[/�;O79�#��:x���=s��=�����t�<#߻��h;��\=x��=4� >0mL=$�x=7�<gЀ�Yu������c�����?v��XH�l�K=��-��=�=�^�<(��:P���b"�;��1�����put=�ǽ�{=�8�W�=���4���=F�.> ��=���FO���ֽ���=��;�ͽZ�ѳ�;��=��=vM=⨹����=h#>q��>6��=Wt�<ϥP�� ��,�������H����=�X6��E� =���p�=g����	>�l��`������<-��=R�)�=_q=����{�������.�B[��!_U����rE�=�)ʽ�K7��e	=ç >�z�<�>[5>��?=��|����=��n=���=>�q"�=�3<4nY��>������=w�='��=/(��mev�{ʽJR�����tC<��^<;�<�4���`��섽�Y��W�=�v,��=�=}��:@/�E�����=hx���k཈��=.�=����-{��,B=�)�=?��<;��{4���=߼W=3r-�m�=.�X=��!<�&>z{=;�<�r(��>����e����3=�]>"�=rPֻ�pڽ��*�h�G=v��=+�*���A=b��=x��lD`�>�=�S	��t�=����<�=��}=��v=�B@��Q&�=/��oc�Mk������)�
�sr�=��<�!��Γ`=�S<�����;�f��V��<��>���=f9<��#�*�(={Qk=y`4=@���ڶ=3����5�8><&<�M�����Γw�p	>�
���d�k�p�����	�V�>��N/=P���<�l'=��~������9�=��=��<�Ȅ<��_=-N
��=���"�=˗:3�<��d�Eh���J>���$=ӯ������q.�@3���ş�\�1����c�;=�b�$Y[<E%=o����6��N�
<L�<>������3�a8=�����=>�[�4��=�Ly��g��A��� �=��U�؀�=��< �ٽ��b�<�*<��%>��D>��<�>�=�z\:%}R����[ޅ=C�{��'�=:���9�=��&��޽�����=��<�z�%*�X}�<!�=p H�zf�;�,r=��a�����*䷽%T��4½����V��=��2� =� 2��!�=o~P;�
&���0����<d�}�>�4�<�<OO<HK�=�H׽;R���s?=�v=��=��a=ҩ4<�r=��_��(=���/w�/�<��=�*��P����V=�=��_�<�[<�㦽�]q����>�.Y����=�9=���=�iN��˂<���M;D�4�����<6�����;,C=n<�Uqb<��R��ܽ�\�=R>4���>�ֽX��<��������񭽖�>)ƥ=N�\=-�����<� �͎w=~z�z̽�����>|��=�$���@�=Nx׼{�<�ý�!���<!�݈(>�1=h�>K��Q���_��Z=��������ܕ=|*��ˇ= ����'�6>�l=��>�A=ݏ �bm��F���Qi�ע;�� Q%<cۨ=����H>h*!���=�H>TY���)'�@�>x�g<᯸�6B*������C��U𽾷�=�p=��ͼ������=��I��Ч�[�!��'+=�(�=�.�=k
�=N�*;�6��蹽��=� R��ﳼ���sb�Nz��S�5>��<��7&5=!��<B|��4��cr<"��>�<֚j=�=�=qA=��j��E,=���8{��<�2���=i�|=; ��T�\=��;#A�=ֆ�=��==��� �<�9���=�3�5����I˽�<���<+Խ�*
�D��؟�;�����^<D[���¼�T�=
G�=<#�_X��u���� >�O����������xʏ=�=�Ⱦ<i�@�҈v��Ę=�->l0�;"SC<�@�=�=>��p�5Y�=,4ҽ8��>�<�fQ�����.�<�^�=�d=r�>��=s��=�+��!^�=�������m�<���=�sH<�4����=���=��b��+�=�U뙽/��ms�=~I2=�g �!b<��<��<��h��� =+ZZ=*�f�DԄ��u<�SB<r�½R�>�w�<$q����rb#>+L�]���ᇽ���<!Q�=+����N=�ɼ_�0�sJ>�=yV >�h�g�u=�J��/�8=kP�= A�<\����i=�90>ׯ�TVڽe�Ƚ5��=�a>���:�n�=KW�
w�<��>�=�)=���=�eټι��:�;>��=q�9oK1��̸= ���D�8^1�{7������`_>��m���"�
��e�+=ꖵ���=��&>hǼ}�ϼ�|��h�n��k>=a�<S�<�.ż�l!�Ev>��<k�=f���Y����>�'i��'���s�;��?�f];f6Ƚ��u=���-Ȧ<s�Ľ�5P<���<����)Ƚ<?t=}�=4�ܽGx�Hv��� �=�4�=�?���W�=Q'�B��<�Q>_F��Z�=��g���8=���=�� =��=���*���=�=A=�tZ��v>�8Ľ�᧽ê��� �=#d�<G�w=o�<>��A>��{<���=c�=���=F/����<!������:P?�=��ֽx�>��O��۽u��_!h;�|��@��"=�}�=Gb�=O�	�;����ѐ���(������<��x�mW�=�%(����=#;����f��<���=���_��=�s����=�.ؼ]�=N��=ZU�<D�=	"���=�һ���Խ78>����i�<����Ƚ=?!=��\�<�=� Ľ">�oJ=�K��JúG/��(�
���>ۋ=O&<t�9���D�d=�;=��=b#��S<�����M���=��Z<؆��
�����=.u'�&�T<؄�7�뼁�ν���=]�-�f�=�4н����IG����
��O������^�=�,$�� =��>�Y3�8&۽� �;Zy�='��=v�^<��%�����͏>���<:�=��U�=2��=�	���,��i&�g�D>�5����N���m��=�ڽ�հ�ϥ�*�i=���S�">I�;>]���%ͽ�s�/`<�|�=F7�=S�ֻL�����Ի�$r<\g�r�t�ަɽdK_���=�F,=YR>�^�=wy~��;�<&�S�C��Ĳd=�y�=;k�=fm�=陭=�O�����<��=��
�{�=�]����q��d=x>����l>U=b��<�u>lQ@�vخ<Q��"<����M�=0�<J�=`]��.{N=ev
��y���=!
�<�=��A��$���>�wo=B��=�譽�a��ܚ ���.���=��e�NZҽȞ�<��]N���<�=�&�51T=zp&��;t����`���פ�.������v���=�Q�;m��=2�}����椼A�0��ˁ<W��<�$����J�N�E>��=�W��(瑽*�w=B���8G=�fT={Q�=�\<�i���� <�,ռ�X[�=P��W����	��Fz��z �O�����x��;�� ?<W��=VӼ�G> ظ=(e$>��$��e|=#������=v��=�u���4>�q�=�M�<�!��V�żM�%=h�;0mS=/�f���=)��=��u�~�\>��==ԟ��۾={��<��*�m��X��=	�'>?�=���;��Ƽ\��<T���TJ�]�=�K�<����*��p���ý�ּ4hI�&��=報<� "=)⟽9F���p�=��v<�f]���t� ����=�X�j�;-e����8M��ц�=�$>L�=����=��/�e@H=��f= �ʼ𶬼�Ҁ<a�޼O�=��A<;��=7c&>m�,�\�=��=�z(>� ,=�Mǽ�>��><Ch��*ɻ�q˽Np���+f>ç=���<(��=����1=:�>=�a���T[=q_��t=\R9�7<�(❽�V��GE��Y:n� ���
��=;�����8��ԍ�,�6=�=H_�=��=(�=�]�E򴼁go<�+>դ@�./�=�$�<�8�.�<hW�<}�$:�k��'>(Y=�6ػZ/��(�t=0��<0s�=
���<�
���-�4����X=Bv�<�#Z�5?�f�L=d���֔=/]4>W����=���ˆ��5�KNA�nL�=}H��C*�������R��=�W�<}6>��<��ͼN�>�n�<1��X�+��ό��=�^l<�����=��$=ɒ�j��:��/=#ᏼ\^�=q�=��<9ý�;F=43={�;�g~��>t��ҧ�=)��4+��r�=�K���Wu�6����h2���,��n��_g�(�%�Ymu=N-ý�P�������� �@��X��<�Ԗ�����ǡ=��=!KG�Q�=>��=�#<&����`��\�<���:�X�=�C>m.�g��=g0t��Y�:_�-�Ӿ�={��=�c�=�ܼ�>jH��o�=�m�<��=������=�R�=2�G���]�i����v>��">����=�3��=<fJ��=`Oj��F�=�  =�R�=��=�&i<IP�=e�<�Z�=���J�>=��=fDq=�~���)��=qK[���
>���="��U��=�|��
��狽7�*�E���B
%=h}�;AL��=����0A=����U<���V�;��=ي�<&7�<xo�<�5�=����ˀ�Ms�=�</^�=�j�(�=�S=)l�=Yu�<Nw�=�`%����=^��;OȽ���=������=�va�Pv�*;�t�!���/���<�ej�{H.<�}=w7�����G�=�i��=T�R�����K(�����@�<�<bSx�Նټ���B$>�\>4:���Z=%ݟ�<&����Խ�g>��>]+>y���B�=�O3����ؿ<���:�rn=�l�|C�'��=�ü�%��aȻ�;��X�����K��{C�; �=� F�n�ϼ{�S����n�XZ�=u7=eK��V >�磽�>v=w.K��U�< 5����<tr�<K�y=�4[<� ���<kв���};�&7=V�q�9���2��嶽c�������3=�
`<���<��ʻ�)�+��<>zݽ�^=����=�
`>�o�=�b\<�|��H�=�����<7�?��r�J�=[9;���G=�F�hж��v��57�=m��<x|=x�&����;'9���/��t$�������_;����
���e�B��=z)�=�$��K���������b���V����=|!S���<�˽��%���N<�ǽ<��V"=��">u�t<�wd������C�)/=���<pc���V}���3=^����=#ܪ�?i^<�1y=L�I�O�G>,r��.�����\=�A���r{<x���Dg���	�=�2=���<յ�= !�;-=1�k��&����2����=�����4�|=I>f�e�9v����D�F�$>��F�S%j=S�$�(Y=�B>�cK=��,���=���9^���xC>�<�����5�9>�ߪ����4�>�1C<�c��:��=c��=3[�#�=
>�v��<R�=��<W~���뽏�����<_O3=m��2�����]��L�=8��O໨�/�@����0-��+�e9�=��=�Z=q	=-2����> ��B;3����%-�t>Z�T>�.l<ޏf��'�=��0='m���O���]ء��A���[=&�=:`�=#�;�H�<&V�=x�6��߽�9����=8�����dѓ=�n��\Eͼ���<3�:�F����=	��=�Y!��O������<�'�=��׽>�!�II=�1R=�½�<�/�<X��=-_�<,K3��XĽ��T;[�=\S�.ʽJ�轑~ҽ���=���=8�9�ް�=����MU�H��=%⼤KO��=�r�a">cm�=,ݔ�:�ѽ�m����<�55��*��b=��X2�=�8��}y>�D?�><)_� �?�!>���|">�����c=�`�=	�O=�f<B�=Ա���[B=ΐ=dy�=b;%�=�1>h�1��F���=.�<2E��-Bc;��=�T�<Ǽ=ϽսGf���<���=:V߼�o�UX��{��=@b���g�==��4՚���Y��)=k�<�to�iױ�(�:=�"<O��=�c=`���׽����+�<=^J����D>���<��B�cQ�=�H�=ګF=� �<�UR<k�q< ���&H�=l=�~�%(=��=�#�=Eʫ<�C�� �y�>4�=_٦=��=쮵==���I�ҽ�V�pt~=�N�=˵�μ�=��>.9�`�ļ"�-����j�=��	�$��<�">�}z�R�>��>�����-ʻA�=���Zc=Ax�=|t�Q�'>��T<{*��]�ίX>�;<A���~���>-� �=�m�ƽW�;()���댾��2�����z����'��-ս$=~�ý��(����=*���W=u����d�={�"�D=�f�=���>"\v<O��=�]�<R�v= b˼Ԕ�=�!=�ʿ=I���==�'ܼ$J�S���G[A�� >oս��=}�F=Hr(�9�����0A���+���=,�=�;�<�^<�˼��x�
����+ ���h��!�;�rN;�Wu�L��=BO��=_>���=U�������\b�Z����Fr�[̘<i(�<�1J>�,=!}�=�D=dh�=J�(��M�=����<��̽*��ҽ!]p��z���.�<��>�N#;�[���s=&4z=�O�=�g=]Ũ����H��u�z����џ�<(�s=4^y�B�>DC��b����=BX= M��=.=���=e(?=�_	��++��[|����=w�<�*��#��_t�F���w�c����=1	�=�5��ݘ;��=�����{��c=\��2?�<;��K�<B�"��b%�%�=3s<�!�<i�6�vh=��$���A��p��x���ϼ��ѱ=�<=q�;ա;�R�[=�� �]i�<�W=+����<�F���ڶ=���=3pt��ṽ�>½�I�U��<�w=� ��ኽ�#>���z��L���H*����<�>�GT=��<�K=�-�F�e=�3��}�=�}(���D�(;��H���l��=b$�<f�=U@�<o��\�<2��<a���5��[��tf>3�>e�y~����=sl��Խ+�;�l=hZt=sޔ<K"�"��=��
=����_L>�,�=)5z���=���`���.��
�*�Z=��t;Z,G=Q��;���=��Y=�TH��x$=����r�=�̜���>�����<�d(�>����=��_���-���<�q�=�9p��f�=���=8�&��ֹ�X> ��;F���R���3�Ҽ�P��e߾<ܴ�=�,��b=n�i<ߔ�;�=O���+=P��=?��LD��n�<��X</?�GQy��:�<���߯���7<�N=+N��'���+�<Y���8I�<�5ؼV'�m�V<Ϲ]��DZ<�xZ�����zT$=�߲=�<�L>���=���@�{=sw�����<9]�<�8#>!۽�1�<��������녽�N���Q5>��׽�X<=~;k`�<4�8=m�i�iX�=���=_�c����=ӑ�=i�v�錟�&���d��~�#=A��������K<�]9=��b<KY���=ng�cϑ=�T=�fϽ�->�*�<�Fj=�v�=_�~�3��=�T��X���pE�����=���=9h����P�����=,�==����J����<Մ�h;��PU[=~�=�쵽��<�it=V�������}<��M�R�O=UAh=��ν(�=��=Ԫd�_=\�=3準5o=弗���B�֫=<������/M���� =yI�<wp�=������ý�c<��=�B񽊁�=ǟ\=�<|	4��=��:����Ž�ƛ<M' �M��;U��<�
6�r(U=vQY��^��5��T�<U���ٞ=��;I�����=<D>�vY����<�ｷ�*>���V�o��=�'���b��>��I=�;Z=R��w�y�)>=��=�H�'#�=����֔���=��<���=�Ŵ�n� �	�='~8=j��=�l�=����Lޙ<c��C�T<w=���=��>?-��6|��F�_�}<��=�<���굽���/�$�<�@=��ڼ���=5�h=k����I=%��=���Z+�=�h<8o뽍48�
u4>#v���旽���=|#=�y�G<9��:�rO>��e<%e佳���7�<��<��<��=�K��(=��D����V0�=�~>� x=PsP��>H��=�]'=�h���6��i=<�i=�_;�%����>=p�=n��=�_>��u>��!��|f=䮲�3ۘ�(�0�Q��=��ȼ����m��@4�#2���oȽ�̥�����;Ow�Y��f<��=7
B�խ!=�kb=)�����;=A�>)i�<1���	�<�0��Q=�g=����	ڸ=���ڒ�	ýC���0*����)<�5a=��R���<���= �=��;!_B��/>p >tQ�<����_�ɹ<�-���h=G�<v�7�<e�:�p�� ��}]��҆=���;ܫ��_">�W�fZ�<�B=0G⻤~<�����4�b��=�Ec�R=�\�����=xm�v��9=Xե��tk�bE>G|�w��=�)�'�.��f��$�}=���˩J=�tǽ�@>Ep�<޺�=\��Yѽ�Zj=So�_]��G�v6���B=TO=��=�0�=r����;��)��¼�p=6=>K~O=IT-�����:i=�|���?=�Ed�� ���Cֽ�n=�J�;��ɽN+�<'�=��p�� >Qh=6�=W;a>wtj�%d=>>��?���:=�6
�	���)^�=U�i=���=|>�=7SH=L�漁�=2RA�FHϼp�=���;�=q�g�&����Y�=ƙ���~���=�����q������4�=]�漏� �	D,�/�=����v0��k�=�</�'9�;�8��m��8i>����J!��}�>��=��8��<b=�1=��}�*O=�Ƚ?^�=�ܽ�ȽOB�=i�o=p�\>���=9�>�V���%ӽ������=K�8=)Ժ�K.<֞U<ֶ>,B>j��a�>���������0�/�,��d���(�v�����>Phr=�4����=tԘ�L�h����>�<����`< �t�|
��@�@��=~��<�{�fc=���;��Y��mӽJxƽa	F=��<�ې��m߽�-={혽��B=J9>R]�e��=�I=^��}S��T��=��+���=�,Y�B5��$=�>�����p�Խ��p;��;�/z���#�����VuQ�Jrx��o=�:��>���l���觽3kT="�=��=�U�=t�=ǥ�=�\�=FK����_�����J�y�nK5����+ѣ<�z�=T�����L<�n��oy��x�<�P�<����������t��ɭ�߂��{<ߩ���R��H�M<�0�<"��=�!>�<��<�`}>X��e�<�B=<�l��0=���Ke=}��=�q>W�U<�`(� �;X��=��>�T߽�t���D�T2=4�=>�����ŚN����X	�^(�=�J4���<���=U4�W���d�=4"=�3�;N�F>��.=~&d=b� =*t=�	=��;�}���&�<���<oܘ<�Z�����j=Ǽ�;�Nr��S�=�"5<Rj�}��=�`��H�I=;V���y�:9=o^޽="�[%K�%�ɽ'#�<�t=f��<�썽	j��ݽ�C�;�(�ZN�<8�D����<�<E8= *>��w��Q=� =SQ
<dt��+ᇼL��<�ڼ�jM�@����9�<'�mM'> ]�<�L=d����=t�v<�G�ҾQ�U=o8=���<v\>S{�P���!��ܽ�����t=��>�8�=�86�ʠP=	��=���=J�4>�1y=<��;=܀�zW�H,J���N�bZ=ZB�=>/=HGC�)=��D��o�=���k��3� �6\�=�ԙ����;S�=Li�ˏW�QH=N���L=�#�=PJ�(�}=)���g>c�<��"���)�&?���㽀�"�
��'���\�y�����='������� �=�=�)��Q�=:h<v�<��8���=�l=�c�ڇ=E�j=^�ZGR;7}����=���VAQ��s�=��U�iH�8ؖb=�=τ���ν�o=7�$>�=[�2n佁f$�r��=ཪ=Q��=ҕ���0��j%�J|޼�7 ���=1�u�*B <��;�1׽�y��z'=�NR=���o߆=��C<��o�=���^<�54<֝=q�H>�6��숽��r���3���м,>�w佮��ƚ��)��	�=:�X��B4�3��=�EY=�\�<"�=SU�G�=��]�@~=~ʻ�=� �<@�=n�T���L����<��=5g"����= /B>���=�Mi=e�����=yY]��ѻ[d$;�B�=��(����w��=u���z��=ʟ=ص=��<d��=���=��1�ܽ�dE�!�� ;�輣.�Xvu��飽:�S�f�m=ɟ\�;�<��=U7����==�O�D�;�(��?y2�z~�=y�B�{Mؽ���i���o7ȼ���<����_�h@==��5��Y=4����z`�D�B=��>�7<s�=���<�𗼁Ӌ= ���<=�Y�<��Ƽ`�X���+=��S=��\��@>
︖�O=qH�=���=n��<�b��݈<	PŽ��=CM�M4�����<�;��8H���A�1����,=,b�����E>��v=I���f����z=7^�=�)�;ڸ���O4����<١���+=nj|�1���z>� q��8�����ze=5һZ���W	H��|���:�=b`�<�z0��u�;ha�=t��˚#==�<����qD�D6<\.j��aӽ$�R�*y�mle�V���佩� ��޽/����g�f�<�x�=>a�=^/5=d��F��"�L\"��y`<�����U��>=����Dn>�N�W��<�Ϭ��儻y};���<�u�=�[>���<�s�<���нP�R=%������S�?�J�/=� ���	����9�������h���V<P��=�U���ph=�g��f�ee��ۚ=��=�����ٽ����Zxi�ˑ����t<s,8>�=�̓�N!h=vB=g"��%=�`�<���=���Z1�*� �_=#�<X���uw�=N�%�Bn�=��W=��n>Q�=�����;<�s�<���<���=)L�=,�C='��ي=o�Q�&
��������Kͽ�2�=��	�GM;=�i=(-3<ژ���rl=�;d=�n)�mO�=�2�=���<�sZ���������;�d=�a�=jw\=ʛT=�Wü��=�=g��f�2=�m�=ނ��j=������;�=%��=�ˬ�fS �"f`=��]�Ql�Kc=U��;Q�	��&f=�c�;�;�/l���g<h~�щνt������8g��K�=�9�<?�_�Ӟ`�u�����.�"6�=2_��'�����=���<�o���6�)x�� �>��</꠼\^�=*��=��=keb=H'm<o�6<��^� �k<=�<���=����+z�=@��;0kN>�E(��H��ٽ��=s��������۽t֙<a''��(=2͉;�^�<K0�b�輢K����K��Ի�.�=��<�����u�?δ�g��=��>��S�A��*]�C(�;l�=1�,=�I<�{�=����N$=n�\=�ԃ=؏G���(=_���ƽn�<}ч=��+�	��=�/�=���<��R�X�4��� �7E�=�m���(=�P���f��le4���=�ĺ�)�s=��lI>�_
���*=
v�=l#�=���<|�H�����:�<�f�<=�>�I�����[1�=�r�=����$ <��?=+��=Ĝ	=e�=9�U�j����3���A
���=@�W���B�÷j�'��=����G��S �=a�L��5���%���^���V=�`���	>3~�<����X�J*�=y�&���[;%�> ��;I�鼨x=��<�_T�,�~<��`=��"�M<?}=���#F<=��>|��>9��]�=���=��!:�����i=Md�=g<L=ދ�<=�J<��j=��*=��\��݉�g��=F�����>0�=�9�<|>�=�ݐ<���=�@<%�=7=r�=X3��?��ϥ<�MV�M�;���<��;����V���5X�U�M<�ͦ�UtؽA'g=`g����t��2�<���<�a�="��=�ݎ>6�=�"���uu<�J�=km���>�E���8=-:A=���=|���������;Ja�=�)�ҭǽ�e���=��e=�e�=r9>QH=��ʽ��t��u������]��=ȷ۽H�����A��������@�|�������,>2wi&>���j�o>��
�'l�=��L=�s���y�<���Ήr���;�CT>�u�����`�Ŷ���8���-�<�e���a�S����oI<���=�?��KFڻkrC���=Ҕ�Y��=�����i< ���Y��<�Q:�R�:6�<H�!=��ܺ�#���(=�l=[I�=�{��}�>3OĽ�T�=��������bs�=�]��.�>�@a=E�=�y�<�C�<�o��Af��� �B������<��<W��=e�=H>����ὖ^����=R2+;�%��g�:�	{y<_��[b��s��< .潻5��>�jz;��S=��5�!�=&[{<dbԽ��b='=	w|���xq�< �<�{<ܯ�(z> �s=r}{�uQ߼r�:G�q�M�?=tΗ��"�=�{�;�k��<!�`m=�� ����_����|��xԽf��<Ø�=����-����^ɽ�/��+=�#�<�ؤ<��<�ŧ<"}j�H2c��,�~� >x�ս���<4=(����WM�[�:=�~��G�=�Rp������ͻ<��?=�F�<YY��p��;�
�nl�=�1�<��җ���
�=�#=R�� �=BB7=�Y^�ypZ=���<��>;�!�=&��= 6��DR>��{�
X���y�=p�H=�ح�y彶����}�����J�	���T�t�&����=�h���->~=e�WK >�.���'^m=�m�<�p%�[��=@�3���M=��7> � ����ːS=�җ��Q�=�!���G����f;R���?�>E"��E��=/U�ג9>��	�@�G�K㑼H���=�I|��b�Gk<~=�s+>-:>�ۓ<>��b=T�� �
=�b�/���)v<#�ּ�7"����K�>�z�=�56=g�r=�ͽ�F>�)'<�9(�	U��ܠd��װ�����n=`ƙ�>,�Qؔ�7�l��� ���j<��)=w�+<����u��:�kP�H�=�9�=�Y5=�ټ³ʽ�O�=�X�<T��<(�9����=����d�=|�=ن=���#���2�p<mޒ<��=�	x��	��V;b�=S�<�B�;����,��0p=�:ݽ֗�<9���;��;nG��������h8νj4	�����+��<��=��m=�5=`=|<Ň�=��D=�nL�f��;>�����W����=��=��>���<�_2���ڽ;=´Y:t
4=��`�s�>�6%=����QƂ���@�|��<H��=�∽O�غu2�������;;�н���9m�;�}�=���oXa=�ă<��������n<u\�֍�=�`/��q=5�2<KD�=�vʽܑu��<��;D��)a��EP��g<=3?���� �y=��=]u3�H�Ȼ.Ӓ�?�=�������%>����O><Pn>O��=n��=3��<��x=\ܽ�y�=�FI=OJ<c:�<�Ҽ������;E�ȼ�z�<,yM�+w��� >�~;<�=u`Y��ϓ��-���*<��i��p���'�>�Ƨ;��<�e=*�<uK�<�*=�/R=m�]=v��;q��=��?��Î=�J���s`�^v��L��z�<�Ԗ<O�=��a����<_C��p�F��{�>Y�>}�}�c��=J�%��x�/^�=Q������f8���=���;w���f�>��=~�>I�>���Y�U���Q��I�<��.;կ�>>��=�9L=����(�ټN�^=�딽�Z�=(RB>S����>��۽�)�� �]-��B�>�L-��У=��=&�X����=p%��:�*�a�*=�K=#���v���5���=����҂S��n{<W=��<j�f馽і���.�����Ne�y�>>�a5��B��+X=7�������4����<R�>'�5>��-��E�Í>�,c����ݠ��"4��2�3�9�g��<U����M���KR�c^s�t����x�=�ϣ�j����?�=����d�T=3��=���=�G=h��<��>��@�h��=���^�B��\�=����������=�n�=�7�=����$��;:�z����={x꽺刽7���(���S��<���!v=L��;��<��)<Qȥ<\"�P�U�9�\=��p���U=�r����=�h[>���:�|T=�/���_?�N�X��%>C3���+�zɿ<d�ǻ�[�y�=D�#�_��M�=����W��O�I���>4� >�r�]D=�r�=�<��n�Ǽ��=�BD<|�eZu;���=K� :E�;	)�=�f~��ݾ�½Э<n�y�@�<��+���=�k��7=�L�<4;��z�d=SP#=�Q�=Q�=XA=/AϼV<lT�=;ˆ<"9�S	�=s&v=�R̽j��L>0�Z<24o��3���~Z=��=;!�=���;;�Q�@������=�OQ�o�{<�6�<,�*��l=���=3<Q*=���<�=�~E<M��=�eG<ڼ�]�<r����A=8c�<��9��Ƚ�ҧ�B��=-_��ʚǽ����=��ֽ��<o��Q�$��&�=ϙ|;�p�<�w<���
T@�s�ß�5ݽ�C��
�L�^b��y=<��<gO=�@i=�A�=��wuX=]�p='�>M\��_���=��)=��=1O'=A�I=ы!=���<��q<���=q �r<̐��R�<�}̼EС���t�>4/��#%����=��	>���=���;�˻p����BQ��q��$�;=M����	�	�/>r#*���/�|&�>?�K|K;h��?O���8=�{�=���b>��=ę��]s:��@>�],�忋<j@-<�Ί=��	�g�����<<��D>�#>e*>yil�_#=��>ҥG��,��F�=ً��9�׼�Aq�d1��	�����>���~����3�A5�>gW�=�����#e=�Q�=��>���� >���=��=�;t=�T��̞�7��H�Z���<��ļ�8��2ﭽ�.==g�=���=���i�;ޟF</�B�Q���� ����oy5=��<eG�<��H��=%�s=;>v؅�� �*�A=�>�Ƽ�Z��s�6�v���nR>U��o�!�卄��麽k+���+���X=aJ�Z=�k\� =4���2m�����:�;_�'�,<�=#�<y��=��;&��=�	���O�ڹ:��F�=�U�<`u�x�C��?�x]���U��	��&�=o��<��?=��̼)�����e=Y�	���R;}>=�8>�#�=d|�<41H=y��<�=��>=t���qZ�=9	>Ռ�<����k����=��=#���,>���=|o�;�ȽVu���ޭ<4/>�<=i�R;� $�}/���,==�$�=2pS;<u���Aڼ�����&=V���̖=���� Ii>2��aZ=t�F��+=
��=t�=�a\>hV���;�����=X���o�/=Z�|=��;K��{l���ݍ�O�4:��H=�u�Fk��&�l7���������;���=�*��V�$�=P鸼�s=�õ�C&c=���<�]��5d8��_'���0�DA�7�����}<t��<i��=�b-�.7��V>��<RX���y���޽�d�")���4�=�(=<�L���2>�gм<�ͼ�g����DսX{�=��;�׽����W��|�; �f= �>�2M=ur=.�@�!m�=)f�I��� �E���3C��W�ս��:�j�=b��<#��<*=}"'=uV�uS�!ݛ������u=ݮ�I5 �ar����=܏ɼP��<ψv=A���f���*�;{��8>"�9����Lf�+[��ļ;	��=a��<�	>���=�ߜ�k{y=�':MF<>KC�9R=��<�>�/5�=��O�S>�J�=��t����<I6�)C=��=|��;�r����1����Gü$;�<��4�͙�=����\A��K�;�Q�<���d4�=۶c����}\��di��)��<|���=���=��λ^�e=��s��'<��<�������;��E<�y��8n�V3�='L��K������So��촽W��=E̽��ֺԒ=.܉�U*>�L�b��x�S�E�f����F�����5;"B]�̠��5�;�h�T%r=����*�����=9��O'���9��F=����G�<&t�<[��=F�v=�K�<z��ͻ�C��<w�ڽ�=�F>]#�<=���?�/5�5��=s_˼\�,>�ð�%�=��3�9G}=q��<�~��?��<����D��#�j=��v<�Ȅ��
>�6�=U+�������3A=�d�Ua�=mڑ=ݪ�=��=�oy>�)~��g�su3�H�n�%K=9޽=Vmv<����)Ӄ�h��A��7�{; �޽�dڻ]C�a[>	'�� >sY=���<��=���=���=�>���˪��I����=���<<�V>^�=;�`pJ;�)�<}�q;)��T����Ľ�⣼�6��K�1�<t =�v^=�䎽���=��#<���1�=>�'�n���=�p5>a͇=�.������Km=C˽�p'=���<z�@�em���3=sٙ=��ýa�=��ý��h����:�k=�K������<��T��t�����>��y��(>��S���=
�D<��=�-�<PHͼ�wu<fm�<�څ<6t��K=#UO�u�=N����X�=�1�<���=�>ؒX=����A�>Ã$>�1;��D��?ǽ3z�=��d=��=7�=���=Sy��o۔�$��>�p����<ơI��ڵ= }�:r^>|P$>�Z?=�3!=1�/�ӽ=�+<�V��J�)>�����Ͻ�]�=v�$�F�=��ܽ*�ѽLw���(>I�G;��C�F؟; v=����=�>�(X�<�(��P�1�9>�&>��`�����w!�=��:=���=���H'��N��y��S�=3��<ի�:�3���7=s��<�:<IټU$>�;�=1�b�I<�;���=��o���V�+���.�h�T�����V�ü��`�=��ƽ�H��6�ZH4��ڪ����+ߺ=�,3��%%�v�>�w<�0%�]"��Nb>�W�R'�=� ����2�^�=nJ���5����|=8Oͽ���p�=^S�=�<ڌ�<���;���A=�寽bF=훓�N���J���#T�Z�K��U�=`�8=C8�/D��:x=u,�=6z��{�;͋O���>E�2�K�=�ݛ�>�,����D��=��+����Ǿ=.K.>.�K��l핽N.�= o������d��+�(=˰��j����=eS=���.x���E=F?5�G)�_å���=�c^=ԛ�<3`;=E8�T
��������|=�����+>��=��Խ�LǼu:e:Vy��<���I'�=^'���{�=�?U=V�˽�{Y=��!=q�.>w!:=#*(�ޞ�=\�=���L��=�_�=��M=޻=*�<�pK<L&��!Q�<;|ʽ�7�<��潶�!=��=�'�=�j�ZM,<�x�==$����0>>ke=�J=6����	m��y)=�<S�0��<( ����=��/����=���=�4=��%�=��;@����Q,�fB���Ƚ���=��3>:�<�i���=�=tf*=am�:�Д��+�'L�= ���� �~쇻�K�:N�����	�u��;�o�(�3<����� �i�>�R=	�C><�=3!����!��͉�(��<��%���=�J½���ǽ�Y�|����!���:6=@�=X���)s"<�Pc<�2ҽ�C��Q=�1��f�S�G=�^�=�<�z��;8�����<AZ�;��\=�b��Da?=�L�mU=�	���ҽ;��<	�r=�T=0p3����=Z��=�{v���.����1�ռH��=���<l� ���$<�cb�q����>d3�#�=�Z�=E�$�$=�H���a�=�X�"�<��X��t��.f�=�-���_<��N=�g�<W��<}�="��=@���������Z>;`�=�����5>��<�)ټX���:g���G�
�w=c�I���[��<�n�`�Ƚ�o���O��l0�d�G=�\����A��a���Ď�,ُ��޴��X=�W��ͽ���<8��:�A���	�[��'�<�.�=���=��F����;�˫<��n��=���;츽[㼖����<B��V�2>�+=��p����ވN�l~J;�/j�L�=C@�=$�r=�(�[�2=�#�=%�;9{�bi(>����=����Av<�9�H�n������=��=��>���=I�-��O.��,u�Sq�=0:�9L�f�0�ؼU �q�&�SА=T�=��ƽ��P<,.���p�=��]>�l�<;�=��;�mư�s���p�a�׼�s=��a��ͼGá�_�=�Z�=�)Ͻ6��=/\�M�ɽ�P�E~z�� >n�>�.<X�->���<,���L��G|��%�=�O9<w<�=m�9�(�=��.��Ò<�E��>��m=J��=$Ǽ[�9=Yφ�vb�=-�<s�>�==�	<����7F�<bp�<�̽d<�C�H�M���>�v�aT�<cs2��Bӽ�?�=M �<U�e=��=5��<s�F8=���=��W��b�=>�	>|B�,>�׽�>�Ǽ;��=�G�Tn�9�3�k��=WA�6Zi=�I�hP]=�8#=|��Ŗ��=�&>��ý%
=��,����=)l�����=���<k��Y�=F���7�Vym����</�s����1� >�����g��ŗ=��'=����<�䞊<r�x��(�=�<�4)�=E�~�2a>�i�� v�=�N�ã�=�<=O(=j�����)>�l��Z��51ʽ#	�=THʽ�R=��E=ł����>
f��Ob=�۪=���=�C=�߽B=�T=���<�żSD<���;a#4=T)��>iV�:K���z�=[���=͹��>~�!<r7=�!�=OY=��'����<���dg=�����>G��=U�G��5Ҽc�1<fUT��)�<�e��<����J��753��9=ũ�<3i�=�D=�E[�D�ټ9��<�/[����S�W��>c-ý��= �=��_=d�=�x�<����%�`��?;��͒�NO�=��.>@������=��=�B��!=W�9=dM�= �=��㼧^(���'<��=uP>=˥=���<|h�=�h=�	�=�d�=[�������$=aM=BCu=)^�<�/>���='������_jҽ;^�=���j�f��k�H9�-�=w�D>���S��<�B���=6>=P_���=sg��8�=}.>�ӎ=��k=�=:��M=�s�χ���O���'#=�v��o/��lƫ=����͜��n��m2>P;>(�߽ƺ�����Uh�<�>�/�T1=o�$��
�=}�p���W�b�\=is�;�k�=z8/�'ۼ&w��F�Q�=ȥ�;5��	�sW*=v�ɽ�\�����=�!���|��|�>�t<�J2=F����������"����̋�gQ�= ˄�˒�=Ip,=��=2�L� �=%��=*�<3_\�ڣ�={^������*>��=ڙ!�M�x��P=^��B���V<6�;��:=��=aEN=��=�yv=ՓB= �=.�$���<���="��<�����N�=��ͽ�����k<�Z�8î���;�C>��ٽ_*`����=�d=o�.>�.��`�z�ث༆�<�[+<�T'>�,N=�I>ގ+�%J��cҽ��aF5>+mL��)�<]˽<�W�ɣ�<g�l=�
>]�t��M��aL%���=�.��k���ī�23���׽�a�<��ͼ�u]=.Q=�K4=e���}�F1'=�H��~C>�E���֣=�hݽ	|����=:��������<�⽀�2=M�����vQ>���=z�&�!'�=Q|ýi���!g�=�ƻ����ĵ�i֜<i���Ҍ<,�{��b�<�ؽ�\�=��ͼ���d�>%�A=P6�=��X=J�Ľi�e=EWm��姽����Cր��J�=�����Z=i��<k+E<��=����<��6>�ԇ���x�=2D�o��<h�
=i�>�&���aE<|M��_.ͽ�6�=�m!<mpz=(RQ�������;�Nj=/� �f\>_=Gkc�]����=�g�=�#�;)��<�ޫ���Å>=����i�=��t��ɼ`¿=�TI�h��	h���<�[���:�<i�=�r���+޼B�:ƨ=�v�=Eh�=z�=��^���ʼ�eǼ=�ƽ�ܚ��j�	�<(;f=��y=*>I�=o���K�=2��WX����=��=����S�=.0=�Y�=�q�=$��0��We��0Yټ���|�=2uн��8��*y=*�������!�8�KP�=k�A�G�N�8#�=�ײ=��;��v=g��<�@��#L�;�E�<���=mL�=lJd<g�ǽ��>�{���%�@�=B�	�O��=�G�=�+<���<E�3=\�"�=5w��1�������x=��ཆ���0�>T1�9b6��W;�<��~�-�]>�o)=�9�����9<����=9��^�>u@�=�5�Ãi�虴��H;���ڑ��Q���徼+@!���=켩=�'W��eW<�1Q>�)���#�SVl��˓=Fa[�DfT��c��h5>|�i=���5>�b!=#����>"U=�鮽�&��U)�=�뽻`�<I5=�=/2�=]�>-�<�9�=����|=nǋ���
�e߽uV����=��4<f��?k8>>�|���ӽ3&��;����=g�&=t">��=ꂻK�=3[h=u�<��$�=yŦ��%���A��K�H>y�7�c��t���<�Q�Ͻ�Æ=w���S�=��{�����S<�ڼ�';/�=��ۼ��㗂��=P��;�8��-V��D>/�><���=j��=���<���=[h�;C��=�q?>��r=�V�d<� ����O*=�	�m��d����->EE
>i*���	�=B���F�=ĝ�?�<��1�<���<�m�d�=2�b=�-=O��<�8��Cн4ݘ<�Ib�v�=һ'��M��|��=9{=u�=r
�RS=^$F���0��l��S'<0�g�A<n�>���B�k=�����*%>�h�<s骽؁=ޥn�=һ��ҽ�nR=!$�=T��Q }=��f=�\
=��=���O��m=�}�Я==�S��7ʻ����C>���je�=>jV=�{ֺ��v�]t��=A�<&T�nʕ�dK�=ڋv=&�$>�DB=�������<I�n��S���9������.|�l7R<�oܽo��<}@�<
�R��!&<�^=�*�=�!Q�h+��U	=�.�]�Y��⎽&8>N�<:���@���� =�ʛ����<�� ���=����nq���P=�x$=iA=U}�=��H�@dF��(��3�q�2=����=q�P=j*�=#h�<���=�2>uN�=��=�R��|-ڽ�W�;�>����:���=�=��ؽ�ϖ��=wž��*#>��<��=.~�<��̼x7/=h��=�����=�m=�q�=�,�E��=dn�F�z=z�*=���vP�=2FM����=i`r=d�/>P9�=�����b�<�]�=zL�=�d��_`��R�=8ܥ��.�)k.�K����C=�e�=�[=����s����].�TH=_U�=Ȍ�=�D!>n��<᪞�Ú&�q����>��
W>�+Q����C�O>c��=�9�=4��>��G�'x�m����=ny^���-�������=�v=�8d��	>R�=��"�於$�<q�<�,!=[pۼ*W=�w>���9R>�3l��1o�X⌼�q��XZ�/)�<�����n��ɫ��_�< �A;��!�v�-=�J+>��K�q��o�o7<=x���5>gG{=W�˽�I>Z���3:o�V����7��MH<���>l�=�9�r@�00�!�:�=DH=z;��54����=�`�=c�G<^�9=�ߵ��4O=]ü�5,; dż!A>0�=zk�	����=d]F=�'=X�)�X<σ��k4�<Lȼ�o>�� �أ���>�9=<����ٴ�֗$�])P�k�}�=�>o=��ؼ��6�ؘ\���'��RB=���-^�<.b�=��=��O=���=���{���-��[;l�=o)��]Z�<���=��q=AS��s<�8:s	��e�=ǔ�=�AZ�D�C<X�<������e��vY�vvH=q���Л�aq
;�
&=
���R>?��x>L��<�$߽��h=') ��ο=M���4ه<x���	�=�%��$��=�	��&=��}���="��<�٩=NԂ:z�r�И�<r�=�J(��M��,��z���9<t"=��>�L�'���(>�����8�Y�T<:=<��̽V�==�>�U̽ҵ�ZW�����-�1�<TG�T=�=��Q��^ �~��=<�a��lj=�	&�bQ=h*���>U���lK�s� >�4=�	��� >i@��T�=r�T=N׽4ы�]�>(8�=��ӽ�-V�,n�=����OH��$���BG=�Tμv�$=��a=%�s=��M=s��=����)��PV޽���>}��<z��=�n/=����Z=P/�=�9�U�;�|b=iC>��@=I����)��'�<�~�=A|&<��T=U����B�*Խ��<Rի�E����=�~&<L&=k�2<�P1�ɂa����\m/>�ޭ�|��;����>y�<X�>��C�C��;�}�=���� =�s�s�
=�����=�}=)y�=�h=���]m5�.P�=�b_����Q���$�<$;=����w=�0�;^�<�.=�P$�VY>��=8�M=O��!�
<̳(=�=_܊�^_Q;_���[	`=S���WNT�鑖����<�U?�h́<�����ZL�SHM<@Ad=`�<݁=>�=e���]��=]��=U���UD�=Z�=��:�n=/t½Py=�����T;uD>-��=ɛW=4A�=�i1�v�=K��=ـ�<>\�^c<?J����T��t�<BK=�@�=O�Z=`I�<YӼ$,�<m�J���=����廻eG�;�P���.<���<�5���Ѽ�K=�qC=�Z�=�I��L�=�^=~u�:c�
<	a��$�c��jM=�R=;�1<Z](��@>|��<��=%��=�	�=�" <6�(=�?*�
6Ǽ}O�=zb=���p�;���P��P2�=t=G�A����<}UV>�aؽ|�����:��[<t��g�5�d��<pB(�HY��p;mC���� ��p�<@V�����=w˻�|J=���=��󼫮ٻ��=g���='m���=$�=�>�ý���=��j;�DüR'_;������;�g+=+��=���vr=��Ľ��*��:=��<X�ʽ4G/;�U;Z+����1�$>��]10=2�5=���=K�>n�=��<Y��=��>�s���촽���=*�=̊A���M��s��qF��{������r�(<����h=3|����;���`=K�����>��P ½:}=���������'>�4ͼ=n�I��r�;6:B=
%�6�Y=U1=��1>��n�7�>dtǻ6%�����=�ĵ=a�>���=)�=��=}3�=P��=롛=SY
>�$�=�ǽJ/Ž4� >Eh��ϖ��Q�=q2>Yg�=�����<EÎ��M>���-�x��	�<�>�}�=(�Z��N�<e�>Z�=�����n���Dν�1��O=��>�
=j�=�9�=��">'���<-��L-���7=��<��=�˲��;>@����0ҽ�{{<��y��S=����^��>`�}��iq���= /ѽV��=��=����/�5��3漊��<��L�Y��<ڞؽ3��;NԪ=��:�f�:=I>��R>il.<D&��kI=f��)'<Ŕ�ZU�'�=Zn��D�Z�wD�=��*�2��&#B=����4��k���=ٚ�=�#��s�=��iK��߼��@�K�-=|,�=I/ҽ`9-��A_�����Ē���+�K�=�g�=(����3����<�>��:�)������p=�蔽?
<�L4>�%e�G_=$~�8�=
��]ͺ�;�4=o� =���	K$>뚽�)n�����B=7�A�m3�;��/���'�
�p;�Q>(2�=?M�e�ý�}��C���=���=�'==�b�=�����ӯ�#�̽P��<�ý^I�:�@�<�=P";�>ڽ6�=�6ǽؐ�;�#��>��3>�n1�ո��R�Ƽ2�=�����1��4=�D=5(�=��=����<��M��}=�n>�~���dC�:���=�a�=X��<�d�=H0=祻��=�i=jń=�(�<狈����=�nĽ�c���z�=�հ�2���z�!�v�*���=�L��������=U��<t7���9=z���\L��O`�S�b=^����2><�dּ�������J�%����=o��w�>x��?��f�f;�����3ڽh��=��}��	���>􋾳e�<�v<p
κ�W�=�j����t<1#����=�Z�=A��<[��;@�4>
(�=A>O�=�c��j ��x��6<=_����]<��н�ʃ=�͙<b��<�Ҽ
��<rʼgΦ=�ӳ���q�c=�j���L@��,6>��=w�/����9P�ҽ�W��~�<�J�<��x���=?'=�<��>�0F>�(7�d�=I8g=!{��f��=�D><Ȯ�=)��=C�6��#U��z�<ō�Ԩ�:�ɽ�۶��p�=���Ov(����PX��a�Dʈ=_�%��g��s9�<ǝ;m
�a�^�X���=-���.�g�a�	��=ɿ�=ӡ6���>;ν�]���e=���M��=jb�����<��
=�A�=qZ;y�`�˄u���-=�ڹ���_�z9=*��<���RC �(�����O=�g�=�H=X3>$�=�ن=�HF>�3w�Ъ	�1(���1����<�e�%>��=���= �H<]��<	|��R��<�2ǽ��>���<���;5��=��<2>ܖ+=�����{���r�<�s�$��=���=<��Ԧ>�̻߃">��N�����U��=��-=]�ɽ,�">Y�#�k8,<�=��">�b#���*�2><3�=�[=���=fL���=���=^��<TL�=�X;�>L�K=�M�L��Ւ#�3m�����<W�н���
=�����=R%�=̰�=O9��0���wUi<	f���=��;�6
��,�=��R�'d=��ƽ��%���C�<�$�8�ə�@Ǟ�^�=�� >$@��I�<�o��\o=8� �3ν*]�<܇=i��=>=��w*��*}�=U̷�H�j>��3=��<��E>~�>��&=~-^>�= >�l==+&�=�8��I���j�/=9V�=�N.���=+�;�=�f�����9I��_�=�y�=Xs��#zw�J|?>"s��O���
��H'3�3�;�s�=��(�3���^��=T���E<ོv+�==�=�����Z=���=��}<��<�d]>`�������d�H��<�i+��p=���=�r��0��=��S=��U�X6�=�=0��=x�w=�w��s���*��ڀ�?x���Լ�Db��W.��Z>l$V<��=9�:c���� ��u=|�e=*#��&���M=��>�<���<i׆=��=�Q����\;�02=�x">����M�Z�~��:�#�����k��������=q�{<G�;� ��r=�>6�#=Ym;o�I����=�=�o<捠=�2i=Yor�I���L�+�^=�,�����5f�2�
�6��<&��=�ź�tk�=�`<=�W���>X#���[{=�!hA<t���K�2<=D� _��>�==aE�=˓�=� >�O2���;��f�І�eq�=z�j��ᙼ��=ʙO��Y$�x�<>��<��e~Y=�ί=���=&U�<�Ž~:/=х�=<j�=EY=4���ռ�d�=^�b��<�<3=.�7��J��Jb�M?�<�o=�&�:��=�=&@�=�S����
=����� >������������ӽ!S=���/���g=&x7<�bǼm^�=ڱ<j����b��Tb�AtP<��U<`��<�ԟ�Z-=���=�iu=�t.;~0�<��m��4j=A�=�Oད헻�V'�Q3)�R;�<�D��K��=�z]�fA���=��,�;��	�d���-� �4=(��=A��=j�ý��ü�W���=���<%Y$=����S��<�J=evD��==3����=7�N���.�l������������g;��=��|<|.d=�=�|ʼqg>=�Nb�qe3>����9'/����{i�R�Լ��g�#=g2>^i?>V.I<U��<��=��	=��׽Ak����W�{�����8^>�m��3"��7=4��=��=��=���,=2n1=���=�	�)�w=F��Ol�=�rQ<�,�1<S�J&=�7� ��=��,>�]�=du.=z�p0�<��[=O���K��/ݽ+�#=��=1L ���=�Ͻ>��oK�=a���'�F�w��=�����o�=�=���=�+㽼÷=&���w��ת&�g��D���ܡ�<�3ǽr�<���<ʐy>E4�hCȽ��C=���>�_���<q�����<�ƽЄ�<DQ<l7�=s�]>��#1
�2�\���H=m ��[-��W.��6�<9:�BY��*�J=(u�<�K(=V�=�����2�MX_��B�<\>>�+V;Mj}��#<�8� �����Z9��^���<">�<�����R=Mٽ=�.�<k�>���,�i=���ݑ���@&��b�<�=n<y'=ңT=�u��+�O<Ŝ=m
ǽ�{�m' >$xN�� >|+$��$�<���<;ý�M�K=c�=�	��+Q�6dH='�E>+b�=Eʽ�-������=|���մ=/��z�c=�� =�«=�a��!<��*����=%�=�}�����:�=�Nx=l�y;������>�\�1[=I%(<Ω���>��mq�<�j��iő�Q~�����#�=O��<Gc�<"�>�
����H]�=ڊ�=�-�=��}��Y[=>�I<�o<|D)�UQ=�[��`�=�q����=��z�������Ƚj$>-�WpB��,�<x������)����=ϵ>���X!��r�=.�㽻�8�ӕ��?����<Y�<�`�=>�5=gQs<���<A��_:�=�������6S��=b�=��J�����:���m��6�<�����G=Ӷ�<tWG���+=�?��_���9�:
S=,F	�/������=`���Լw=�_+��?��������\�=ㄽ&��}�=:�<4�"=�dD=�3���g��p�Cf&�	�6<S<��Ձ�=4�<��<��JY�|� ����=ү�=�'`=6T����I��<��1��K��=A�н�#>�x�;MI�=D�=	���*M�W;���ټ�<A�1V�=���=H��=(���>��=�=����^Q�c�S<"�B��"��6>[��>�3Q�ze��`~�=m��<�)��z(�=�{Q=c&>Q�>�N��v>7@L��>6=���f�=��'=ۚ�<��S��Ƕ=��
>A�S>ƅ)>�U�w���E��%��	ν�/�z�>�<��$�=#$�`s��d�=SD>6��;��ýJ%)=X��i�<���>�=�<Ɇ�=Cw=��
>��<T�K����w�<B���X�=i��=ȩ�=a�=Q�㽓�;�o�=}vF��h�=�g���gx=1���l1�|4<�n6=2;G�ꛧ=fD=�T�:P%j8�Y=q�(�[8=�Gq<t�	�?s<0[�=��=3�l=�T>r�ǽ7N��3��J���0�<e��A���Oe6��~��;��<s�}�Xz����<D��|�w=B�=D�;KI�=��>��ܽ�^>>ڌ>>�Ԟ<8�W=mP�=/މ<M���n��N�=�f�=�;���If�T����e������F���3=0�ʽAp�=j>[�_=X����f�{C�=�w�<ѽ�=w�f=���=c����֦=Qͤ��C!��Ż!Al��]��]������=�������� N�����9����>r�м��<�f���񼱈=0`�<
�=j� ���H=B��<Lq�<A��<e�<YI�=J��<.��=�(`�D�=J�< @<�#��t^��m]=d=d\
>�ʺ��eѽ#*|=R.=�����zoi=��O=
���೼���=��>j=Q��������=s�x>@��<[��<|=CѼW�;�TL_=y�R��!�=���=V�����>>�f�A��=���=zr�=�ݳN=��T���<F<���<!~��/����e���ԼN �p9�=OK�;��#��4��K�=y�%�oMe��u=q.�<Qσ<k>���=X�a=��I=�x��ߢ-<��<|�轝*�<�v3>�����J	<ߟ���L��G�=DW�=������<���=��<w�=�ܝ�￲�[��
�ɺ= Y���╽񂄾� ��%=n?=|s��hy<-�=����B_���K�]��P"�=9� �f�>���}�=o�l>;��<�=Y�Q��D\<�!���R�=�VN=�/���?<$��<�yS>�l�<�=7(�<�6<��J��r߽��Žed��<5좽*�_=5�=v�o=�L�<�ʍ<�*]<:���J�X7�'�">yg&<V�Z=:�=�m6�d �=��O=*&O>Y/��i��=2o�k=F�=%U=u%G:L ڻH�;x�<0EֽAa�=�g ��>==@�f=��;��ś���X4�=��i�أ�=�S=SX�=O�D�DE�H��	���I�=c��<MЁ���.���?�V$�PWٻ��<��潻�.>u@$>�V���z�=�򽿗���ĽE,��0�=d��=p�ĺ��o�gg�<�67�N�I�/�L�:���쳻��w<���<x�K����"Ļ�(	�J\&<`�����=����<5��n���p=�+��5</>~|M�<;>�?>J����:��}E/=ٸ�=�K�=�Y�;a=w�U�u�G�=׵d�Ryg=0> ;^<�*�YQ<mY޹���;^&�����<x|Y�@ma�T��=�b�=��P�Qq"�,
>[���=�� >`޺��=��=��>��=/Ъ9�#;��z<��@=�⵽	ϫ��p�=��]=@�c=�
.�j�B��N�@;��6<\[���l��=P�;C��=����ݽ�{�<�6�=����4"�և�=_��;��E��L�<��
>0	�;_�K>�ۼ=��r�iYd=�<@��=9#6=�:,�B�<ﺛ=��9>�a�oK,=�n=X��=�-��B=���<�fԼ1�;�7=���ɋ�?J���=i�}=��=�_�=�2>��>R��D/�=��g����k�9=)��<2���M��H�u=}O�h��3�=��
=�(�<���<��=�x��!^u����>��=�4����=KZ=\�x�S�����ͽ������A��P>��M>����
=CGt=��@��t>)�
=dn�=G<Y7=��`=�A�=�2>k�m����=T2=d�r��/�u�R=��<��>JW =��̼W���J���l;�0�=�=]7�=�/��l5�;�܌=l4ͽ��0>#J�<���=��o���=�O�=�=�L]��5=�n˽[�=2G:�����+��ؤ;��:���=�|.;��>t �=h1�=���J����F�<��
=�=�6x�M�=ޜ��n"¼��:�t�7=�{-��Q>�^�;M��<�B⽚���}�<���8H��q8�;�H�;,�彀��:��Ņ�=b>>��������vq=&�v� ��=Pw">i�=��z=5�"�.,����"=�d=�A�1���F��=..�=��<͹(=��3>��#<�(8�ܐ�<6�>�=a4"=�M�=T��=(����(=ڙ2="X���W���9��S��&>�J����[l۽R��AZ���	��	�[i7=n�#���<�)!��襽�!4>-����=1K��&<;K�<ɢ�H�\)=�<�=�:F7�=Wu�:(���%@z�x�<M�]=q�6<�Q<��>�/+=��;Y
˽PZ����	>��>r��/��E�=�ue��{=*k	=_`<�E��j=,U�<Zo���:4=	��e�<�.�F�3�+�=�<����h=r�\;�>���=;�4�=�ζ���X=�Ɩ�kP=!N�>�Y)��"�T���"f�=+�q=\�,�.>�L��=d�=~l
���@=�c�=��Q=��=Yy=h����G>M=ttq=���;����;������B�i?��}\<�=�&>~��=�� �U{=��ʼ�>�B>�<�N��=�=>� �EZ���[��Gz=���=1=��޽�|���c<�K�=���=�:�<=�>x�>�w�;?�e�83�*|G={�F>?�<c�j=�I;�%�ڥl=��=�ǽͥ=��&�q��X=�8:/91= [�����=u��;� m=�}	>g`��"�<^b��n0"�G]&=-<�=R*h�}��=�2.=�<=cݷ�r���� >*��=Y��=p׍��'�����ƒ=(��=��[�����s��ZT<�m�=��
=U��*�d=�=�=E6���n>^G�=p�$�DX��O��@@=(<�ӯ���ļ�臻aq�=a�<�q=[��=8Ξ�x�录`�=���5�<r[w�s>�=�`���`Ҽ�. �cTs<#B^=�U=֍�;��=�8=j��=�!�Lm=��<�fC<���=O�P>��@����:F��*��=�=�*=�9=�0:�)7̽�Ž��E{=�(p���8>y�=xk=���=C���BR�[\��Ͻ2�=Y<rFŽ˴]=�V����>�)νj k=Sͦ=e-�=�$=a��1g5>���� @���T>���=����j�=	�>����sn_��9~��<O�u	/�WL�=�V�CD==�
ֽ^}Kf=���%�d=��½'���7t�;@Q:<h{��0�d��\s=)ð=5ˍ�G�<�-=I�T=?�>�H��l�3>��
�B�w��/��;`��Λ��f���+>�y>�<�v=!{�<ⴼ-Ԡ<)Q�But=�f�=�5�<�=�n=��=�i=�	���-V=�.�<��=V���:�=vl�<3�,�>�=u_�=���~� =�H���f=*�ʻ�#�;�]�=�J��v�;)/��?�
��jv�<9�{�i��$D>��<~g�:���=��AYA�B��=
̻bӽ�l��������=�Ǵ���==R =����L�<Rܻ�Lp>�{L=�x�=7���>iɻ��Ӽ�Ȼ��w0�v�f����=F�׽�=��Oӎ<�=��=�d��7��J	G=�<�='G�<$GQ���&��a�=ˉ�K	����r?;> �Q=���*���1��N�{M��&����k�ؙ�;l��<�*q=�rp�X�=��X�:�=��~=Qc�7��=�V={e/� �U�S���P1>�Ƽ�!ڽxI��!�*�@R>�	���׼-%����=@�H��+=w�D��֚��=����<=y>�:c�ҽ=	=@��=�1�=R:����=Os����A%���C�1�<p⯽��V��f=���=��=AFz<���$>:��=��&=u���$Z1��R��~A��V0>.A=!9�	����W�~+=��X>���
����q����=��=�ؙ�ú�<{V���߷=�t�=��ĺ��=�K��<>����=8g�6�=��=�'�O����<�s=핽ᦟ������"�R>��wÀ==)�� �=4�I=@��<��B�L�����ƽҜJ��>�q�<�P�2E�L�x<6c��>���&��ϖ�=�Z#�D���"sٽc�&;6⻽ڠi=�?*>J��; ��h�=DeH�7(���D>�5<�"W�<�P<��M���<��6���
��i6��=��� _>U��މ��<�9�]�V=�)�=��x<��>"�=p��=,0��q��:"BļP�ܽŶ���A�KG�<�;O=r�����#��s�=B�<�ı�������"�>�<�8��O�C�^��;��=�ϡ�5�ܼ!��=��=*G+=�G=�^�=��h�aw�=��<�Չ�s��uQ��W&�U�0>q'[>1�F=��Ӽ^�K��-Ƽ͘ټݚ��Tʽ �>�e��dn=�=�>��;~;�=���e��=<Q�=9��܀<~=�M��F��=����5�=���<��{��1="�<�Z0=2�=y&=�^��@#���=>��<��?=�?=��D�=�e*>�<�)8>���/0<�B㽴����L=+E�=�<�=�K�<Wˁ�z;k\�<�q�[pd=~>��(>�ֽ��=�d�=����>��vʇ��ܹ=4�=O�ǽf�F=?�;*�Q���H�V�= ����=�.=YMd=I��<�`l�����PGW<����&������t:6>rH���v>~�'<o�;�)Ͻ/�]=�u�<�D=	�L��Y=�����'���=�߄;OXk=��ڻ��<���gԻ��<Z��;���=ZT#<�ܘ=����o%>2��<TU��R=�gs=�į�=��<��p���=gЃ=�:=����<)�<*<>@l=�:;�m3��b�_B�=rӎ��\X=J-�<�K���0=-6=;]�=?:һR��<I�<�$<��|��E����'�q�<-�"�Dg=�-�,��= /D=�CE=yE��F���u{�=�\�%2]�Oˤ;�`T<"b=~���G�����=�=��W�[昽�Gr<�A��6P�!�&=��D>�`�o r;h ==C}:=M���IA�N�<�<y�z<0��%�y=�|=�F�=��8���=�ω<��.�+���m=�`w=І��F��=ٞ���V�	��=��=���=������F�=��5<���H��h�>/SO�,$����0=Ȟ�;ʝ����<���7�z�L੽�6��1;��
���6�%u;�\=�<���=`�/=�]=�2z=�e�=X�*�gܡ<�ң��$�=��E;�_�=�D=��<�F�<VKt�5+
=�)2�S󳽂c�U��>P�=�f>�-=�\'�B+|�U=姽�O�w��>3�K=>h���=>.üwF����(��x��X�>`�w��Zb<X�oP>����|�ۼ��;�ŭ�4���2>$_����=[臼����� >�尽�}I=�#�=O9/�X�=�$�<����FQ=��<��o=�+���	�'����C<��� =#��#�=��-=v����w�]�^��_�<~��=�=ڑ7����<��=���<�;"<ޥ�Y=~�=;�����W>�<ͺ�=�aH�4)��sd>�İ���=az&>g�=+�h�V"��d��=O�=ݼ�;��-�:_/=vL=�Y%����d��=,-��lL�=����=�U;���ֹF�����#>7�S�M<x�͟���b���:;�gg�6�~=ə<=̄S�{�=pf= ��=�=N��SU�*6ͽ�ة<j�뼵:~=�����3AQ�6Ԗ=�t/>bF����s��=��c<c.�D=t�V���Z=�%ҽ]<������=��R�L�=X/��^��9(>�~�;|����<���=�:!�m�N��E��(7�*��<��s���=!�8�Zˁ���=51�}��={-�f�L��U���c���(H=�Os�H�Y=Ǌ1�)�<����=�Ϊ=�t�=�N�=e<Ř<�H]��$T��N��<�Xw<�6>鴼l>g�Q=0��<�$.=���i±�Qy�p}�����=��<�!=�y<���=�Z>��>�`���U=,�=�U6>m�=�T>��l<�x=�ʴ<�,=3��3���nd<��>0��;mIļ?��5�/�Pn)��@�㺀�j�<}��'��ϱl<��>٣�=t�=;�=^�۽]� ���>n�<�A
�EwϽ2�5�/��"N����=Y�j<��)�%�<ì<����l��<8�����;UG��~�3>{"�<k��e<�E��E���1��<q؊<����]�<He��Z��=��x�w��=�N���~���N%>�
���z5>�1=m���,�=U�4>����\�`�P��(�����;x^�<^�:�ٳ�=%[�<���=\[5=�V=�!=(�~�8�<A��C�=��=�D�����������v=�#�M��<�#r��z>�Ȩ<�E}�~��<�Ȓ�p��<S�#���=#ס�22�����hq=�!E���	��-q��c��s=GAȽ�g=v�=�N�=���c�73]d��)��켸���Gw�w�C�9x��q��j��$��=�]�=Bt)��ñ�ez�=����be;�V�=�u,��(���	����G>0{��"�Ž���<������>4��>H�<���>�d>}�&�2����r=�|4=y0ǽ��=r�H���P=��G>t�<;��=m�=+M ����o��9p�_�'<����]B�<'����v޽L�>�۽Gz/=Ԫ_=�9=E8�<������� ��T���;������������������b}��c�=`.
>[7�<����B�<���=z�w=^����]�;�͝=F=�ϟ�;�°=�m��_�=����f����=�sL�f0ݽ�����~<<��e���FD>�/=�L�=��
��7�ޔ����=S��m�=����y���S���}d=w,<��Ҽ��=�V4=��=f蚼�Z�:��$=r�E�	S�=D�Y=�F�=ߜ��"*��A>K^�����y>�A>���=�E8l�<��"�0{=d�=z�����<.V�=8=Q=�i5�=.����N<<�F>�S���sO=}���r�<@�<���=��w�ۼ��=�ͼ�K�<H	=8��ڿc�r��d�H�=�|�<�ͽ$4a��	����=�X��jރ�i]=O=Y|v=R짽��E������}��χ=A���>=a@ϼѴD���D=��q=1��-0�=�94�g�<g����a��\_�B��;_�*<��=�i9�ܲ;M��-=�4=�X(=�T<c>��	<��<��=���=h	���G��1���4J�� F��>�=���0ؤ<B��;&�y�.=q]E��y���{z;�K">�~�<��4=��d�M�={��>@T���=��f=���*��<��ҽL�G��r��N���p>aɇ��+��W��<��t=�q���:�=��;E��b˼��v����L�<�==ȣ5����=�f�����:L�����p�,�����<��<䫼pU==�۽?��<�S������+�=FQ���|�#�ʽ'�i�V������������ao=iJ���Ͽ�X��<�����;=��w�� ���y="��Mq>��C<c�=S��=�>�
>��;�Y=�F>M:+>���)���%�<�H��O����-��iu�<
D�=��=ׂ`��Z0=;�����]���S�!i�;dM<��	>�٢<A�k=�O��#��Bur���;`Љ�>R�=��<�넽Aˋ=����r'��f�=�f=qŻ��&=�
O=�]7>;�=�B>7~���3��6
��]��B=c����:������'>hQ�=e��ZCX=��R�d��Ž����F�8� ��*�=+�#��"���R��=È��A�=aX=h/D�m�ʼl����=�߽\��C��h�W=��d<��q)��ך��ޟ=� ��H��=��4=uھ�/\P�3(�����O:��(�=L'��������� 	=�^h���=CT�:�����M�2��_/ӽ!��<W�s=f����~I=`s�<��S=U�ֽ�����1>���;��߽�(^=-C�ԓ�5�<PNĽ�%~=-q�=��j=�B>�U����=�\�=�uԽ^6->�>ܾv=�3a=*J��=��=VŽȨ<��>�O�0�Խ�>�a>S'����<�j�<HS��et���\�rh[>�Vf<�SG��	N���ɼF�<&oD=5=V����=sc�=�<9�>�;ƽ��^=��>pG���=	ш<"�<���J9���W;�M�=����fQ�c�L���7P>Γ�=�7�fdy�\�=��;��=�_^>E���c��n.y=�C���<�I����=y��G��>X�r�-�x��G��2f�;��<�C��)���B�=��<N�>G�н��ڼbO>3[D���i���Q���= ~�=��(=b�=#<7=�=�=�0r<�����{�Za�<����SNI���=��k��=������;=��@=��=�4�O廽�+�=��=Iڽr0��Jh��w�xq>�fh=r	+�h-��O�=YJ��N�a<��>�$�����=�M#=�S8=}@�m�&��v0=�}̼��:o��=��$��=���=x�ϽL�/��?F�E3=���>r�f#;�SO<H{G=͓&=dw>P��=�S	���[=G�F<)�����=M-T���=(y"=����������=�>$��=��+��h����W����g�>���Qe�=Y�W��'�g�h�һ'>㾴���#>蟜=��J��O�<�0�=d =����@���>�;,����{9��/�,�>uнA�ϼc|�=Gޝ=i�������1!���;��~=��E=�ļJ���=�2����{��=��=i0�&ƽ��R=MI�=eӽ����|G#>�|�=�_�<�>� �<�z��4E=�齑������1�����]��c>�[|=n�����⽴�!��r�=S_�=<Q#>�=��m�I�O������n���^L>JHŽB}����=p�t�h��=���9sޑ<�P۽>�ݽ3E =z��h��<4[=���=�Ͻ=��$�(�DԱ�Br"=���<S��=K5�;���=�\�=t����=."����]��=oVm=KD[=��ǻ\�ȽrT<��D>x*E�s�𼻾��}��;
�>�������=�N��b=����W���4<���D�c{����w�sJ�;<?k=������1��:�<e��=a!E��W=��ʽ�=o�L�P��9�e,���,�� E=�C�����>J���Y =�[*����<��\�W^<}^&�j�y�\�5<��=c�=�|��kν��=W<Խ�������B��:9�=5{T����S <#*>��켆�=��=@^���a���b`<)%�<~2�=��L>�c<"`��� ^=���ڟ���8>�W�a��=D4�=�e�<����u�����`�<��=�̽�r�;?�����;��I@>4E>_���Ā=~2'�*��=��G��D���=s >�q�����g=s��A)T=�B,�Жx�TYc<�$�Ʉ���-�qi��/_>��Q=df�=-V=N�<�R<��#<�X�<�3�='�I�;�ܻ,�$��^�xRd�C�����R=G�=����g6=xP >Ɠ�=E�F�'�(�qm=\\<�C�x<���GX�=����fļ�p��1a���B��">- 6=Y6;3n���;�S��ǽm��
�������Z5l<\N�<�;Y�=
�<ZO=���u7�=��7���>��,>�.��J'<�`ؽ�<�D�=l�)��fżK5м��\<b�ռ鲣<�Sd�x�=��I<�$��������<�R6���<$I������7�=��=!|�=̅�=�>�gL�gS���	>����5o��O�_%�E�=b(&�s������=��=���V4����=��{DX=�V%���=��<d��=-��=���=f�<���p��=�0;��'<z�>z�a��h�����>��>�fC>v���c��L��;��<���B�:c�>�C�o"�<Љ*>�;�=S�=&e���{=��F=�[�����{�y:��b=$�=� �݋��sQ�"�F��M=i��<!�ռ5uӽt�\>�Wl�Nw�=z��=�ְ=+n彵Wj=a�L=5,e�ꊄ�>����S>k'�;R�<	3���o�#Z）��e(����l<�{�&�=�Ƃ<�q��/�M<�>ؼ�=!�ƽ~�<֔��'�=jȂ��jk>�g�<u
�= �l�����GJ�=x׼<����hC=@ɹ��E�hj�q��;/Y�����r=���=�ܱ<���=��f��n>ǽ?�|�$����7h<�?�<�m��=/q��&潘�W<�l�[��<����=�#�7��� =�F�?e�;a�R>����=�Wf=��h�# 1:�L�2~��4�v<��=y����q�<9͹<[5���栽��U=�
���]C=zq�^��aL�<�z��ÑҼd�[�;Q`>T�(=�|�����l�>qK��Em=3ʚ<]�&>]V<<�ͼ���v�|</���b=c�ܼ�#�=[�=�m����I�A�+R�="�伺T�<�J=E7=e�m=�B�<6_Z��A�ɿ���f�=%w�4�����"��O�=���=cB=�Z�|_ܽ_�g=��-=�`���D�PW��h���bz��<�!=%���~�=&_��$�=�� >7�o�=��<5&�^s��'�Gf����=�I=i�y���Y������]�: �$>t��ͧ�<��d�̽C�<`�C�0=���=6�>��;�3��\����=�q�<K�ʼ�佣�m��fԽ Τ��p���Fҽ}�����<��=�:���1�:ݦ�vn�=�Ǩ���f=1G�=˙!�>�=T9=~�w�p2�-ͽ�T�<���5���l�8�{�{=��=*��:	������=g��=J�=	e�<��Լ�8�N�0�!w�=���:F�<�b��(�>��x>�;�,>����{wF<�ޡ<p_��uy��R=�5W=1�<�漒�<�=tu�@f���
������=��E<>�=�Qc=�܇=:������ϭ�OE<��;�u\�������=͊r��P����;4\��4>���,���$�QQ�D	�=�Pӽ�(��L>=����*=��Ld9=��{<�G�<�����NE��Z������b`P��}�<7��=��<������L=����&�<�%3�ϐ����=�^�=���<��/=�݃=GJս{��=H��=����a��ZƷ=g�>����4>�r=#���Rֻ��~����!�<'���ؽ|���:�=�=g���K��%P��^?�=���V�<��t��蘽��=|<�}>��L=�"V<u��A�=�@�� <�޻�>#���0=������:-(�=����J7������9>Պ�ׄ㽪���`�мvOP=M�ɽ�& >W�� >��\>n�;J����1=e���s��(I�=@�=	�C=M������J�+��<�ӟ&��X'��\=V'�S�n�a�N��<����>%�<|^=�Q@=�u½�/��ꆁ<g��<;탽籕��s^���-=��A=s�,�)q3=%=O����=�T��t> �Ժ�Y&;Mn�<v�"=�־���<�]Z�^<T���= 6=�O�:A��)<U0^:�c|=�*�;�W)�pq�V0��:��㽝d��&����y�=�ҹ=�r�=�'�=[;=�7�<��*;��i�(=u�l<%��#��`�;�W�;vR�=�F�<�6�<G�f�v�d�	�e�=�d<������<����j��=����;={�I��N����i�<���'��.��f��ֽ�4�<��<��=�^�=E|F�Ԯ�f��"N�<�G=vD�h=֗">�y�<�R�Oo5<A�һ�ᆼ���� =��>������żI�o>mٙ�<:�<iM=v˼��;M�p=U�����5C������m�%LH=��ͼT���6ֽʲ7�����V�=�����=��>7��=�n�q)�=U���א�h�ýՑ�;'$=�'��J[<�����k��9>"0��^�SB�<t<�:��@O=5J���\�=��<]J>C��U=	=w�"�ʔ�=�]m=��:�dϋ�-�ѻ�<j=�<�N�K��=�$>�����Ȁ�W�q=M�Խ�Ϗ=ak�Gw�=\��=�/�e-��a<>�,3�I,�= !μ\N�=����b*
<?�=Jj+<��=)
=40���e�G�=����!>�[+=�k>����De�=�=f���5��vG����>vy{���I����NzE��&�X��?ٔ<m�<)2�=�Њ<
�=y���̼I�R=7i�=��>��v1=��x�n[�=�^޼o��=�x���#=Y�9=]g�=�aJ���켉������=%�`�pO;��=.����<|��<xm
>N�R����	�E��.�<�NL>19��� ��==3�B��g�1[4=�����t,��f��_(=ČR=Az��g���>�b���<Ɖ��>���=�b<᫹�?�_=􎊼<�+=Cн�����u���=���!���c�<<>@�=�s`=�� ��aS=t�_� �Z<f��gtQ=���zb�=h�4<B���G\8��v&<�����=>`W�=��x=Ed�Nd=K�<�O^=�V4=�������;ಛ���/>�p�=&#ڽ�><	`M��[=��<��=��>b�>���T>;�'w�\-��0����<���P�����Ttû�l>lVu���=��=�w �lཻ��>�5�=�uQ��z�=@P>��=}<4��<Y�;�:��,�T��i�<���=7ߋ����pϽ�=�b�ۙ�<]�L�ܫ�E�"���=�D�����=���=�G�=~�d�T��=8�4����<���=8�= �8>H��=�g���8�=/���䕤=E�����:Έ=2���Ľ�ݰ6�F����۸�״=�.��n>{P�=D���yI�=JB���v�g�»�����"�:��������[=�мВ�=G��<I/�=�h��^���V1=���<Z%�	����^=s =L��=۸����p�����F
����C��ɽ�i=%��=0�=<N���=9k=$;*<���=����t���.�s�e��LT=h������dZ��M���o�>��'�oHG���ܽR�=�.ѽ�E=�=��Y=��<If>���=D;��7���ؽW>���V��sN����=C�̎o=Vә�GE)�<��̢
�J�*<�r���`{<�b?=v�������t|�<���=���ܞX>�M�=��|=��<n�ܼ�Mi=2����(>j��O=�Յ<�?�<���<�$�Դ��̪ >������=:�<�̗<��<5�b<a�U�gnb���1	��[wC�O�2�ڡ�=\����=A�=y��<�=>�1=�W����v����=���=���Ȑ�����>� ���<�f�S=NO�= ��^ʸ�[�ἁ�>>P|�7����O=��=�	�<�մ<�z������/���`_+=������=ϼ��Խ90���<�=;a��!!�=��K=+h��"�<M����-���TZ�M����ԩ=���on�s���[z�"%�</�B���q�"�n%���½���e�#��=�S��fM=0D&��Md�B��]!�����ǽ��=�w�=���g��<E�C�"�����=��d=�=��L~��c�;�=0�Y�ξ�<Q%R=
�8��^�=n�x=ϭ�<����g�<zg�=X�=�;����%=.ef�����������Ix=)�<[�=o�=O���D>�y(��pT;�f&=��"=k&= �=�>W*��	�k=���A=�&���5>*M=@hg=Ν=�t�U��6�E�Y�>�f�����Af;�<亂۞��$>����7�=��Y=��<���e�>���=��>�z>��ս��T���(=���+t�<�>�/�<Λ�<:������B=6Y7� 4e�ǒ����<�8=D9;_��=���=�!�� =A&�=�/�٠�=�Y&>��ɼLz�=Z��<�7�G=9��1=�;S<�!>�5̽�K�����<�}>R��bҒ��Y���kҼܭ����<�Ұ=�ː<��@>*� �g��F��{?�3�u���C=L��<��:<�7<���^M�wuE���ݻmy�QW˺5�=]��=r&F=����Ǿ<i)�=!<:<
6���ټ�kZ<S���9��>��</m��û�5��l��6�s���)����=f��=����򼔣h=��<Kr=C`�T�J��=�n+�#�*𠽮���߅=��ż@F��3>�=v����.5��>l�I��P3���=KSa>��E�8,=F�o��ӽE�j�o����[=Jk"=`���Խ�aT����=�Ȍ�HI��f��<a��=}��=h忻H7���%�"I,: [�=�¼H/'�:n!��C<OV�%�|=u���c�=�%=�6=tm6�o��9����K=�@R=�̀=��i�6����tZ>`�$=8+�=���n&���<D���Z��Y=�A =6W����<91�O,мb�x>��+=g�9�y�:�C!=���jX=k�m���=���<�)Q����<�<����=�sG�)��=���=�(5�'�6����=�G�;85���
����=-�Y��[¼F�=��ϽPK&�й+=��<�l��8e�=��5@��a>��0>��=�(��:}������>ǻ���&0�9޼4	�a����K�y<TG�=�q�=��ļ~���ջT�<_�={��<g��=0��x���u߽:'�<fz<��<׏Z=�Vn<Ź� ��,q�=:��=C������%L
>]�<Z3�=��=�ͯ=Ԋ�;�s��L��m�o�����2>E��sV�`r���m=�l<�	��:����!<�dd�����O�����=���;�&����0��7>�O=����;��>�R����j�B����<� =+��7��=�0%=1���Ǘܼ�Х=x�I*����< �_=N}ٽ��=6t�=]���n�9�e;V�D��֯l���<��=�++=��<�k2� 3�gH��3����>=6�2��.�7�;l����C1<��^����<�M�=��<b��=�����-<��B��;<��<�����.�=���q4_�"9Y>����9O:k�9=��A�ٚ�=���[�=y��=��X�*�Fᔼ����=�4q���=k��9�������=nH=���<3�<g�E=��=���=G����H�=��">�Xͽ�q�J���I{��
G�k�������'��k,�W%�ٕ�<5�>��=��
���1���`��=#c�e��R��H5��(�> �p=Z��= я<�K�=�=RVP��8 ���]�8_Ž��=��ּ4��=Y۽���{��Ȗ<=y���=�;H�>�ڼ̕<Ck�=+!�<���=�.>�����<���=jBX<��&>�L[��'�=��>��ʽ�w�=y�=k� ��ԻQ�<�U6��V��ϙ<7�W=��ּK�=l��<�~=@/R��vֽ\D���6���(�=N�B������h�� ^'��*���0I�+�M=uh��`��g5h���"���U�!z�"�	�Xm7>+̮�K��@�мE޳�g�<T- >s�޼8���8�x��.{�V�-��ټ��l=�轳U=�c'��8�=W��<i�;>̙�= .������܆�<U���o�=\��S]=��=#��=�+�ț�=0��������P�<�re=,�5>3X�=[�����������=Z��H�,�S�/=Yd�����Q.���;�!>�$��=~��
8=�=ci���= r�:/Խ:)5��נ<==���=�;���*/���j���p��zA=�h=��<Z'���f>/$��hռ��'���6���k���,�2>(I=���uA׽)FƼ�Rм*���b�=�j���S�<�[��4� ��	'�ݜ=�ɋ��^ؼYS�=m��=����N<��_�񁋽W����-�|?�S�d�F"=;c�<�7=D8J���=���=��==�����c�˻Y%<񸞼�y=�x�;%->M�f=L�=� �=S[=������@�(8�=\����$]>��)��Q=�<t�X��D=��n=ri=V.�=H�O=7#�=!B�9���;�m=�y��r=ؠ���9�����&H��F>lD"�v�>�-��;v�h��=4�=���<��������1�"n��6�/=P�=�ӼD�=�8��(�<H�=�Y���J��{��=�����Y� f=�q�b�}=O��=:�ټ��\<:�u���F>�0>n��<�E����=�Z3�]�=������<3>��T=i�����	�v�=Ҽ��wNL>Q> �~�(}ѼC��<��h=[���?Ѽ֒ �����g���4=��&=:B�<!Vh=�½q�0��=ژ4>[m�����&8<�V��\��|��ˮ���Q���2"�P��:iC�=��M;䍕<�*�=������<W2�=!1e=�f{����=p1ֽFS�=P������j� �Gbn��¼�)=aA=v�>�.�<6���N�ݼ�O<R�l=S[�����=8+��*6==k�:I5��Z�E�L%�������{��:7��a�=iu	����=��ҽ� >ĩ��l�ؽf��M���"ͽ��콧\ʻ5(H=��<�-�����<Oc��7�F�˽'(-��K>B����<���<�ث=��9;Ӹ�2�>�_)<D�<�k%�1������;l�A=QB=�>Q=v�@>�M2��jt��z��,�l:�`<��ġ���h=���`mT=\a���j�=�=�P�rA=O�(��d�=���u����Q�k�6��;��e>N�ڽ�Ϻ;//;ٶ�<�`��� ۼJT�!�=��=%����=%qx=���=�#R<��<aż�9��J!�PT����O��<qs>�V����D�,��=a"�=T�N�Zd�i=�<���kR�<Q��l�<w{�=�E���� >�Լ_�=nW�$%��+��k%�;�_=��Ι="��<ۻVX��8�=Kֽ��=�`
=sJ����=�l��A巽�">XJսޛ�=m��=��5�eXýo����T��4���='u&��
=:�=�$Y��׃��Y�߳:�>���=YHE��Ba<�O�=��4�5�=U���&m=��{=,὞�<���<���=����N��;�g�����Eb�=����0>�p=S=�<N~^=�A���d>ڪ��*ռmB}�c���<ü�7Y=|^��w�G=��(�ր��dȬ�e�=�;���������������d.�a9�<��o<�W<��	�*���v-�;l@�F,)�ت�;hN�<&��=�3���,��_<Q=�;��}���V�=e�=�=|jo=i�u�)">˗<6�O�@����4!���w>=�S�<_��=���=�b��z>�������63F>W����R=Ϧs=q˽�3�=z��<��6<'��=�+=�mp���=��<�'�I!�=X��=]�=a��H��m�*����;��N�c,=AӽQ�>�U�=��^=	0׽��p��W��!=㮖<^�;,=�)���lt=}/)�t���8#�;���='+=�9o�<	�=3���� ���<�H�J7�=�[u=
�*�e��<����{Щ<9��=��<�$����=R�K�4>�>I=�&�=c�_���L<�"O�HA$=����6)<��=EJӽ�d;�{�=�  ;C�=P'�=�q�=� �<�p��I�=�e<W��<x���2(���-�<㹽���n�=8)d�%p^�(#�A=��=��=�f�����X>�Tɽ'\�� �=}F=E�ͼJ@�%r��/L��ZAN�I�=N)z=�dc=�AP�8�B=Ɩ�]��<ָ
>t��<+B->o=�ꔽ�Z�=�S��n�=��ԽSS���>��#��B��wb(<΅�;�Fƽ{���B�<��.��ն&����2���6U=J�2��E< ؍�Q�0�e�$�K-�<y&=�[>��ۻ�)'<�P==y���B<q�>�XJ����=���9AG=n�}=�^˽�{ۼ�h!=��I��y=Q����;M%��W�׼l�>ـh=Z� =�qK��J��}/�at��	8�:(���
�=)���'�W&
��,r=���==�=2U�3���lcҼ�K�=9`I��}<��T>����=�)�����#��=����;���'�>�G�Ἓn�u��=�g��՛>�Dɽa$�3%'>���=��Z=MF�8�!=�V�=�n���i�=��&>�=*�D;	;%�Fk�޷�=\�=Ӑ̽D�>��;d@���x��ҡ<�e���=O�m� @�B�Ľ&+�:�脽Qͼb
=gW}�_�3���߻+D�5�<r=R�7;�@;�֭��9��=}�����B;�{�%�����=R�C��5�=��;�5>���=}��W<�v��=��;�h�A>����I>��Ǽ_�;�<!�	�>�K�=-��=4¨�N�m�d�^���Ӽ�,5�o��=�����H�̷@>�G�=�G���x>W������~����>�Q�=N��*��=�U���!>�F�qSx�Bݡ=v�=�!<AĻ��1�}��<Dv�v���<Cؽv��F޽ ?=?�պ�iZ�k��=6O-�4��t�=^��=�2>�ۼa����ه�;�U=�����H�����6=֋A�~Ů=��&=�9t<��=o`9�i>�ӡ=�}�D���1�����=T�~=R��ڨ���x>�`��@W�E揽�ڿ�+
���>=������y�<HP=p��=���<�"�<V	9�nq��*��ڙ��/�=����@׼�½?~�ܘ<�#*����=5%>fs�=]�A=8��ķ�=��=2�I<�>���K��6i�$K�<���=x�*>)ϼ���=����u=�,�<挺�OF��v��=��@�ԍ�:�"=�ݽUq=�-�=3z��_���ד��8�<G">:큽��ͽF��.⽽{2>���v�X=KY���O=ja[9�O�=�HV����� ^��P��K��=.m�=�jW<(�.����=P�u���<K��D��<Q�=�A�<GX��f�<%j�<�4s=\�=wX�����=lOd��˽�Ŗ="^I���A=2��<����K�=�a<6S�<{´���>��h��5���=G
��$��+�)�\X���������=W��=��m;�AL�eĔ�l��=�b=�z�=9Z� ��5�z/+���5=w+u=V��� _w��/�=uou�^�=�>A�=���a� ��� ��H�n=��=�d�\=Y�soF<���Ի;����2�<K�=hg��V���"������ ���������~�f>�x����#��Ҽ� ��7�`�O��=i{|��Rs=FC=!�<�1�@9=J��i<�yB�[��=|�<9A�<2���� �<���=&�>}g=��|=V<���t=��ټ�qͽ��o<���<�ϼ�.=���=7�><u�0A�����<��ν�z�<s�ҽW)D�ܦx��(޼�SV���b=�:�<��<�Uv=�/�=�;�y��G�'����"�=i��~J>��<H&P�D��Hf�|v6��9�b��=c�3>�Tݽ�c�=B"�=dt<r�=�G�%j?=�!���F;���=�e��W�W>�����½�^=f��;�:�=��0=�.���&�E;�=�í��w
��%<�ȡ<���<(�><��=%�= ,��	��;���0gм���<�x=��&��<�g�=��3�J�����꽛���kV1;nW�<J��<ˆ>�G�=RR �E�7=-G��;>.R�=O��<�ּx9���1=��;�3z=�
 >�����V����< ���i$<�W�<	P=Q6>�K�<c�"��:�;%�(>G���%�;|=L��R>>��Y�G' �V�W��,;=��<h��=�p<�C9��k=���Q*�=`����=W�'�-TK�E~<�s	=�)��\��{eU=���<�@�<�"!>M�<ɽ>w'�Y{�<q;�H^>0����:=gI)>�р�t��=��=g�#�o�<vI>���=xbk��2=�����>��=�O��� ,>8݀=��=�����Bw=@7l=w!��ν=������=[��=�5�����r�����l9O��0!>ىǼT��<6�4=�R��oM�<j8t��b8��v��U�#�"���i���&�^�Y�JA�=o�!=^\=+6�<���^�y��nN�ˣu����\�/��<�T>D��=J8>=��*=����Ht�<��>��6=�"y=έ����h��l�$�*���\�s=>�mh�**=;qY��,�=���pz�H�ýo�=r憽]��<x�R<b)�<�7�=��i=F���T�=�="�|bd��=��{���=44<��;�k;>�q0��Y=�7=vʵ��m�W �<�v�=u?��i=tV�=s=����A <-��=���=	�X��p�	#�==( ��r ���\���R�.MH;?�����:H�	<=Ti<�J��Z���*e��z<��4�U#�<�}��:��<�9�=<�=���<Fj*���P���,>2��=�ƕ=�g=BQ>�Z���뽔�½��=m��<�p?�&�u佸L�=l����=xq4=�����d�;gci<��g=��%�=T�=���=w�$��ы=Y�=~��=�X>�/�8̽��������RQ_�/�ͽ����R+�q�8�ZN.=���s�<�: �Yق��"�<֛=���="#x=i¼9��z��<A���r��_���g�=.��<$ �4���{8���Ž��>~�>=��=��	��q=}�*��Fڼ@R=���<�Eܽz`v=>ܫ=�jM�P����<�2V=����I�W�=��B>���%$>�L"����=�i��PBA=�`=F"\����=!�>�)ڦ=�8��:@��P^�=2�{�8��=�cR<ͻ���5
��l�=M.�$[9����<sh<	���?�������/�=�h��QJJ=Mx��I%)�m0�M��Gō=�c��L�����*=jQa��8�<��=?߼��	<��t�=̞��J=D���N7w=?�=�]4���<=�:=�\ʽp�՗�E��p�[�=����*<oI�=Ť=�o/>�">'|�;�Gi�5�>3:>�%m���j��,d��Xo=��{=sY�<|��
9,= 8=��W=���=�N���7��l�+���7=�t/>Kյ�K��=�U>C�&	>o9g>������<�=�=�=�к��O>��=VW��G�ﯽ�i�����<0�t� �œ=v�TQ=<ȇ��z=�[>H�ѽ-���'=�&Y�p�F���!=���=�n�<�\Һ�R= ->��=��=����9ַ�p4�=�~�=���g����y�=q<����X�<�����<�J
=�W�=E"�;7�,�=�ѽ�h�=le=��Vm=�<"��=#	W���@<Y��z$��k����=��<����P���o�7�~���=Su��!@�<�|k<�;�<��=ژ�����=�W�Ś��,,�w3Z=HM=�B�M�!=���<��L=Q�ͽ�>�=K#���C.=���<v�=l�E<���<�u=�� ��n>�����q�&սwq��cg;����e=朝=�<?<>M��=r=Am�<�1�=��.�2��<l���z�f�R@a<h޹=�=:�輡�����3:�� �=�~�=�Tռ!���H�K�!<���=��%=�L����>�2�R���C:x���漸���z�%=���\5=A�&;������8�G�Y�5��<;��-��x�7��RܽbnC=��>ja��P�H�;
�=0j�Sl��oZ.= ӌ;V�>}�;�C2=���=X�=w5ʽK�h�k7&����=�
�;G6	=ǰ6=��<"��=�&=S���b�W���S�#f�&�����<��!�_�=�ܽhJ㽵e>� 3��R�:���¿���7>���<�p=�9<��<��=��c� ,�=n�5�нO�;> ;����6>�����|=s\�=�,R��q�D	
��b��:�|>k��=C���o����?��*żP�=yD�=R��=7Ȅ��@>W�@��2���i߽�#��#��=I�=Ϸ2=���=����S����x�n=[Mv=�
����=)�v�DI���`R�=Z�S�h�X=�U<ܽ�A)� j@���r�p�1�>2���ߚ<�.\<��g<�f<c� ���<�[�)�ս��Ͻ8�= �=��=�!�=&
��,�;�Wr�^C��'�ǈ�;!��=�9� �!=�e�!�7�Ҿ���`������=֠�=�h �%&>_{�=*L�=�ZV=
��;*����ݽ� I�}�K�'��=�n=���=��F=~g4��s�=V?>�C>x��=dv<�-뻵eл�s=;�P�ݼ����	~�H�7�KQ�=�<�=hɾ=ڡ�<;�j=V��ZY���q#�E�!=+�:<�T�m�w=�F�<����\>L�ǽ�S==e<�"=�7c:���<p
>�����Z=΢l�����	�=�W�;�k</5 >��M��6
�=�=�r=Qg⽕ݟ��x<Bj�=��U>깽@*��)�=��<�iQ���HG0����=H�=[���)����+Ie��h=Rj��O��<�� �J��='���y���/�@|�=�'>�;t;~��r���%"=} ��g';=�y�q�s=�� =v}=�œ��½̷��:�2���@=к=�B��½,��=<B=��=�/%����=�J[��w�=�"�=t)��䯽m]���G=J�>K�<�|���=�ec�� =q*����P�<�2�K���..��c�<'F��, =ӑ{=��ܽ�쒽�s=�0O��_�u��������[�<WxU�ݠ����0=ܴ�=��=��K>���=��>=�<n��<�*սh�㽒"]��9��7�;��4�;��a=-�v=Qw�����l�j̘�X�>�.�m�=�=�Ѽ<#��<N�->�=f���=�T�=�!���8�=�Y�<5Fi����=��������g>L���ʘ<���<���<�=�=�t�E��=�!Ž~����wh�
�j�w��=���=M>���;�{�=  J�h��;�:��H��<fμ��,����="])����� �"=b�>>����߉����>�8$=���<�`C=��=���^l=�5�������� >�傽B�'=�1%�3���>V9'���5� Y��/J��C'=�Ғ���<|=6�F���=T}����=ۤP�&č<\v录E��WtK��SI�H"�=�׽���<���<bC>n� >��4��m=?��<�C���m=0��#?>A�.����<"�q=��>�ܒ=U��<�U<+%>�z->i�l=���;��G��C1�� �;���=B���w��<'R�I.<���=����2U��o�F*V�?��<|�¼���<=h�E�=4����F�}�<Z����ƭ=�k��2YּQl�=4h��.7��L���̱="x���w�;���=Ǚ��3�˼n<{����<���<�d�=@�>	��$�`= �ݽ	&���<<�끽���<K\m��@>�y�=��m=Zf�=��bս=fD����=fwܽ�)��&	t�B�~<&2��>i<���&�3=-�3=����c�x�.>�ț;6;�%�<-D�;�E�;�t�=z�����O��^�=�ǼOT��]�<��C�X��=�����r=�=I-�����+C$��T�;�D½ZI=jl:=�O�=	M��֪�G Ľ7�˽z�J��=�
S==�
���=8�@=	��<�۸�~�� �=4R	= �!��C�;� <�(W<=Nr��S��<��G�2�=2p_������<���V?��^D��sE=��:r�>:-��y`�=B-^;(�%�=x���^=f�><$�н\����h�噻��>"���47�Z�V=C��=j�!>��d<�쏼밳�h�t��+���q�|��=��<�tQ=���kѻ��X=Vz�/컽�E>
��=c=��st�<?CM=������;;; 湻C�����<��IC�6mo��IF�A@����>��H��#=��ĽGh=��<�њ�d��3�=`��<l��<�=Ba*=r�/<�ʻ1<��=�/>���=�>�
�=�ȕ��i> =@>�ҁ<޿J��ף��tX��獽��L��=4='\=j>jr�=�Ľ��k�q)���<i���<X��j.�w�T�N"�Mx�=3���ʠ�=x�>8vA�f֗����<���paI=\�F<�'�:�����=�n:�}rV��uh�R}�=� =�>*�W��<�p;+?�;��;'�v=t�Z=F��'�=��<��9=�5�=@;�=mŞ��{����z�-�=C����&�D�M=b��=�yJ>�(��'�����K輱��=� >���<�kH=���=q�j�;)%������E=��C���Q��0�}�p=�>f?=du�����=cd����ý?�>��ǿ;�0�	�=�F+>�����M>������=�D:��s�=�;�&�Ck<� &>x6�=9���w�	e��3�gء�B�u���>��=��a��a={r=NI=#
=�o�;8i�Gd���{7����=i%�=G�۽��ٽ�=�����=�N>�lK=�i��ct=]x�Z�,=�/�d�>�0n�=n�Y�d��7B���i=J�=�r��x �W![��ۼ���<�vm:s	�=�w�=���=�ص���-��hֽA�>����D���~=ԙ�=�o�=vm�<;�����=�
>�L������:<4��݅��ߞ��p�;¢=~I��僆<0��=��0>��=����f�<���F��=���]>��.�=���=�}#��Ӂ�c��H��=���=��=@� ��%�����<Fb=Z� �x���&���j�s�� =c��=7��==t�=�d8��6N<�aн��}<����x:�:���f����n���;;*/-���
=:��=8�L=bQ=�� =�M���ެ���=��˽W�/=�/>
��<��ݩ=� �=��;��]=2K�=k���0�x��=\i���h׺���;�L���R�==���5�A�v���r������펽r����w=��=�<�ƽ�t>�n�����F��K�.�$=	i�=��=�����w=H�=��X=�g=��#=w�=͘\=o�=���=��=fM��<Qh����'o4<8��<0�$�80��ț4=}���%j����s�F�=o�l=n��<�#�= �<�X��n�����<���p ��L��=S �;���%�a<�!��M����=�u8�D"�<�|�<1&�9r=�_�=p���n��
�^E`=�B=�<��`=R��i���z䄽�w�=ߑ�=�X�= /(�2:|>m�k�x[o����<�����2�=��<9g�=���T7���<�����:�̛=�½�fԼgA��kȞ<�Y���{��\�=�i����;s�߽~Q��C�=�>)v�=��v��>�04�ko��vW�=��={f>�/���=V�8>��	��뵽0��=�1��k�{�RU�;p���v@=��ٽ[W9����D�����=����z�nY�=�����Ai=1��=���6G��x����W�<�ū<	>�]�T)l=7�=�Ic��������9n���\m;_�=+���;	�=�x�='j�=������zr�=KI�<D���5:�{�=�%���И<م���$ý�!�=�XѼ���w�C�8н~4�=c%�`q?=��Ž8p���=��b;���<������;��=������"�Ζ�=�-=V��X�~<�Y<�� >GX'�����zsL�l�=47�=�꒼���=gy��㑼�����>�Wk=�+�JA=���;
�<<@@Ἢ�ɻ,?����l�XT�=���=X�<��򽡒�_6����:�Id=_��=��Q�B�;Ј���2�L{�<x����)w�I�=�=7�|=�ֽ��=����:��5�?0罃�����G�Z*�<}T�*�����t�������B�Ľ� =�{�=m��;R	�;�}�h��fp=<�	�&�j��a�=5�n=�`L�ؖ)==�۽E??�c?	=��L���"�[�̽�ꃻ�-�=�[4>��L����=���촼W��=Fn��JG�;����9�֘\>z���m?>7)�;���<JO��V�= L�N����4C=⛼��S�=�ȼY��<�=��>ɷ+�fP��O�=�U=t�B<�;3��=���YD��'^�=�=��2;������񽭽��)>_l���{�C�ս���U;٪�<QE��J�x<��j=�V-�2_��v��.Q��o�=�W��fޅ:���=�쯼�੼�]t=���ǽm� >Z��P�����z�8�`;�:�<��Q���,��M�=v�$=���h�=��_�,�2=O���">)+J=�z�=�Ƽp1+��3�9o~�_�P>����K=��Q=u�G���=g>�H< ~�=_K�=V��=�̽�ʥ�@�����x=�M�=���=�K�<�B�Ĥ�<�=0����!=m_�=X�=j��J�q6>����D.<2;�Hp���}�2�;�w�2] =N��=�H>8D�=��L� ��\���(z=5�0><*���3�[<]�<��=��=�������W�<]h�=v�<��=bq̼^c��.Y~�E�<7>�/��E�����Lý!E�<(:��_=�!�=�g�?����]=d�=��'>�����de�T�V�x<ِ�<T�+<Z*>os׼翏�TV;����}�<O6��蜽��l�P�ý��=$����=7c���Ƚt4��	��$�k�jj����<~+ӽ��z����=-/1=!�'� =ϻH=�6>ܪ�HU�;�Yp� ^+��y*�ͬ�=�G��n�;3WC>��üX[*=t:#��{��k<G>`�U}��6j�<�/=���ր���	���o=���������;��Ҽ�^�K��=�-=&�<˺=˵	�|>\>Y�����\r���tǽM�o��y�=mIb=���<%=�lm�'J�<����vż�y�=?�>D.�=�%�~A>�Q*>�@�/����=#�3��[��V�=x$=M��^>�q�=~�#�0������S�	�D <H��=4����	��wq=���=m� <ë�<ϛu=�T张V�<�`=�kh=�>�=A>���=�p�|I��j&=�=?���Nx=�꽼M�e�ӽ,I��]E��q��P4~=n��~��=p1����;����2 �t�� �~>�=M=�����V���R�s&�<{��:���^ۯ<��=���� U�����=�:�/�=pC�:��佄q��m3;������=*FV�n�ν6F�=h��ڔW����=}�r���=4�;��;�c=��f�#��<B=��з�<�C)="�[=cÅ=��=v�����=���=��3=�����Z �6R�<�W����H�:}A<��=�h��h�=����4�=d����=���=��d��4=�ŽX��1�>0���������P_�z5[=$�N��6�=�5=�J��L�<��;`I�;�K=(�F��Ͻx$��Q<�㠼	�ʽ1w�=y�}��-�=�ү������$���ܻ��̚�<\ҟ=�p��1eٽ�	5�;��<o{�=i���;*<��=I��=?ʚ�����}<n�l�W�4�s�=���e;�Ո�7fX��M��`�^�>���=�\G��`;`q�=�v��Ц=�=͸O��_<o�(�q�<=
�=����2�=`>=Yk���LJ���=��"��=
�v��=^Q����l=��P��<�v<~��~�=�c����<�_�=�����)����G�"��=����e����=���Q�$��=q_%��Ew�v���ν��K=�>cn|=lB����̽8ڇ��e��)�<{�1�	x[=l)�&39�O�=���=H�!�=ۼ�2����0>��=Z���1/��YY<�e>w-˽�3<E�*>��Խ��Q�C^>!J=��ڽ�R�=����*>��<0���&��pnC���>����jv=�&�=6���/�<N���/�=�B�=Ӡ��F�����=��<?����=*�7�Ú�<�(z=���93�=l�.���=�߇�`���@O=�}���=W?=�w۽(�0=�4��'*N=��=^�k=�%�e��U2�<d3�����,���GE�l����ѿ�:9���[�򅳽Jt����`<�;=|*}�Ex��g�	=w��=(o���?�<����"���WH>�<����v�Q
���t����F�=����D�<���<	�=4=���Y����<:ύ����<]6>�l<� 3>�;"�;����T���TȽ��E���I��= ڽ#սz�=޹�P�=M����C�6E�<���=��N>O�\=�{O�?�*;�"�d���9^����<4ʻ=�>a��C&���`=�uļ�$��P=����=1>v=�h��3M�<��"��]e=�;.�_»��H�K�=3�d��=�!JP<o�һ��=�	ٺ�s>��#����=�\>R�/��8O�2�%����=K]ҽ"�����4� u�=�\;�@3�='[/=t_�s�ҽ¶��Rp�~YW�K0��(�o����p�w�=Y#�<�3z�'��=x=��=:ۂ<�c�]��<�P��N ><�=�F�=��)�\�Z����=��b=%>s=i^^=���۵��#��R�0�ڼtW*�^7ݽ���70�/)ջzּ@������s�<�,E�̭�<v i=�*�=_�$��`�t����Fu=�:	>�x0� D��#��Z�(>��2;i�ػ8��<�Q���80�u� >jAB=>�	�<����ʷ=�W7��t���<�;2�>�c��ZŽr�={�>��;U�=��=�h=��ż��=r���->>�<N��<Vd�瓽�O,�����2��=�Ž��U>�xR<c�Ѽ��Y�O�*=�/��L[=s���k�=�Њ=�t��%�=~X��h��Q���*&�Z"=VS=FՎ�m
<R�>LW�=�2�5n�Y<!���3=�d�=��;�K=�	�8 �����$�X;?Z�<-�<;�^=ժ�=4ν�bG�_"=��;=hn\<���=��=���3E�z�=���<���{ǵ��Dg;��p�uh'�������O�
G��J��HF<�{�$*��E`�g�b�%~�����A�=��G>q��=�>��<+\?�j,y�����;;\�<4A/���[�=#�<
}ɼm�񻡊�=�6�=4����91�^����м�RT=f�<�-=���S���C�R>�%=���M�<=�2�:KA�=�u+=H�
�+�s������=Q�?>�Z=�<9�Y=�J�<~�-}�<���=�>��ƽ���<����;�?�=l�����x:��=���}"ɼ@y>��M;��.�=_��<���K���Pv���1<����*��"ٺ<�!�<>���bb9=K]E=U�-=�j���D�7�wy=�h�<�����!=d�6��t7=Y�ɼ0�:�&F�<^ټ��&=�T�=��=:2�<�
�^�=�.3>�~F��w_=ERݻ��S�%sƽ-m�<��&<[m�=2=F���f�NV�d�hA�=n[׽Ȼ�;�=n#=ٛ=�%�8d>�P�a¼q$=���=��=�ټ�j8=�?ʽ�e���>ԍ-=��4�C�>j���
���� �J�r���a=�=��>���>ݲ�=�y}=Yr�<hב>h�=��<f��^ �fU8>87=�.A�o�ɼ��.=�P>]��}O��ԻQFt�N|W�=���G�d���f;U0��_�O:c���^�ýĮ3<��=���<��Y=��;m�=fFƼ��=�=�=S�i�?=R\=WX>7�k<�W>��<����K�����Th����=�罸q�:u��W�~=/���������Z�Uu�ބ>n1g��w!=?ఽ��<��[����=��<<��<;oL;q��:1N�<gz==��½�O���=��<)�<�E]>�f׼����	��<���<��6�B��=�R�=?����i_��x��P�>�\��DD鼑����'��b����#<�N+�G���6w=�뛽�ѽ�]fQ�;��=����y���N=>�;=�彏�*>/=�{�=�d����o���c�v����"����=�]T=��?��?>`y�<B�z�^պ;ҧ�="p=�#�;LG>S��=k_�<F1��b�8�U��r]�?��=hv���=�^�1���-r�<�z�������be������I܂=���=Lw�<i�>?�Խ��#>��f�ղL<�%˽��
�t�=����Ұ���<�m»X>W�a�]s�����=���߲�=h��;�ǭ=��=N!<g[T<X_4= ?$>O�l��'?<`�O��d轏_����=�`=La����=7�=�Ę�/\��M�=�>�=waý�G<)���K꽟�߼@󭼪�H=��u�E�1� ڥ����=P�J=n��D)>`�k�� L=�?�������ﭽ��>=|-�=<��=��=�0�=H(�=H�Ż�8�=�St��۔�ܚ�=F�X�|� >/�Y;��`��"*=�B�c����:�=-���U�.>h�>�ܽ`�s�Y����,=V�=i�2��:��k��4��=������ס>�sa<��g=!?��o�`ѓ=ɿ>�m�=3��
V)�m������EI�GAD<y���� ���{=C9�=.��<��Ӡ�X��I�'=�����w�]�<�K8���=�Q���m�=�=w�|m�Z�e=�B�<� �=���ѓR=��ͼh��S�۽+�.=gl�<L"��>K��=��=����#[=3U�=�i�ٕ�=���Z/�=�D���ֽ�:��Q=�0>� l��U,�j3<d��t;�;b׼}�<;t[=Z�h��J�?��x=����v���ֺ�\�s>y>p�G=%>�>�	���0=�=�kT�l2>"|۽-���J����]����~
<s}A=`��=cİ=�a>=�S��ٜ<��>E�!�և=^]���?�<���<��">����Cs���z=�{T��{����=��v�1+��>��=���=b���E]���=�E?</ۗ=R>�#�=UlD��G��e���;�;V�v;m&c�9��=�Z1>��=)��=nz]<n�=�w[=�������_��5G.>���=N�<��6�zP�;�%=ȴ)��D&=0��=���!�M�a=
�N<ZE��	k=��o�(D#�N�|�������=�I�>����<�G�=�:�=� ?<Z���=+�T=����#=��;=n���$�=?#���hv<��t�M��w��u�v�=5�<H��=�t�;�����O�4�>�삽
Q�7�	��h=w�o<pD��!�=��>�S�<l&��f���H�=xz�:�O]���:#�����=)=�ܶ=`�<�q<Hے���<���0�t<n�m�籠=焽���<���=����)/���=��>D=-4�=��B��pF=�+��W4�<�q�=Bo=���p��R4
��+=ʩ�=d�>5k�=f�̽mR.=(ܠ��D>�]�"�F���>ּG=G�w=h�:�T�=�ע=>�>�n�D�z����q�ѽ���<i�=]�<X�,=��=�@�|>����=�3 >���=�_��üJ_ҼbR�=PÊ;ܖ���6Ž�3=���R>Z˼��<�D=(��=�/	�#0<��
�<������gؽ�g�=|��=?��=N��=T��=Uŧ=]�<|+�=_�n��=��=��^<ѽT=C��<�b�=��	����:��(<��3���r,�8c������k>�>!=Ӟv�-JP=���=~ ;>�?�<��=��Z�`�=�=ҫo�����.�F��M�<U+=@��p3<��]=����S���:Q�Z�4�}���=𭀾��=߯�=�Y�=��ս�~߼���=���i��|���W=�= $�������b�Up�<N���R�=?i=��z=�ن���>=8H;��*<0bz���x�'�1=髝=+8_>����.>�G`�@��<h�2>�lg�fI���G�;�=ǩQ�4���s�-=��ν�����L>��>�	2��Y��=ҽ���=�b:�u�<�|��h��=�^�= ��=�+.=P�=�> =��=P�0<1�=��ݼK	�<n\w���D��J��t	��B�=Z�"=�!�<_�p��Q����@�3YZ;�w�K�0�ER�=�=x=b�C����;��ܽ�+�;�Hz���;�V��76�+V���7�1ld�:ټ��<6
�=8�>�BT<�����+�d@/�ǲ.� �bnC�O/:=[j6=���::j���=n	�㭝<�+ ;�)�;�Y�;�eg<Ñ�������_%>���;8����e锼�U��u���{=�[��=��U;=!����=�!j:׼�=Ɗz=���=��g<(K)�&��;�4>n��<G��=��<q�=��=�h�=��"�[� >���Ȗ��z��>��=�G=K"�=ҵ|�8��<��V=�m�=��*>����>r<x}r�Mp(�cH�<.���8��ջq�3@�=A��=G��<#����j�s=.#��hF�����D=	ߛ���V������=�=�螽�k�:%h��E==@����=��>��j=�3C�LW���s�=Ϝн���=�2�=79'��Ur��@^����<�>�K����ڽ�+=8=�=��'��N�=�=!¼�=_.;�:=֣R��B;��=�A�o�X=qq;lU�=Dr���?<�/[�^�<���1= �{�Ľ6�=JZ=�sM=�9>q �=������<���¼���<��.=+�ƽ�Ş�<v�� J_=�"�"�=@j���O(>{�ݽ�ᄽ�����2=@�
>A>N��?�z=;�j=
 �:�<3�|�=I����O2�L�� �<M4��a^�F�>=��==��=��=�6���`M<����>+���<Y�������=Iɯ;r�L<��(���B>u�=
��=+���4�=6PD=]ߨ����==�x�:B]�<9p�=C���RN�=���n��=# >o<<�� ��.����@=�Q����dM�=Dw�;��=_���C>À�<I0{;+��;����EX=�(4=�׽b�<w��=��<���<���=�ъ���)���;�I�=�b��D#���Q3�u��<��4�c���=���
J�<�>�_�=���n]+=���=�� �����Ks<4�<+�9�x��=��#���=!5�=��B=A�@���py���D=��=X�˻��>�o��Z��=��Ļ#���ؠ� I>�~�
=y����f����<Y㠻�*;2�_�'$��}ֽ���<�o�=��><Ma$�L��([=V!k=��<�4��(d�=�Q�=�?����=�j2>	x���t~=�@I���=d֟���=�J=\>��>��鎽Cҍ<K�>�%�=�c�=��8��񑼑�>�Z=�a#=]�O=���<Ϛ�=sZ����=p�ҽ���<��𽠮o=��8��R�	-�<�]��K�<5Oӽ�b6<��2��R�����:��,��� =Ñ���c�����u*�p���8=Vp�=5�=�o0����=���=���<�� ��E=`�=�|=��=��t�M�4�T7�=�^�=4�>0:�=� g=�04��n%����bM��h%�:&ż�����^�=� =+��<�hؼ��o<�6.>�0k=h��=�����N>˒�=�䈽֫<�p���S=�H��p=�>�ޛ�Ӧ˽��;`[=�\$=M0��X�<�]����[<���3�-�r�:>~YP=��=�[�=2�T�:�B<î,��ah=�7�#�=�/��ż�>I�=�Y==a���!��TD<7cG�4GL<:��=15����"A4�1q����&=��ӽ��M�U��<��<] �U<ü�U>��*�$��<{�� +����H��צ=~l-=N�6<��K=�=	�n���	>OP=�񕽌���>�M=n�t<���=�:=��=��#�
)"���3>H�m��9h�yך����<�S>��ལ:���t����ٴ>=�%��0Ӊ��	��6�=���t�/=U�T=�=�ս���!z��<��I��<�=�,�.O >�
�VG>��<�D�=��N���"���	��>o@�<�3��r���>U��n0�=���<��>	!ּ@�>�u= PV�����h#=Lv���C=wJƼ�@d�pN��� � ��=�ʗ���=@�;��}=��q��`�m|�;q�g�baӽ���<�ȝ�݌���敼=������Q��=��P�=���/�qH=Q��=��=ӾY;*�սt=���<�}D<�Z���ue=��<��'=�Gz;RX�<��*��_ͺ��j��;f����P���9��l���=���=oF9��>�=$Tν�B��R���l=lœ��6ѽ&G�<&��=��=�����S��L^�Kf��`>D�->��;k��O�]=Wn�=�p��dk�� �=a�=����L��<�%�՝<H�v� \
�n�U=&u[=]�=�t߽�{n��\��:�==�o��E-��,N=`����zM�t�>w�)=�,7�P==%컄j|�*��:�iW��HJ=���=�s�<�6>�����޼�/:��^�6��<�1̻�}�<q��=��L�ʽ���L�.���=�ؽ��.>�B6>����=��L=�r�P�R�}�Z���Ѩ���G>���=�[=��3=�tƼB+
<����cŒ=���>�[�=�p+��ֽ����c���>.̼4 ѽ+/���/�=/e"=a�6�)V�j�D=�m���Q��f8�F7=��ٽ�2����=�i���>������w{=���i�< g����<u,ļX#�>D J�F��=�P��7\=��;O�߼Ez<��#=�q�<�j)>[���p=w	���a<��=�u�=�ۡ����<.���@�I�����>oO =�E�=���=9J����!bڼ��<֟�=�1=h>��U����[�;���<`Jɽi�ܽ?�$<DNN�|���E�=*��R>�Wh�[�>v/2�*"l�3穼D���:9��;��F��:<�2ἄ{�<��=X\=->?�B����=�F����=������<�3#���d�#>���g����)=�Tt<��"���<C&�s�½I(ʼ�3=IP¼K�?��]���}=W�k<xE&�6�E=ѫH<V<T��J=-���*c�l�>~l=:� =��� Q����=0�	��@_<rB)=�o�<8�=�	��{y�q�/=�";T�C=��K#�������T�|��<~\@�Ȇ<8��}��:�=嫽�j��<�?<�M"�P�<~;���52>.kf=�S���;���<63>,a4>�G��e]<)�=ľ�;0���J=D�=p�<.ٌ��8�<�T�_�Q��]h���=�0=>2��='*<Y��=m�=��f��<�^9>��P��e��=�81;�蜽:���͎=i`�/w�=<��0�4=ж#���q<��ս�=�ty='Wv=������<�AT���>K��(ӽD��<�|�fw����;��Ž�`W�@��=�=i]�<�f =q�;����=�8�=Jg���Ѽ�1z�N=w�w��'=TX����=��^���i�=l�D�W�z=u>>��6=W_7=�Kὧw�=���|�y����)[�;Ϋ�=+��Ʌ������⽑�_=��ȼ�������T<�w<zڗ=ؿ�=�������D�<�����<<%Wa;��>}�<���x���nH=ű��і�b�W=>��<�!�>���.���<��]�<Ct�=Jz9���=��>r�$����=t�g>"jK=�=�=����U@��b�<i#�B��1��=�K�=��K=vi=V��=)�x=�н� ���=x*�;)悽�ܪ=�H=�}�jj ��̭=�Cýg��=��>5_=�<��۽�Lq=~9�<��<".余���.�>�h�Q��=�6�V����:���=�� ��D_�֑=��c�]�>=�������WG=��ԽN���1L<��|=m�)=���=*Up=[ļ֛(=���<�����H���7=���;��d��y=H���W=	G4=P<�r���><CG��|<�_�=F�n=8��c4;�2������ �ڎP=���N�
�Ra��&2�=��&=>s&��EJ=�2��Y9W=$"=Dܜ=&���^p=[_8>�Q�;��=�,�=�4�=/���"�<��N���=ڬ�=5ټ���˯J��&�<[KI��X��4�:=rI#:���=���M�\��2;����2!]<����.�����1��a�=U�Jڝ���
�����;i<�J>9�P=�k>r��<G��=-���E0>��k=�ե�M�(��}�	=Z>꿥=�{A�&������<�����<3��^�\@�(����=����}i�<�`�����<I��=׳��T��fnU=�r�<eՄ�:~��{l���o�<���=
�2�9=��;�d��]A�E�޽�
���x=�gg�8�]����=�����E�=��=��߽=	�=�P�;�H�>�<=�S=�@�=�p/�Ϛa��|=X������<������&<��=�]��v�cн�\=*�Խ��<��u<tю��;�<�B=w�����f=���Q=���='Ȳ���3�,��=᤯�[�O}m:D$�=�+�=OD��ܱ���{����<�/��J@��`�&�ܪ�=����⼐�'��[��V>>[���q=U񹽖~>Yb=���=���=�o�=�s�����n'�=mp=)4�*�0��V���3>�z����=3*�<j>\F�=�#���u��Gup����JW���$<|�K=xmս4�j;�9Z�~���$Ϡ�mW�=W�ཷ=��;�.�=1��=_�O=����_D�h��d��:\w>燽6&�Y�<�.-�U�,��H#=���0y�����=
�>]ג<ȾG=z�<<lcؼ �� ~�;�L�=�4�<�s=Iu�=0P��G��=�򂽝5&��3��dL��34�<�m�=���=��P��=�]�< cǼ�����3�������]���d��ό=9�>���<y=aW��;3 =�����\>a�y�B�@��2��M��Zaͼ�GL=g�XG��Ŵ��Hʛ=l�b�X�����A�A�代<R=Ĳ�/������� ��/=\�*���;�i򼅌9�|=	��=��D<Q���6C=n�W<�W<��*����� 2���F����=���vL��G[���k��H�J�΂��%t<�!���)}<G�M�����oy����>=ӑ�	3��R�Ὅb_�q2?���D="��=B�;�Y�� �&�9^�;#���
_�Hƌ=��[=�"��X�<s0Y;7"���V���(�c�Q=SϢ�������=�)Ƽt��==�=����������萶<���=ňX<��:=q�d�/֑�[_/=(�=��j�L���}��==�̽(޷=�r?�C��<��=T���=�x�F[-���ֽb�d=���<"�����$=�o$������!�#��=�-�=�W=$��=�b��<���<�Q=��&=)�=<?=V�W���<�*��#�hU�=	�J�pE7�X�J�}Ԣ<,��=͉��j�H��^=\��<�F� ���:>�:��+�*=�X�;���~+o>�=ͽ����zf �%�+<w�T���>��=�
>8�>$��幽�o�R<����-�.>�N����;T\����=��=�. �! ��;^�<�,=|�/�p�A>��w�R}N���}��?
�Z2�<5��=O�)�+�#���=ft�<�Cm��l;��>ȁ����<���=�i���B>TO�<}\<Ĕ��a¼�p�=z�Ľ�<��=��=x���=K��=���=��=Ǽ<bٽq%,��͹<4��=��;�.>��'�w^(=H��=7V ���ƽa�F>y3N=�pݼVۼo�>	Ch<\�#=H>8���Ob�=ϙ>�C��ɗ=��i�Dp�<�=�U>�߼.P���>=�k�:$n�=�'�=i���7��Q4�ѣ��$�5<r�=M��<�5�;[|U��*B=M�<˕c=L�=<��<�DR=��A���=&/�=�n.��4�=�f����=��4>H�=�g���� 衽$���c��3W��P03��h���>G���|X����d<ƾ,���;|��=&��=eaS=�A�;
��콼���Ӛ�<��D�=*>��=' ݻ+�=�N��͂�"'~;pC=;��ü��>��c=��=�א;�:��[;>���=J`�;`iۼ�v#<�2=Q���=�ϓ������s-��c��(�=}��=��@�v	�<��8��=�#2<�+���{�G�n�LCS='?H=މ��Wƽ��=�ڙ=�E=[�;�%�=}��s����=x_d����<���=dk<Q�=ޟ�]�>*e"��g�=��A�B��<`쭽�=c�R�W|�=�g��s�_��"�u���,<f�V<w�<���<JDW��.�=���=���=PC+�²�=1�S�uLq�]$>ࣨ;E�<����=���]!=�1>E�ֻ��>�"˽�y�=G��=`XS={�Q=i����=~��=�G[=��=�����;F�0=E9�=_n>��9x�)=�*��Ӝ���<>iWi>�Ҟ��ͽ�y�	�G��c<pIn=�u�=�����N=����2��=�}��e�<D�>�,h>�&��%��R�>W �D���#���W���k<�k;��N��0>3�]=��^���"�C~>Q����k�1��x��=uK4�áǼ@b>���=�1:=.>��_��O-�����>�#�=f��=�L=c��V����ۼ˼�=F�������=�G!<����,p=��=��<��Y���<P��>�=}��S��X�o��:���=���<��=� =o\�����ڨ��cx<0��r�=��Ƽ ٽ��I=���U��U������a�=��>�d;a�]��eq=���=-�{�`%B<Z�T��E��<��A�:��,�<_����*>[9E���ä�<pO����b=�c!<�v�u���ɳ��t½ � �(�"�&�p29>���=�Bg=J�Q�+=�P�=1��8����T���z)>�A�����<��#ˌ=�PH�|q��;�=T�.<�2����=�������'{=^\��&=ٖ8�����X�ɼ0Y>�;=yN��&y８�?�T-<��.>��0���a�ӷ=� Լ���=�1�V��<^��;H�����j;̼>������K����=��=G�>as��毻���:��F��z�k�t��=�d�=� "��w�lm��I >A�j��nڽQ�e�s���(��;l��LQ=�ul��Jt=ª�v�<���0"U<�=�佽�.A=u��=��K;�:��H��y�)U��^;���;��=O��<�Y>K+{��\5�2�J���<	��� �=�]�=a�=Iwz<�^_�ѱ(=n�aQy���>t��v�%<ݟ�=J��=ڪ���@�<�1�=�Ɖ���=6W��H��j걽�d=5h�<�w>��=<kν���8P�=�x�=p��<��Z���b�t����=��<��߼��8=`�=k�;j��;^+!<˝��>#]��g>�(=�l�����v��qy�=��(=gY<&�ƽ�� �O�<�=>yl�;�=$%������+=�4��ų��cT�N�Q�	�{�3�N<9�c8�<:�>�\>�rI=9h(=�c���7==j >O�<��U�; >,�|���ü�q�<u�=���Y����qE>�-�wT�������=5�>�<eM�	�;�'�<��`��{.>j֪=��;���=̆Y=:�"���۽>��<�m�==����zｏ}���/�=]rW�ţ�<d��=/F=�һ���j=vѩ����'���v�=$�/=YI�=�'�=�ڧ=y$9��.��oO(�)�=���=J��;����ǵ<#���OW�3[>��
;�ْ���<�y�w5��A��;f�;���=�|
����;�	<�L�=�ɼ��C��4�\;�
��tj���G5=·���J��<"��x��b$��XǼG��=�t�=����/=�=���һ!>G�;�X�<�	�="��=� ��&�rā��<���н~��>s=�OP=��<4=�4Q����=�=�M�e���-�����=���z���7,����)>Ovҽ���V#�<Vϼ�%:=�=�wۼU�<�υ����<λ��+4D=R�<��'�|f1;� G=���=�cw<?�`=�;�<�p�;���L�x��Y=X�)�)<��9=���zc��K��]X��!��{���`"|�{S!>g	<����Ӆ�=�<��۽߶>�3���!�=|��d�=��2��c�=�K��f�]�!Ep=PS;t�A�]@>vU$<�V���+f=x󽖉>5?�<n}<� �=�>X=��-�ť=<�T���꼯G)�;����|�<e�>�QQ7�|o��ۊ�;��jXo=z���$
�Z:>�@��3�0>�v��W+>�����伤��=z��ື��c �&��=$�K�%Y�=h&=Pͬ���>��&>K�<��>�*����<�$ν���� 0<��/����F^�=MO�U!���^����g�>� m=T�w>e�Ѽ@n>��ڼ�fȻ����/��TӒ=���{�m�@=(����.>vv='�4���<����`,��4�=�&���=a
1>nC��k̑=��/���s=,�4��=��=w���7<|�=>����h��=x�t=ڀf>䲲����<��������H;��=�k��O�1>�;����e;ť<>�͋':�/=��ʼ=%�م�<|��>�<u��+(��*���ټ	�<�7�|H.=�����$>��������<�7@=�z�=�=p�;��=	ƕ�>i�=�Sr=m��� ����9=����C:��»�`�H"���*=�%J=���l�~.=$��=�=� ��=��@�p�=�>��T<qi������V�<��v;�*M=�lh����_n<�Gߘ�]��x?��4�=L�{;�)I��ֽ�>�Z����U<�J�=X=N�>v�����P;�i!=�3�v.R<>�<|��=T��<���=_-y����=z��#������<%�#=h�U>%~�G�>>i����=��=�'<]����8�<0�=���m�����'���r�=0j9��>Ri�<-"弄�>���=�YA=jb��7�=��ݽ���<��½�=ۿ,�{����=f�ռ��>���=N�����B�Df!>
��Z�>�|н/�ݽO|�=�Ǽ�ޗ=@�=-Uм�}=�&�='�=c��<�#z��a����b��b>=�>g���>�E�=��O�m��=����֪p��*�= p��4b�<���=��B=B����f�=������=(Ro<R|��%ݽ�0���=�+ڼr�=÷���=>�v=(),�H_B=�L���=�A0;kች�/��:�<:`=���<�&��|G��p����<�*ǽ���<\�H�r���8��W�<-S�=m�=�;�D��;v�^�;�GE=���=��=L>J�ɽ���k�ƺ�ǥ�~B�<��}=6�>=�F���M=D�����h���S&^=�f =���X�=�컘}&="�=���<L���qIk=��v�[�+=\qS��oa=�}����<
�>�Z��!-=
�5�5=2�*�E��:*�=h�6M�2�g��\�=-;1��ث;x�9T���"y�~>����q��M+<�ی����o>ܷ���0<3� >GJ=����ѾŻIVJ�"�=f�����C=�y=�ͻ�o$%=\�$��Ⱥ�U�>(�=��μ��E<�Ɔ�L{˽L��=����M߽ӊ:�d�M=,��=p ����ۜ�QJH�s�&���=�����8A��k��א<�Ն=۽���d�+W<��\��e���` �ZLi=m���S�<����Y��<J4���y��5��Cb=~*�;��4�%}���N=ԅ;>�=Y�>�߽Md��4�=���=u t=>ٗ�����I�.�����=!�;�����@�T��~�=�~퇾���=�.E<z�h��{�]e=��.�{;�;�g�	>��*>�6�;v�=����[����.=z�5��݃���F=̣�׬ �u�<�<<x�=��<	r��c�e�=�L>��W��=�k���y��M���=��z=��"����<�x��bl��^�'>���;�?�<��H;9S�=j�\=#��Kռ���=,P���cy<���=\�>���=��=%�����=�V�]�< qE=@�>_3H=3�E|����=�Ѥ<k�=�>=�b$=W���<��YԽO���E'<\ �;�)>�$G���vq���D;Q��=}< ��X=`�N����/>��<E�'�3L���i�=#n�=N�[�H.�<���/� =�2�=^ӵ=;gY=&�ݰm�=9���ܽ�N=����:���"�=���ju>��<�{彯9 =��=:��<���f.
�L֐==ӭ����=�����T���nd�=�y�;� >4�����=�*�<Fb���d�=J�ν�>�=%x>C�
>��x<��ļ8=�ӽ�D�<��=-Q�=`�ɽ:�X=�XF���˽��	�j�ͼ�R�����s*����<�!�����he&��B���w =n�=�b��Mi0=��H��݄=��b6=-��A�=���=5ҁ=~Bƽ`��l���D�����=�G=��l<}�9���=T^1<�c@=���;� =��ý��=�g�=�O��׽�O=lE
�S2.=,�> ලo}ּ��%���:<y=5橽\�=AGI�8���C�q=�E���߽W� �w:�����}	�=��ּ��m��@���Ҽ;�<�����.��a�V<c%L�+#� ?�08Y��!����9T	<���x��Ѐ�=�+=�J=d#>�9:���=��a=��ټ;:<��/�<9�d=����4�A�F%�%�=��y<��n=Ҳ�=Q�z�>=�ڝ�"H����=:Z��F�==��!�6�8�ּ��ʼ*\i����뀸=ب\:��ܲH���=���s��=�IG�A��=xe��<k��<�;�����v:�~�'�8ݬǽP���t����a=��=��
x=_��<��<���<��k��@2�j>���7}�;�	�=��uLr�ȍ��%˼���=�[#��3�o��=��O=yE=dX�<�ŧ<����/L<�C�=��E>B?R���}��k�[[�=���=d#>1��=EU򻁛�<����6N�;g@j��'�=}��=�������<t�<^w=x�<=��OEa=�C��^5�@�ۺ��i�{�ɽA�M�2�R=̼.���ʑ<��r<��ѽ�Si>��=��$���Y[��y�=�����Z>��ռ��=�X�=p��wٻ�U>�e��}-=�ψ<�s��S�>>��=��=Ѩ����t=�lڽn�̼߯�<��=�p=����=�~�=$F�G�Eͤ=I�`=�q>P���.�����RQ*����=�M=���=�O(<�&=g�=Rl2��iĽky`�cR���U߽�I<HPܽV>g
�9��=,�X�ޜ���0J�������&>
�	�o���m>݉�<[u�܏=��>RF#���Ӽ�����=�S���|J<�����T��{�%=���9��;?4=�r���r ��-�:Ґ�=���=*�=R�f�y�K����= ��=Pν�O]�q��=�J�=�>=n�G�D�c�ޕI=
G=u:<B��<���91*����=������<v@A=깔=x� =�f<�mg���*-����:��C=������a=F��<��=���=M<�1�=��9��]==O��:��<.\W�p��Ñ<�f�꽫�����=�l=0<��ӽ�>s٘= ���ܼ���=�,>�=<�΍=�>�=H���Kj�=�4�=h`�;Z5>�a���� ��v=֒=��;���0߳;�Խ����1W����-��Tk��C�=���'�=\�r=h�̽�D>�Q�<��8� :�=)ú#.g<l_z=${�=�,½�%;��?�<1�u��Z�����*o=�^>1 �=��+<��3=XB�<4�M<ݩ�<��=P'��K�� �	���<����� ����=rٰ=^X�=�O<=�e�-浽Z˫���=i�[�^q�)KF��)=�Z�=}��=��ݽ`��x:���l���^�8LW�������)=k|^�Fu�z8>7^�������>!�F�:��=��3=Y���G�>��>.�.�ٲ�%L=�f�F����Q	�B��= ��=�A��P�N�M=-龽�2�=7;<�Y`;5�=k����N���y�'ʘ��e��7�=���<��G=�O&����=�N=젲�Aɻ�i=�X7�skC>*��=����:�<ѵV�%�<Hq���R��ܟ���=��H;3��~��=#��=������i�=�����"�rD)=xݥ<���C<zAW>���=�8&����=F�LPҽ�'޽����׏=�h>��=��½���=���<lk2��D�*ҧ���ͻ�4W�
{>7���1	��ߊ�+R�=y���f=nG�=�Vռƍ���=��e�>l6<�ߗ< R�=����[�Ӽ��>�(q�,�G�3Ig����9[2#��H�`��������b=�S�=�z�Ԝ#;'�,��Ă��ɽ�c�J ��#���+=��Ľ!s��7S�=��]=�j�=�����<ǘ�<�u=�]��>=��߻i���É�=L�=�(=DJU��9>1��=���ED=�R컣-b��"v���>��8=�Q=LNm���=����b3=R�">��%>�ˣ��O�=�<w�<�9�=���s�~�_F�=��>�١=��"<+;>�w�T�+>��N<J��=S�Z=w��=4��Fv��-.��J���c��<��&<hs:�+PǽA�ݽ��U;l(=���ƌK�nS���aټ�q��wP�=!�=�E(>a=F٭=�=��j��3���f��=5 <=J�L�V�F=���D�E������H�j�I����'����<p�=vɯ=���=P>��<�z=��q��s��qͼ��<8!��p�)>�n�]H�UC�<�=O��=#,�<p������=	��=2�����<�U˽w��=�\=�f�=g�p�B��_/>�=H��BY�<sn>��޻;Ƚ�,<p)�N󟽚�>���n��	��=���<�v�=n�=��#=�F½e2/�J�6�]�<k3�=�"=Xmz���(>Pf���>�;�3=}1���L`���=w�E<�ϻ��y��<�6ٽ"9{�r!;J2=�p��d/��+�Ї��F%�=`��=Û=օ�<�M=𸀽��=/Ng=��<�?�==�t�쪍�%�H��~�=m�y�����8߽�i>.��=(��8,>�ؽ����IF�=dT���G!�8�ҽRB���%F<��`��X=��H=Q�-�D.V=WR3=�(q�XBl��{ܼ��<B�!>�!=�o�=�y	<�[�����ٷ�=N�ݹU�M����4<>\{��f��g�>ۗ�WMt�X;�w�� =bk
>,,=�;�=h�ƽ5���[�Ǜ�����%3�=<,<<���:�ȼ&�ļ�z =曝��!;�F�qc��!/1>��=݄`=��>�`v���n<�\:��=b	�<���=��#=^<z^�=�#�ܼ,<�Zw��k���5�=�y�=x���~=�fm���:|��<���4��!"���e�=z4��=����=�
=�&<�H>��=��k�'��;�ӷ�B���m�<m2��9L=;��=fU��Y>��Z=V��<r�=���~u�=�sP<��=h��;@�<�幹=6�=�iN��!����<R�½��ؽH��<�
�<��k�\��X�<���=�>n���E�=�л��]=��̽�eU=�T>5�#=��=)VE��P�c��=!^'�>-����=}}!���6= r.=���<S��ٌd�,s�0��~r�����<S��=��.=�|��*ؽZ��YЋ=Z� ��->�e��=a>��=C����>�a�=�R�<!�����=�Yܽ�I=E\�;0�{=�:= }�=���=w�8�}��=��=��S=�z�a��8��=h��=�����=�N><��&�8�>t���A���XF�<N���*u>er޽͖:��S�d��<��<�;=k;��i���#K=�V =��޽�Lb<�g��D�=v@�<7ʋ=�D�=��=0�=R����PV(��%w=�R˼L�i=��ǽ�ż��=�V�C�Z�������<�����ѽ��ʽ����D>�8<d�=ֵ�=/4�j�>.�=��^=aS�=o~�=�{@=���=�,����%�����1%:���<nB̼��=�[p=H�,>�x�=��ںK7��ʏ<e�	�/t>xݣ�1�2�O���u����ѽQ����sZ��=	=��:��h�S�ܽ��5<�н��y=H�����<c�=����I�E ̽��P���l����=�WB�5��Y�ż�p��ɻ��y����-=�a��D�i�3/8=88��H��=�۽���<�C>�C.=�>��-=�����C�e�<Q�p�$/<�,=���	SD=�J8��9�l>�����=3��<�=]?E����V��;����Q9>s%�����'=�J��a�5�=�	k���y�N����\t=,�:�R���zt�T�C= a=�!��.�<^�*<�q�=�����@6;���="�>�[먼yr�<�:p�L4�H�������.�b�<[�����H=I٦={��<u[8�S6�M�V���f����;Ə<=-MF=�^�=�H%<�7V�o��~�=:j˼�\ټj��s;�ŧ;$N�=���DP^��>��0=p)�$��=�{ϼ �=���[�=��9�T�DI�=�>�<>m�Yկ���뽏�C��=��f=J	�|#��Y�Ž����<>p��<�����{=5�C�׌[�j u<�Q�ܣ1�m)C���=+�ϼ� <��~<��
�55�I(�= )�Θ�->�+�<�v><Ӹf��@�=�ŕ�V����>��r�=87�=}8��]���d�=���\��=8��=Hv�� �ɼ��Ҽ�u=�O�B�>l���k�t��R���!�p�'�1��<�y>�0��iPq�{�:�
4<��׼�{g��g�=x��=�?=)�<�V�=-�<���;�Ci<��j��嫼��m���c�=�.�<�Z�/y����+=c�=.�=��n�:g�8�O8�=��>�+*>�x�=��a=S�޼�+�d��;v�<�ı�"W��N����a���>=�����@����}=��(��N��<O\3>��)�vW<�zӽ�I�<�f�<�^N�!1�=�"㽜����)؛=�`v<f�=��;�����qY��>/:�*�o����5��F=�CX���=F��=ݜ�����=>Bu��{���>=�dK��`��U�+�(�>��1��O=_�_>��=n��ư��}���v>�T$<�g���5�qj:���d>��>���=2��=ɦ�=���=>p�=#=e�=)��<-1e=��s��=1�E<�=�<���tޟ�m#��>o���I�<!�|<ʬ=0��<��O��o��3��B�_�h��=T�?�Y�;�Lӽ,{�=��t�y� =z
o��+���6_�Y����z���p�X=ِe=0�=��"=��>EtG���=����)���#�<�$��~���}-H=6�<��j=��B<EQ�<f�-;T�b<&�w���u=RM�=�/+�r	�=���<�W���Ӭ=����=rü��ռ�/�<ć�[-X=��I�f���M����m=l�j=h ��ˀE�3�L=�t/��B�[q=.�;��.|=w��= +)<�х=�p#=�k~=	�Ms�<h��$�ͼx[�=q:�;��n=�޼�`m��W�=䥣���0���1V7�ٮݼ���=���<w C=���
PB��Z���u�����,$�=����C�{|>c��=�q=C��=-���]=��v������o��xk��T=!�;��T>�=)y�=�m�=�U�r��{:n=C;;u�<<�W��n�����=1�<�D�=��^=F��
I�<�m�-�����������=�a�=���=��<��=<ݶ�+�=$⌽��W��� =󬦽�;�'��=;�=��e=WX�����=w���V�=&��<�[ս�`�<k�����=���&ܽ9�q�+ ɼ2S3�]"<���=�9�?Խ����c�����i��QK=?�:U^��`:�=O�=GI����&=�����=�pbI�h�����;=����l��J]=�9+��BA>$���L7=� =��J=H�q>����l��<M��~���Ӹ=�gj<���rZ��\S��==���9rl���ʽ����=�@>US��o�<<��i��;e�H��T�����<�SL�ġ�<�����-g<@�:=��3��v'>|Pn�ŋ�6�F����}�p=|ȼ�գ��H3>|)8>��0��?Z��k�?L7=�=}��< >=� T=��� K<�=s��{
4�Ȱ��D^>>�+=������.)L;k����=�P콜P=�c�<�O�#�O���P%=�����9R=�p�=�����f�����ɻ��nݽn"K=���;�� =1���ڏ��� >^��ߺ���.�=�_~���<��=��Z�b��=�!�;��������ʽ�%	<��>�N�z�#�&J�=3�*=�ͻ�:��?�d䚽Wy��H˨=�fl=I-���<���X�<dQ<�m��? =�D�;Q��=g+���=Z���<�=�k"�e�<"���P�<�LN=]41�ʹ�=��C�Q��</v[��V�=�x�� �	=�D��,_K����o}�<ו��/���I$���=�+j�AI���=��C<��ܼ>���sb��1��%>�3B��%�����ד=O�"��n�=�y�=��>�ޥ���=,���$=7�ʻ�r�<�]��٠��=��ػ��ֽ]���}>�kͼvOռ^�=l�<�E�7ί=wX�N�.�'8<�D0�	zf9�Z��+}T={��<�%=�l�7�S=�=c�=c	��꽿�>��$>�.���ʽ���<�#>}zD�\a=U�}W3�-&]�m>��{;�" =B?����>�`����{<��=�6�=���=P׵�'<=dT<�?!=FU���P��O��F�:a�E�T<�9���:�������<轸��y�`a�=� ���=�!�=��1���.�[�ѽ��<t=K���'�=�Ͻ���=<��+��"�=W%��n�=u�y���=0�=X0�������wc��ռ�'�=bw>K����<0�j�X(����=$�w;��J=&��u�<�W������༼!�=�0�=���=�u>/�=�<���=9��:�G����=#~K<�v>=�gj=��N�6�Y;�*��ˉ�/�}��Z�=�>���<��=���=��=t�Z>@�F��<�D�=�fC�֞���y='��d>�>f-����=��=��=��>��d�-Ȃ<�#	=
������=�h�y=�X~|=���=+�>������>�;輽W���ꭽ��ω;���=�{���<�� >d��1�37Z<U��������<I�<�J����;N.�46=_�~�.�:>~4��y���L��Wb=�®:�������(Y=��=5	>:�3�X�����KB>�ӎ���G<쩅=1�=��
��k�������͓�uIc<�=��h>
�=�8�=SH���k��!��&��z���/+:�2$=ZyW=p꛽N˽��=���=�"<G�n=�i�=S��<�=�;���<���x=���KP�<�+#�\j�=݉��e_�b����䎽�3��=�!����ϼ��=���h�s=�=Pq=�e�����D�<�z��2U��f���Z�<�i=Z�>�7��=v�d=��9>�r}��V>l9�<�ֽ��o�=�˼[��:�u=�׃=��ս)&M��I��f5��@�}�E<�*���G�<�6�=ݐ=P�o�:H�=�F���X�=�m�=�3�<v�$�C<k���0�����-1�=�&>N(�<`7K<?�=z��i6= ��'�:`�$>�ঽf#�=?t�=r;g>&��<�;M�=	��^��=�ͽ����|>���s=��]�}���/p=Ql���y���ӽ�,=���=N�%���=ɷ�=TM��켞���t������;{�o��R�=I"�=rH�H���<�h�:e>�=#̹=�� ��v��_� >��<P@)��'ؽ@�=�`3�q�<�H!���-��=j�Ž��;>EN����<y��=���=���>�S�=�v/=df=���Qm�=��P=b73=ƕ�=?F�=�#�����=����C�h<�,|�UVA���&>�(���^=�,>�j��v�?�lq���Q����=bqH��F�<�l�=]�K=A�k��΅=d#�����= �Z�	��=Gf�=�=L����=��ɽ��=Z�N>^�P=e�x��9Y���=��ͽ�|=����x��=TJ=
i=9�ڽ�)�;�D���S�?UX=d���`�9���<�_���E�<?J=E�!=X�=h,��ˉ����/<U�4�"r��j����&��2�"<Vc�����=*�	=b��=g:[�gq��Ϡa�#^�=$�>Ӝ���MB=��=Bǟ��9(; 2"<�N�=H��=\ů=��=��Ē��i�~�0cR=R�u�k�����:���<�&t���<��H=L���6a���=�q�=����z_����<x+�������)�=�ѣ�S�f�t���<����嗽#c�<���;���?�$� ��=�o�<������.%X<u�3=�G>�*��K�=ʐ�����1=�ŧ;n�=�3�=v���Eoý������3�}�F�-�������<��=S|��(X>8��^T�J
U�E��=��=[�=p��5�,�0��=�U�=�@>0N�=a�ŻG~p�k����/^>!��q�G�d�i��t=�U����=����3�� Ԡ�lk��b���ۄ<�՟�/s⼵�y�"~�=�?�<>l�=q{;4$��ʽ]��=�<[u��g=�-=��  �<9��=��B��.��ȁ��xk�"sԼ��f<0���ϸ�;�w��QR�<T�j=0�=E#�= 3>�`=� 
���
e�=� ���~�=Z�=��ԽyP<���<X��=e��<��^�)u�=�U�=�G˼6���J<���_}���M�X�=�
Ľ�1��]����<���6�:<���=�eƼا��{wҼ�\=��=IW����<;�z\=2��&���H�-��CH���=��=i���ۀ�,��=��<�7��.J�I�������=1;�=��g>)�J='5_����V�b<8~>'Y>r`��f�S<2��=���=`��=��<\ü:aM=������=�XM�U�=�T�;�n�<�cн��N����;|C�=��c=HpQ=�B�=�#N�S!�N��=9=�=>y�=_�T>c�+>Ka���*����㼹靽�-�=��>�c,������=P���弊Ey;) ���A�������[�=rx���E�=�� =���=B�½�Q�=OCC��K�=�7�ߎ�;ƅ��K�=DW�=���	��!>��(�=�f��|9�=�IW;e�a=�U��h7ٽ!�}=AJ߽�gнs�U=�ơ<�M��<�$<����r���=pH =�Da���>ȆP=�߼��Ӽp�=��l���1��3�-~>��0���#>TyC=�">yN<�缘��<��;>vP�M��=ġ߼d��z����!���½������ɯ;dٽ�:>��5=�荽�'���ֻЗ�=�t���=hn�<#~�<�N�=�P=2/G� �N=,��=��=8��M�=к���\��X%���%�m�>�d�$a=�a���vk��[3=d�A��ϼ	��=C�<�0�ؚ���UU=�P�=�U"��%ӽR�ϼ�B>��==���A>]J>��Y���<����N
>s��=/�:H��k�	>t`�<W�A=���y��)�=+ѽ�*Ƚ^��	�&=��I��?�;�Ԁ�b��=30>���<�	�W�Y�3�Ľ�=[��<�ƛ=E$���d>���3�P���5<�����<!n;-��G��=�_�n��=e@�9���v<}g|:����:�#����<Aʷ=q�g��l�=��z�?�)>�x%��4��+��d =rq��5u=DG,��S�=D�=]�r=f���c��y���;{t[��w�<j<���C��A��;����R�=?��=cD=U�5����=2;=c-���%P�n���-��<t��9�� ��;�=1��޽X���ݽ�Ҋ�s �Zl�=C$8��'7>P�ռAm��6��e�=�����=�/
���ؼol%�rڽ�<'>�@*={o����=UE��q?�=K�>�(=ZZ�<t�>K�<�n���<���9pI=�%��H�6>C��<�i�c�֎#����=l�5������$��]�=<3~x���}<�ۮ;濪��>o,ӽ�6��Υ�=Ŕ�=H�3=��F=�7���8�O��9_M>�k�=���=T�5�ˣ��Đ=�MA��F罢3����R���Q>p%�������=�0.�I`���}�=<AE8f�:"��c໽|�G��و=m��� �7�c�<����%��bl�<�.��,�彿��м��R[=�������y�=�.ټ�i6�`�=SQ�*>��>]���;���[���=���;'d�<|��=�ʛ�떽7�P���8<\+�=KE9=t�T�ս	�=u�9>����=���;�i=D����=��7��G�<
�9r/w�� =�f�=�"�֦>�[+\=�w=ˁ=|rj��1�=��ܽץ�=�����<����@	���V��X[=��="X�:��=��u=�!�>#�`=.s�@��=p��=�%=ud�=K���a��P��=4G	>(|ѽt=�p�;����A��׺#ɻ�u�1���2Ø=c�T�6��<�-r=v�����5����j=��7=r]����{=��bG�=M�@>�w���b�Ҟ�=��@����Z��<�;x� X��O0=�'�<�O��K���Y5�=�]��NW=3)��FT&=�D�=4�"=��;C��� �=��N�T�>=+e=��=du�=�R�=YP����=	���B��૜=�񶺰]�="�½�>��=AU��M.����m���M>�u�=p�/>ǭ��������������<���x��v�>�,�=.��ES=���=�ǌ<�Y7�!�c����Ų�=�W�< Y�����ex�=g˄=����c��a�B=<	�:>�<�>�d�=��n;02�<�=���>>���=�\=�<B�BZa���<����=C�F��
归|���I�d�����B�� >0��=`�=if�^O=>b �G8K=v)<�{;礪�A��`I���e��5y+=�Jջ��<(m�;�����ڨ=���D��<�p�=�砼Z(�;BI�=@�*>��y=u$(>�ٱ:�^<���^��=,_>[Ʉ�R۳=�М=���=�A�{y[=~�c=	��<x�^����<!M>
h
>�ýy��=s��=����-���;�������=�~�<Z�=�	���=!������=�p�=��>�D=L��ƞ�;G=w`<����_�(��=�|<���<��N=c���2�F(D�!E=��=g�:�RLQ>]
����l=85�=�����OK��!>;�K=�!�=m��<�w�<E��=�c:�C�<Z+7=�E���L�H���[2>����~;��x>y���j��4�*���>�9�=��=���<�aZ=i��=��G�L�\=5�>H�k=��=��<�RT��22�F��=i %��+�=,�F��QH����ۼ��=X0���T��`5=^��>��=a�=?M�=]��&G����踴���<H=0��沊���80 ���<[�=�q|����e�<#�=��=�ׂ=�h��6>�u
��/=�Rѽ�,�?fF�bq >c�=IA�=-=cK��?B<uh�;k�����=ؚ&�ω=�i(x>ܳ�<Dmo<�G>>h�1��>����|K�6�>���1P�=8o��+Q�w��<��<V�ý�9[=���r��=�̝��u>:�C=�Ɇ�d����vN>k��=f<߼�=Vw�{��= /� ���nʽ���~�=,����~��� ��%*�=v �=<�a>-\��*H�"��<7nM�)���`p>�ĵ�/[>���l�-={�=��u<9`�A�>�����{��'~Ͻ�cR= 콂����7�A��=s��˕:�"�=g�.>��*�H��<`��S=��=H��=���<U�;>}7=KR����=�&��R���ٮ;Q�H~n�O}=\=�=F��Y��=(@���A����:�L;��<��wn���^�=�r;ƅ=�O�����97��f�<�"ؽ�i�=�o;) �=�5ҽ� =�Ҏ=��-<�H=��=����E�I+��)�=�OD={ཪ*�@_Q=z�a=8=p������;�ʵ�t9=�3�=�
��Dyͽ�E�=�,Z=n��H��@�=\�7�F@=�F<{x�="����Y��Q=qA�=�̽�I��7Sa=�f�Cd=���3C/>��=ˢ����=�.>$�<N�f=�!�=�ژ�����G�=���
尿���=�2�Eh����+>O��ӹ:��->m�˼��=�{
>>S�;�O��⚈��K����!=�=@��<��=���=��ν���<���=���<s�P��Gj���:�䩴=�<���=J�w<��=Qۥ<ٱ�=7w�<{H9��	v<q�*=.���>�!�2�&Ѽ+ѽ���v
R�W�T�F�n=��=K��<�f���𒻘=�%8:��~=i��=�4V��E�x�\��%��%�;?&q>E�3�E@��F�n=̟�<�F����!��Z>-�e=��=�@�;���xȽ���>,��+�1��>꽷�=�7(:�1>�=�m��s��=���:x~�=s���)�=7�>oeC=p�~=X��=�G��� >eQL=��ν۴S�J����ٔ<j;�<�e�=@q=[����>���=s'<���ȡ=�+=E⑽�?*�$��=��i>��>d����=�[��5�=�d��8>ys}=4+I�k>��&�Ͻ��Q=�T@:>R��sM��C>��<{�I=%d���>c3нs��=d2=~',�$r7<��Z�'�}��A>�H�=ս1�>�y�;����佽�۽s7=W	�=�<��x�==�{�"�o��>t��U����
>��>v͢=]���j<��<��=�S���伍2ֽ�'l�5����lv)��c~���=��n�Ā�=���=ȵ�<���Z[H��K>K1�=��<ybȽ9>��3b�=8���=Y�=nЇ<���=Ԡ��Z+>����׌��:`=X��Y�Ͻ�����$�K�2=��=�|=�1o=7�
<���<�>l`���C�/��;C��������!=I�*<9�:q̩��[���=�=�#������8C=2�<�f�=�~Ľu�=���<r�"��x;$� ��<ꈹ<.��=nA>%��=}]6��ܼƢ����<�Ĩ�����bI��s�'=�H(=$����<��Ľ�kq�ݮ�<�Z=�D�<;!>5�<yH�=P�F>C S���=�f�=��:W���<�SL�-��<䯱=�`��?�6���Y�jt�Ă�2�&����=����gK�<� �=+�#���ʻ��0;~����|��8Q=�M<]@�<)ޝ��R�<ɵ4=�P��Ȝ=������n<((��d��!��=�:b�C�W<�d��jP>v_~=T?p��p�:�� =�n=4ʐ����=��0�̷�5�=.�<o���P�d�9��=kl�<�@#��ƻ=�;R=��~�n��=�KK=sI�ims��/#�&k�;�e��Ǔ�B��<��=������������3�<v�P��7O�΍νS�+�C����C>��/����<�E���׼=�=��>�H蟽��
���>��=��	��W>��O=�ήi*�fI���U�d#O=7�=�`�{o�i�
<��=���N���
='�-��b:E8I�>��<� �۞<�ta=�I2�����j��O��<i�)�;����Y�ߝ��Q��D�I>Yp�<0o8�P�B���%)˺Ju_=�̑=@��=��$�"�>��Ǽ�:=V���p"�e�>��㏽�C�����´�=ʔ+�z߼'>w��q�2慽qV�=Q�8=��ټJn*>��<���<
"�<S#�=!�׽���=�:o=��-�����᯼1���Yc=a��<݅�=�� >։��2F�=Ss��엂<�n8�6��͛~�ˑսj�=���4�]����<�%><ʠ�Ś��`_>*w<���=���	�aﴽL=}�X>l�M�;TT<���f�k��򀽜|���q�q�=`L#>g^$=�@P�l�=��=�`����=v��fi=��6���>i~����=��F�����H<H��8=�d����8<Y�0=#=� ��W;C����������� ��Ǆ;�*�;��o<�)�<��d=��&�+�l=��ռi�� �=�u�=�/нi>=��=����Λ���f�=�R; �T��<o7�=��*>�!"=�zA=ܬ���B>�]�����)��
�ݼ��*�g���K����n�u��=�}�=�T0>ڗ�=�5�h�i<F����r�=+��=��ɽ����(;��^<������<W�$=�A�U&����<�̭=w�;h<��ꂽ\P);>6�1���l��D� >ڌ�<��s��\/=O=�� �7E�=.�>>q����l΋�R!=\�D<��{���<�Ix=|�C=�<�m	=t=NU��z���	=0=݉��*��=�7�<����~��<?�ܽ��M}-=ҡC�F&\�y���+ڽܟ�=J{��4<=SS=�LU=��=3�I�-����%���h�=
��=Vk��_���	>��v<;w6=~6@;>^��:c��
�=��>�u��hl=$��dG��n�=��⽿(6>�p�$r)=�mL�N���WTI>E%C=D�=����<:�N=*t=�s<=�J�l'���1>�H+�+8a=+d@<?�;��=�N�<Pb	>z�K(�=�n�=��>��>j��<�C���l=�dD�����&���Α[��8�=>�~=1����L�=]V��g�==� �=�w��A�Aө=��;��*>�ܹ����<gR�=�E>��ƽ��D��<q�2�Yܛ<v. = -��m1�<v�<SW��"_��=�'��S�ۼ��t"����齬>:�ɅJ=��G;�򁽏y8�,�;��3�2�4#� Y�=�����U��sZE�V�ܼȾV=�?�4�Y=����b��=��m�õ�����:�=��W<���.�!�6�i=���FK�������򍜽1���Φ�<��<x��<D9=�v=�����}g=�/�=��ս�Nm�"Ԥ<뇽�fF@�����j�5<�z =�z$=ڋ<=�i���<L;�q��Vf0>�\սhQa����9��=�J�<�r0��H���=�T<q�R=�:�=�
G=��)=��;�Y6�`����
>l`=�)�<�l==ȴ;��}�O��~<sQ=�]��8�<͞=��?>4�>�=Q=��u=x��=UF�<�B�7��<�!�{̻��.��̤�=<ռ<�� =�aƽ<��<�E	> �l=,�3�"�=�=���=�h1��^�=�ނ=��=��i<�2��N]
���?�xƒ=x���� <8=*�
�Js�Gث<���=vG�l��T->��=6�q��F�<�C=��=�q(��Й=����+u|���{��O�=l�O�X�ٽ}�=o��[Sl��#�=Yx�<�n��vt��{�z�d6��C약�Ɋ�;P(=�#�j��<���<吽��Oj�=����i�>�*'=�`�=9��T�½�=��̌p��L�<���l5�:�P=�ż��H=��E��M=K4��6�Ľ��@=+�`=!A��5���(�S�>^=~>l��=2~�=i�	>͉0=��˻�Ճ:�d�<bb=n�+�Gj��p"<�p��ww���J=�0e=�k5��ڏ<���P���`��];P�</>�=��뽮>���O�BW���6S�6J>�U���ҽ,!Y�\b�:�V<#���D�<����H��=���<߶����>���;�}i��#�|��2>��ֽv���F>&|�=�̏���3�rc->��׽��� �$=��T�"�=_�ʽ�R�=�=�܈������0�����Ӛ
�L}=͜=_(=m�)��6��>�:�=c�ؽ.8;=��6=_$��T���c�:3�=}��<�ݨ=Ԇͼ��=����/g��K�"��= J��(f��^�=�<y~��%�Q=�=�,=�������^B=�G��������}G¼�p)=Oφ=�x�=�y��\��:�E����ǽО>�p�=�-=�"�*�p=.�=(z�=�>�=��<{�=�S���α<������O��E�>丝=��$>�D�=
�#=e3�^���E�=%^8=��=I/�=DL�=}n):����=���<�ĝ����=��Z��%<t��A@���<6�u��=�	��{�*>��*��Cm9��E���=(N=���<�m�<�{����=/����Ӫ�|B�='f�=l8�=��v��=�!�<�S���v�%=��ƽN��=6�R=,鵽xU�=�(=���p=��;��<f�N=�P�=�(+=!�������4c������D���[^=�r��~2=�=+�e<�����,�;M��z�=�ؼg����Y��Um<cm�=d���X<����8=|���	m�����n���t�j�4Q]=���=/ѽ>��=���=�$�=�">I�z�eC!���xE+=�F��B�=
܃<�����=��\��U��1ǽ��A=���;x4��\)�#��=e<<�+������_<D�=O	��3.>�袽E�=� >7yнqC��N��<�o�S�H����'�Փ`��q=�3?<�%?>�⃽
��w����@�<!O=��!=���<)�$=<*>�;��9$=zp=F�!���=U|μ��)=�w�<���=�9�t��=�PH�R�= ��=G`㽘Pּwd��M�=��,>
�(����g�=��<z��y�
}<���=�=�k=�z�=�Y�;�zN�h��!>O�	���0=8��0ZS>_|�<�\�s�=�ؽr����	=;>���=�A�bb<9Z7���<���|R%��u���q�#i�<q��:պ���<��>�����:���=�T2�%�<�̛<��p=�ʻ�\:�e4����;5���$��a7y�� �<Qj򽕁Ƚ��=��>��>5��;��zH>Nzݽч�<���0=�Fɼ҃�=X��=��>kNi�I�޽J��<��n½8����<��мN��=}��=6��<�L�=�l�So;>�����@3=��j��g�q	\=V��<䓝=��=b1�=�J��i�a�������:��`�=��=`��<���=&�=q�7�a<l��_�}����;=������1��Bt�D4n�N�q=��P=�*m�R62>�)=fԟ=��%>A�K=�+x�L�;��=���=$��=���o+8=���k9���X>XՊ����=���"�������2D=��}�����k�C��S^=H�q�@��B���$س=�!�<�}=��޽�c��5�j����=�����BV���b=M%=E(=`����=��ͼ��y���;��==�}�=�)=K�=������=�K���)=�"V�ה=�`	>RV����=�`����9;^� <��Ͻ���=]�B���8,=�8Y=�*ϻ���q��=�ɼ1Z��>=��[�o,�=���<�j=�
-��F>>NQ��B��`�=��4>�
)<��<��D�9�W��VH=;��<�4(>Q��^���~�=�R��Z�滥��Yӽ W�>�G�=Jߚ���W=�7=���=�~�<A=GU�=�=^j�=��3=Y>�<�;�bҞ��;Z=_^Ƽf>5�=��=��=|�0=s^.=���/�q=��=	ne�It=	Z��v5�p=�2����h�J��<:�м^��=�����(	=�o�=p>V�s=�˽9Y>��>
��|�=V�M>U~�<��?=�GлsB��Vٽ���=�����v=#�R�h�=�ἄֽq0�����BP>��#=��T<h��q�.>Q�<�e4���=H <�$%>ǘ�=��k��/�%"e��F�=��=!�����[�U^�=i�>m��;��=��󽇪>���� $����*���@��+�<�kF=��Ƚ������μӃ�=	/�����<y�=��=�k���l������!���}�<�#I=�3T���>Iⷼ|>8�ƽ+�>$��)>2-޼��3�,n�;�B�;L�׽���=�ᢽY�=��e=}��=/��=\������=/tѻ�B��؇=�Ua���	_�O��=q�x<.sf��&�=г�=�UH���
�ϛ��`=���g��<#��=tB
:_��=�
+��oX<���=�[O�uk<��<u�{=^%ʼG{��=v����= �6��\<��=�<�W�3��+73��^>;��<�k=6 Y9��j��^e=��<�Ӥ����= <�)��=����n*��d�#>��6�ԁ뻉� ���:c�<��X+�=�d�=��e<i��=�k<�$e=�t���9	=M4��@=�N=�/=��������$����^̽����K=%��=���=��b=���<D��=�kڽ4�<׋_��>�ʿ�������<��z��Q<EĽ�k�=��.'����:��V�O���=���Z��4yy�#�>V |<�E�=��ǹ���=Oy���L�✢�ps��
e�<o���W�=�vü��1��=���D.�<MP>�P�=��="z'�<^%=��=�E���A=��6<<��Qמ=$0��B��Ŀ=�>6\���\��)�<>���-��1�>v�=�I�*��=)��4F@�B>VqR<e>B: ��B�=Gތ�)�Z�Σ�<^��=z�Ǽ��erܽ�t���U��=!�=3�>}�=��i�'���⍽�5Ž�d =k�D�,��6p�=XȌ>�����=��<^1>X����P=�~}�Χ�J�,�c�e=�Zs<>�k�<�=b��<$BQ�M��y������<�ѕ�W�������%<����=ɖ)=1�ؽ�B��zlC��].<nt>EC>��o=���=�m��.�<��>�������=��#ü�fZ;b2<ge�=̿ѽ�|@�Gs�=o�U<���<��= <a�7��a<�-�������=C�(=iP�����s�����]�9�4��	��5�;��l�Nm��7�=�����E>�i���~���=�=�͓<���<��>>Y���<��>�F=�M��bw��U=��ü�ࢽܥ<řT������Dx>��X`=Wȟ���-<:6P;�-��������C<�{I=4x�<q�������6>�5:ũ�=$�=!��
�=�L�\�S�T�o=�&���̼=aC=]�<�V=�դ=r��j�k<��=ʞ��G�=jӠ=��=h��<%Q�=S��<`橽j �˦;-�=`|>�Hk=��G=�^@���<�(�=��=�.g=(7<+h1�/{��BK=�y���s�冡��<��ʼNDO=�7=7s�=,�<|0<[�=I��:6����˧<�~V���ҽ�lp��
!��0�D�<ϲe=a�E��X�*�=N��۽,g>v�;w�=��+��Rd�cu��М�P�G��	���Y�<�
=�>�����總��y1ѽ.iO=�@;�~��{� ��	S�<#R�?6��U��=u����T�8�l=���<I��=�3�<�R����=�ע���d=�X���w@>�.=��C���/¼B2�=�����`V<�H��$>?��:�3<�U[�W��8��=�O$=��=��-;� ->�NM���ɽ�K >�<T=˽L%p>gO��5 ��>o="�估�I�遉=	>�:�!���<��<<9�=�:���=��经��ȡ�< �E��>Pi�=.h�=J�M=e'��Q�<E���B%���	>�k/����=��d=PE=��$����<�q���̽�t^�^�<eũ=@�j�m��AR}�@#=}uS����=��R��R�=�B�;�k��;����=�y��t�=]c���켲"]�˞%�CH_��)�<��<ٿ-�,�;B��G�:��1����<'N��f�	�����ϼc�C�\����A��h�=#M<�Zv�	��H�=M���=�s=���<�:;��=fV�<��<��=��<�u=��R���%��\��G>��<V90;���;�}Խr.�<9�0<	�=��d��N̻)sc=zR�='
�=�����9k��݄�a��=�5�=���=���=Ǽ!�ҽ��=��U7�;<)��1�Y=��-��r�=�P< H:�B�=|�,��uV=A#�<��=�C�<�eM�c��=� �$6��K{����ы��[��<I}>N��U)� s������9=&�޼ܑݼN㰼`�;��&<���b��;쎐=���=�Ϸ���q�7��W��e���W3=D=X<+XN�]& ��������;��8�=<�;�<SXH= �=�E�zd���)b>�)���x�V�<=��=a�O=�I3>��<"���,�h�;�i.=��
=y��=.R�����A�*<���=�ٖ<e��>9ý9���I���>�\��dy=��ӽ�F�:M�����=�l �y��������ӳ��w�<�,ͼ���&mO=d%���tj=Ftr�[$X={�������<=}�
��"�Hv�������h���=��C>�2���->�(��	͛<�_N��
�=�(�<)�}=�И= �<;��u�=�^=ǆ_��0K���x=)zX�\Ġ=v|���>��� �,�9R���	ڽ�2���<=R==;�5�Җ�;x ��3k�=`��<dQ<�b�<:Ǌ<`���0�<W#������?�	b��U���[��jڄ=��ռ���V����<Q~Ѽ5룽p����>hŘ=���<�9�=���=Kn�=�>��>��>���<�o�<�L�@W�=�4�;N.O=�P�9�Ö<���;���=��r �<��=\��=p "�F�>Sx��}Z��#�;�� �(!N<��U���=�C��23i<��'>��x���
>��-��.���9�W�4��
��IU=�R�=_.�<*	�<�<�=��==������%����=�����]=S�I�&n�)�=�9<��G?<�	�:��=�.2=��N���0�h���u<߼�S�;V�b�������C�ʯ�<C!�Q��;�-><�­<���9���Se;ts�=L��9��=oL"�^�<���@�Q��]C;�=�Sp=iݛ�]HK�|��=�D�����Į�<�T<7��3>#��Y���O<��=�o�=j��=��8��E�	�b��0=��;�+W=S������=��ۻo���I܁�z]��t�,=���<:?	�6�+�x˽��'�6I�����;�(��v�;iE�=��p�+�ټegԽS�>��>��Z���м���=�`>8ļ�Q=p�}=�,�>��k27�*a�<�7L=��Q[=>d�0=o|I=��B�Q>���=�TX��]�ˀN=�����$��'��=�c�������<_#X=��/>$s0=��<���=��潮�>�v)�0����hL�p�= ���ǽ��D=��$�	{=��?����g=�=>f��=�D�;~�K=��<(25>���<r>r���U=����d�=��v�y=Zd>����ܞt�M皼��
>���m;=ƫ=�T<��<_7��4ᕽ<l�=��n���z��D=1�ؽ���c�/=�z��ҋ�<4��<s�w���b��[> q��Û���mA�����-����=h��&I=Mi��Ed��*>���<1�T�ڬ>"��=y���g�<�$��w	���=���M�Gc��O4<@����ǽ�ޣ��kս������;�6/�D'�<�� =6�J�G��=���=1�=�g�;�.�<�.>�Tl��_��pZ=KP=�֜=�X���v�:vP=͔�<9:��F�F�z;�%��VF�<15ͽ��<��#=;^���0�U�>��=��->s�o=���8J���:���FJ=���:E�=��=�x
>�d�Ō8>��<��@>�� ួ�-a����<_@j�Ͻ��x���;ͣ=��T=�=��d���
��RT=���<��k�>0w�����{=�mm=�3&����<� ȽB��='G���*O=�>���A�.)ƽS��H�3o����$�v��<lH=u������� t�<;I>`¥��,>�S�=k�������=�r�ݮ���$>v|R��ے��'=�2�X�w���=]��<��ؽ��{=�y��q�<�e��b'=�������= �ѽ�1����$��X<�]]<U�= ˾���.=૶���<N�3>x�N�l�;��=`�����=�K�=�g(���=)����=(r��1���+��{���X��=#>��~&��q�;��x=f�2��?=0o��;��#��=L��=Z�=���~��ݼ�=��-���=A�=��DϽZ�����Z>Ƽ�Lc>���=���=�:e<2��:��Kt.�/�=�C-=��=3�>$I���	�P���F>(�����j=��޽�X�=sI<WB�<,@�����3&1=�(�=ǠZ=aav���=_]�&>V�"�L�8�|�;<D��<\��=��$�:�=�����ɽ�K>K�p�����IĽ	8��@8ýv��=4����40=��)=�\�����<�6�?R��� C=��ӽS�n�.y�[/��%���>I�=��A�����ꐝ�1�񽯘�=B�Ω=��L=;v��H��6+/=��=�'�;/��R=�բ=��>0�� .� �F=b7�<Uv�[������=���<G45<~�=9EF=e���xV�=���=�_�=�(�=�B�ڠ�=ˏ=���<�|�=]=B䐽\�żv��lE�=F=��r���<�����<qa=�=�'	�=í;4��<���=Y�fE����*<|@_=ԇ'>_<ڼ�Ǽ�	8���+�Q�<kb�;��7�l�>�v�<���<gV�=�Y=c"�=�,�$=�]ϺZ==>�}����=G>7{E�כ��ւ��W�ܽ�ֻE�=<�%>���3�4���<	��<l�=��=�n;��ޝ���Y=�	G��=�xm=&L%=��ټ*�t���Y��1X</��� eA����<ʊ�=�K��3sY��V�9�M=7�պ51�=ԅ�=,%�<�9��6>)<��>(����S�= L�;vR?=9�I=�17=���=�Qx��,t=��=��/��=CKڽ��>���=��h���N/a=��;	�=X����v�=R�,s�;��='��MV,�.����Ľ{�'����=��$��W�7~E=#�=�����:����t/�<��>�V.<�����)=���Ū(="�=
��=�e����i��=``:>V��=�&����;I�&��=-C�;F!:>3�y��<C;=�6>Fd*�MT+�F�ｏ���6��=�W=F�=c��=H��(L#��:�=;x=�Ȅ��m=�g�����K��@�h���=�p�=�2����P��=Z����7�<㑼��=Ř�=��o;"�=�ͼ�;���	>�ĳ=�QL>0���)�����=�L�=�е�4v����=����<�:7�=~�Ƚ
��=O	�;��F���Q�Bh�=y��=�6�M�<�t�=�5<8(���K�/��<�����8��NU<�P�<���="�=�Rh�iW;>����{>M>�U��%�=��=�5�=�=���=�#z>�_>�2���<�U=>��E�=��<|&K������j�B�#�{��Y�/f>8|I=I�	=�0��9��<���;��=�+ֽߤϽ�Yٽ�f�=��ż%�6����<����R��z�C=}U�=ŝ#��U�̖�=�;��
�N,>�F�=���q>S����6>��K>��=	��<�x`=�M�Za�=?񛽫G�ɢ��S���[�N�=�N1=�_���6��L=�o�<*`'��3�=�,�<�D3��12=�;�=N��<�<�g�S	�<����V�r)n�"���������<�d�=�Z��'��
͇=�d8�l/�=\����=L+�g�p<7�����=6�z�o���>���ZԼ bg�5K��	2�Lc�����(^��]����ۈ�=h=xp&���o=r�)>�+=*z'����<��q���V�=¡>w�;x�v=�x=�� �r^;�Z���n	��bԼ�8<�����F��e�>���<��ļ���.�q=��Y=���^�<�s=@M�;��n=��=�l��/V�q >��<Z,;j���fGŽxB=ɛ�='��=�����z=��,;�S��n���4��{>�%V��	�������_~E�]��sL��{2����=����N��`�-=2?���
�<���)�=y`�=�e=�7�"��<��b�g,ֽT��=F=%<�^�=��м��Ǽ
���S�`�B>_=bA���l=��4>�n���ƪ=�b�=�4���f0=XX�=�����=�F��=�t������a��&<���=����W���V��8�=K/>"�= ��[�TF��7��U�=嗽=�w%�y�|��}�<~Y�Ľ�k� ��=G����=|��=�<,�=!�S�����==3���?�ռ�X=!b=��-=�˫=+�=��<��<J�e>h ��u�=hP>���< �=�7>�7���]V�`�x>E��<���Z�k�w��=�R�=_��A�i)�n���m��E=��;�1><��J�F=�U�=�$<#+���!W<[��=p~�<��=#��\��E�=�y��@�1��颽T��=����:r=|�=S�<�����=�|�<��Ƚ�*=9_ȽQ;��B�=�v�4�t=p5G<�-R<�aA=�;����=g_t=�3���K:��(��&N;&۽M����8�=oz�=݌����=�[ ��9��2��h����`	>͋���Q=>�=(a��rF�>S=5M�=i�I<b�=i���7��M?<S؅=UD�=�J(�b�ܽ�5�<+a<غt<�+��۶͹�İ�U =�5Y=�<%��#=��j<�H�={'=��$=(0�<y=C@�=�r'���<���י�=�݀�9�=F��&/��"�<�Tm=��R=�Ơ�Y�>�z_�EO�<�f+�z�<;�E7�
�����'=�B��X(��@%>9�i����#㽠�=���=���: u>�ɼNs��_>>%�=�$�l�n=�W����=�ت�w�O��©���8=�P�-MC���;g��=��I=�]�<�� �k	�=��;�B�:��<}Hk;1�����@<%W2�y�=1 ���0q=��G���{��<��o<hg4=���=�@�=�"��i��=��P`��Op=6��ݿ:=%�=�=;�%=�~��GA
�;��B��<7�>u���ޓI<Aj=�rB��8;;�%=ь�(K>^�<�;�=��N=Tv�0���P��ȕ<����B
�<B�=�$ϻ�XU��SY=/��������;��N>_� �`�C��,�
��=�{�e�HƢ=+e\=T�<>,�����<�Y=D�2��E�=�|=��t֕���_�P'�<]��P>>*/t=P#r���5_��,ϻ��.=���<��:�x�<Uj�=���<�>á���lR�+>g����.=���
5�Qڢ=����P�<�nֽU8��+>Ҵ�=���U��:�bٽ�9�=��3>��=cJ����9;>�(��s��}-��]2=�5�=��F��70=�$=r*c==W5<�_��w���M�E=z냽���M�=��ѽ�=�Gt=v	���<�#i<^��zK�=�;��Y`�=6� =��<mfi<����j&������]ʽ,r��/2]��pK=�7�h��=ȅG=j5�=�SȽ/L>���T<�쉻_��=�b><M_��C��:'�ۼd��|X7=$�&�η�HDo��~)�s8>��=Rp=��X���AS�sKP=�S�=nT��5G=��M=L�<�;U�\ ��G��=�e<��Z=%<�t>[1�� ��=�ҽ�+k���>fD4�V󝼊��=�Fd=�w=.�H=CE˽CB>'��=ʊ=��=���=@Sm���;��>5Z<C�*;�=��ҽ��=�m���� ���i=I�`��Ѣ��c��p=Ɏ=ڳ�<;��=��<	���P����d=/�G>װZ���B>k�S�����$�=��=���ػ�� �Ǖ!>�K��]��o�=���<���=�������<�$���k�K�ڼ����wt=�0Y�~��;�{�=���� >�lͽNb�����<���=|�<�(g�;B�M���G��J#=Ю�;R|��0�� ��<�xԼNo4��0;=y���OZM=�-!>��=�[Žz���@�=��<m�d<[�D=�������<`/r�>B����½�q���:>��������T��5ǽ�}y���]��I[=�n�%z=�ۻ s=�:��g�'�La<�3=�>>_�=�����9`=��b��;�=��4�U:����kT�5U=�l�!��=?�=���=�b�����:%>1�ܼ8����)q�#����>XĨ�����2�F=���;�y��pH4�~<j��=��6<F����p=lGm=&ka��=+eu�����w�ͼu&�;6�o��ռB̒�Q	='e�ޫe=��b�?�����=�F=�>p�缀�=r븽Hc��'v�Bѓ��B�<ʭ>�C�=�J�={ �<则�x^=,B;>�U��i���~8��x�~=�2 ��*�����.��=��ڼ�z���D���X�|�Z<(��<U�r��>����W�uk�=������ڜ=�={��!��=�V>[5̽-ŉ��߶=��	>w�,������s<�>�B�=$w�=t��<��<�x��|�<9=<"�=��=�ƙ�N��=�Z�<�9|�Y��=+�V�sn�=?�">W�d�=�O�Yv�=�M6=!>.>p��;o6>�l�;�졽������=M��=��f=2�	���=%�½ �=��$�=F޽;gy��2=��ʽ�T�<١��IL���-��1<�*��G9>>��s�<����hѽ[��=�|�P������N�� �<}��=^�9��Y =A>>�z���^<B6>J�����?�N��0l:�;�P"7��ym�R���ڽ�;4=՞����<X�$���w�=b���N���'�w����<6f�=z J����׭w���>>Ke=�V�=�=�H��L)=���K0��n������e	�=e�<v�8<��g�VM�
�Q=�u=X��=o	�=Ѭ��?=�I����<a}�=@i;�(�>����b�>�%���>u�F=�;`ǽ=Y%������+=��d=�A�=��<�i����=Si�<t�=��e�ۼ5��=��<�Uo;`�={��=�ޠ=��1�_�g=��=���=5>(�;�^���=���=!�<)�t�u���:�U�gGμ�]�<�Rp�l6���z=�'�=�J=�헺�h<`�l��i�<�y��#>C������/>�*�����=Lu��II=�ѡ�j��=�P���K�=�g=
F�<o������;��<����=�o�:����o�<6�> w�*?N=��[<J�Q��;�= Cڽu����>o=B^>N.f=K��=ݖ$�I�1>K7=��==lz >B��;���<��d<��a=���)�;㥬=w��G��[��H�=��F>�<"���#g=Oq��&z(>΄�;� �=j��=Qs\��ل�W8�<Ox�=/�=�ۃ=I1�=�����
�=�Cp�i�=I�>l��=�L/<u�{=�νײ�=0�=�p����<=X��1�F�W$�=��=aب<}��<w�(=�'e��Ė9gŎ���;�m�����=ʡ���Ο={�=[�0��y=�]�=��i<��=��ý��6���t���7�_;ѽ��:)�=�T����;�xj=�M������<���<�𮺯kO���=��b�7��<���:��X=ߔ��NE̽�%y��-�=~׼��O���={C8�gw+= 2�=��j=uܽ6bj�p%=���.?.�W�=��T��⽎	�<Uh$=� B��X)��!�gn=�%2=�`�����M�>%.��|��=:&K�N�������o�=k���}H@=�i=$�=.�>��T�s<��r=-�7=ֲ����ѯ5�̿½�z�=�u�<�H�z��={�}=y�F=���:<Q���Sc+>�z����;	~L;c�*��l����<�t�<<{��=<v�=�¼�f߼':�=�_�=C�H�%�L>���ee �-�U�Y���;�ӽB,�+�w<����o��<l��<̹O���=�K���y�t�<����<�O�=_�=>&�V<�+==�)>���=�r�=�xB<t�=C��=o�=�b���8�Z�<EV/��n�=}(C=� g<[� >�l��;���h;��f�I�N<��=��K���<{T=�Ku�9����e��D;⏰=�<U��=G���f����5�C��'o=�,�=`�'=k� <,(�=H�=���<�ׁ�[�h=�c�=��=M�;� ;�����xɻF?=#~y<� >�����;�z,>��=�w�;���������T�{Ð=i��=4���=����8=��*>ˡ�>��W=��-�@l��N�= ��=^�>{��<�W�/D�=��<b
���[�ޠ�A�k={ >����Ǧ=��� Ԥ�s�f=Qhἣ��<�Y�=��A<��!�6&Z=b=g#t�D��=��"�:�7�=m��=��>�&>��>�=��^���3�FD��[��= �_��<�y<��>)�F>���=�oB���>����=��>���<���=;�=����dN;�ۧ��5=ܓ�=�}�=i�=�M��7�=G�=�<N�C�9O>��<���=�N�X�=	#[<k��<v��;gj�izg=f�=u����Q-=�K�=`�=�g����<ߕ�&{E=�5=�a<5<��e�%�Ž���S���"�:�=]�ϽT��<��=��<�����=�8ڼm'��T�;دz��P���|m��D>�5�m=+�����k�@�٣��"��>�fn��=?0����%=
m����=�>ٽ�����>�f����=2I�=��<ͨ�=�@�<<:���ˮ������=�<��=oN�h�=^��=�B��Qr'�5�!>�dE�H��=�����=QA>��;֩ =$���ß<>>���`��={�&�>:l�n踻SI�;���=|�F�K�,>�|I=c�<L��=�2�=�0���k��ss�t�>S>������<N%O=���<�Zҽ�:��Y>Dȼ�|��%#�\4���l<$����=;>�.<>ʾ�=�j:A�0� ���ct�< W�����=#|	�ݼ�=$�=�ļe5�=��<�֩;�躼C���I<В�5��<"Ĕ���A�uԪ=,%�=�8=�`�=
^�bP̽K�u��=րؼ2��<���23�~ď=�C�=o��=ڬ���[=�F�=��+=���Et�v����Wv<��=����(<u�<��$=�~>�߃�~'�=���
���;	�:4��H7���� ����=&@=���0m=�t^�W=��=�*�=����,M�C"�=I�=_�Z=�d<h�	>Lܡ�cV�P�G=�F��F�=g8�f�z�?NC>q�����I(=2���W������<x�輩���[.=f��W�ڻ��>�
5��4�"�=�˰<I�ӽ#���8$�b>��I�<�(m��ݴ=P~���&>��C�����O��"
��r�><Q6�q?�Ֆ�=�9�=w��<�Х���Žë<��=�刼��ݽ�������ؔ<Z�[=0�<����<��=(t���=��<�=�z�;4��<���;LmW=�D�;���rIX<�{l�B�X=1�м2@���=R�=�v���;>)��<Q����>��=#���I�E�>e|��ʼ#ӏ<SBT=�P�=x;�^��C�>$$�Q�=��>�cb��C伢o�=�)>�:!M�X�a�z�>m���xż@�>��L����<���;�>r��N��<p=p�� �N�<�=N�u_F=��(<H�	��g����8�K����
E�u|>W��EN
;|����=~<ǘ�=S��<n4P��O<}�<r��<�,
�]~��4_�oY;썽̳=�+F_<R�}=!C�=,뾽a[=�?�c�-vͽ�[���h;c�B=1G�;gν��U�=�x=?�弁���0����zd>s�ڽ��$���ܼYq�=��8��D>��cT1=�o=�� ��1�=��V1<S�=v���ɖ�=�)߽��<&��=4�w��ғ=�d�T�%�~�=�x�=s�=T�Q�<3�=���;}j>�l#��&(�	U�>�	�J��BM=�O�;�?=��4�!�=Y6s<��=�Ͻ�(>Y޽�W����Y=yly=��=Q̽-JT=D=-L���{�}��=>Ȧf=[G�=�D<# �=;}���5c�� ��a�	�"�G=o�';
>ݽ�Ԣ=��;=x��=�w�=�EH���=��<d�=%؃=/l�������^���<��=g>rEE�y�>�B>�*E�ο:��ֽ�P��P6g��끽�<��R�;���=Ĵ'<5D=����:��>p�G=��Q� �=w�%���=qT�<=�l�$?z�(ڵ���}=H~�W�E<rx�,�h��!�=������=�K��ht[�����G������=4B>��=��!=��&�Y�W�f|I=�=>F��4�8=�iͽo=���:P%d�u�н�-����7=}��=�#X��3!���@=x>����7�Ä
��Z���=��M=��=}�,<.M���,(=���=�3�,)=�\	���=X"�=\z�!N�=a=���=��&>ip�=��m=e<�%	�*�１��=�ס=/2>T���Dc�~9<+�ü�6��^.��)��-9�gO=><�!{���$:�(�e�:ǻS��D���<��0̼��>�i��<��">����A=�Ό����.�=�;ƽ��<��%�<�,�=Nܻ��\=�>uN
=��*�"�->f�/��Q��0Y=���<� g�4����=VQ�<������S����<.�b��<IZ�İ��F������&`>��������+Wؽ͖�=-�x��=��< <�=���=1�L�==�M/=޾X>��J�6�c�'({=U>�=�g����ĽS�\=�cv���'	>��i=&��=��W�N�Ѽs.=Z�;в��3̼m���R�}�v�ӽ���<�Lv�����J8�Mb��@���p=���͂�=G)q=�����!7�O�9���>���=�᝽m;<H��UD���!=�t�m�:=����Ң>E��<��a=j��=�L�=i�;�E�
�>�F>	Y�����Р��i�J<9��@-����=�������#=$��i�%<��@�=���- <���=��ɽ�ݑ<��>��(=��=��>�tL���>���=�E/���5==�.���<�\">�J��0\�Nώ=���<};���+�=�:B����=�r=}��<����!�ɥ�=p�f>��=���;�ɽw��<����b�%��<rh�G�e=n�=�t��]Ƽ�@e�Kӽ{��=��|=��i�=�/O���B��~̼$������BU�_Ž�y���!Ƚ:*��=�lU�������<�Ǽ���J�7<p�=��<������#��}�;1�<V�<�p���P���=��[<�c��LSO=�DT���<iz��Zӳ=�H�<�Ͻ��A:�r=3H5�;���������<=
1<��=s��<���b�@=6'��П�<lZ-=�n�=����)=u���L/=���Y�պ�e��>;���Tf<��>��ub�� ����j���"��v&=,R=+D׼6D�������=��k��pǼ�z��v>B��=%��B=�P���Q��<�3���Ae=G
�>Z$>eQ�=yOǼ�k�=�Y�XJ����7>�^� 8��|<=�#��2�<&�8��=�	���w>v�l=��@�(��<�����=^/3����=/ɽ+��{�,��3��N�=Y�>�p�<פ�;U���:��U�2��Q<�}><�BӼ怴�D�3=�R&��\�|\��4�5�����=5���f�4�n�v
"�	V�.ɗ��{w=4H�������,=z�g�P覽�I�=\���~ĥ=8�ɼ��={jv��a�=���0��F�>}���!�">ࡊ�����轼O� �ʴ�=���=.×<���=��]��bS�˶׽�4�U*�GӐ<�� �8�<{Oʺ 6�xH&��	�=Q�qZk�������<|��=o� ����=�U=jb��a�<%J>��+=���u=>�7&��4���ӻ�콜���(>�/=1	��q�:4�ƽ�8=_��=ٶ ��J�=U8�=�䅽G�ʼ@34>���<��;�9�<5���MdƼ%�_=��D=4���)���<���:���<AN�=�p�=ݥ�=��>;����d�;� �<�1�� =!;�팉�V�W<r��=����h=�5� ��=�9��e��Kٽ�P;:Ym������Eԫ=�><��z=�iu=�]f�OC��?��E<;�G>�Ĉ=3��Dy���1����=$w�u�j<rˡ=?J7�䵒=<�A�=C��;���o=�<�'U�"w�Vv��I/�د���>a�Y���K�2���2�=r�=�M�=K��=�۽J����s���m�<�J;�p�;�����:���(=�=9��<��������5�=����<�B��:nL���:�^�="�<q�E�s�>��a=�(/<������K�	R�芴=�o���M<�!ν�w��1���伜��<�q�=+1 �$#�=<;1T�=���������=�=G(��pS���6=z(���=2��=�&&=��=��M�U��=���.	��+1;�'�faE=N�<�PY;qw��[1�;$�};��=�cf>�&=�.Խ-a��E�C�&k����<_���$�=�pb=4�/=�2=�=�M �d��=�2���	�]�2��^&�a�Ͻ2�=��Z������#�h,>�м�����u�=+�ֽ��=���=�}�=�=�|a�Zٌ�3��=L<F�����߮;�{%<��m��xY<��=ȋ�<c�,�6��=O���@�\<��|��%>/^ܽ�b���s�q�=��ֺ$qz=��,����5>�i0>J+�:id�=ֶŽjGƼF��E%�sF��kF=�֏=�䤽f^<��/=�a�!�*>�U<J�=�h�<����}?��e���'����=B
��3-�=Uj̽z![�z�R<Z�>r=#��;z�潳">��=D��=�}=v��=�x�=�h�c	&��H>����9�C�5`�<�6=&3
�A��=]�=�>�]=��=B�>ߊ�=P�	<n��Fμg�>��<ϐR<�+=��8�R.���2/=����i��Yܱ�pH��r���;��.����l��� �	�=��;p�T����=Jƹ<�!�=*��=�5X�2Yw��5R�%��D[�="}����8=䈨�K�=+��U�<Γ�r�����<,5�=������|�4V�<;�=}�=.�=�t=���=@�¼��:�2����=	�{<��#=��Խ�=��;��=�3>�*=`�����=�#Q<�:ʽ�gý�`�= �1������=p���P����<�w=я�==eT<�E=�T��X��=��"�]��=o�=���H�I=�!=
ĩ��^���>�#O�4��;�����Z=���=b��x8>��@�V�Z�e�>2"-=�S۽&���/�=�����P��=�9O��A�=���<Ӣ��h��;�	���Ѽ�).;˃�t��=$�߀��o��`S�����v�<���9`i��+;��=���N�(=���=k�=��_=�t���`<=M�<��=�콙{Ҽ5N�=��ٽ�	7=���j}ʼ��=8sZ���7�y��<����<�=�Uw=x�'=��.=�=�^3��&`<:b���F�z����R>�̔<�i�RS�=�<� �=�9��[ \="����=�&мx#�=+�｠�>͢^�H��mZR=q_=�i�� �s�W(¼1磽
z���0�ݱ����>=ҫ���j��߻D��M�>>'�h�����"<dy�����=�n���Yb<�)׽.���i�A�5���s=L"���T|���=�Ά��{��-}�=Ta�=��ͽ�����P=�mJ=gQ��T��V�2�j2U�=�->^���ך	�zT�<��<�S[������=�9?�����=u��OM�=�r�<w]�=
=~��=~O����W܋=�B=�x�=;:P<�H(���<V��=�r���%>�����!�J��<E�ؽ��=�-�=�O�wGP�� >)>�7��C弮x[�M� �#rK�n}S�#�>�$=�;ǐ>��<7{��4��=�`��
>n0>��K���>D7> es=+�����=���=�佚��;n��PM=Hge=�5�=��8='���*:K�=K:����'<�1�.5�=�A���S���=$�`=f�ɽX�>�kǽC��= �����I���=��ռ�K �0Ӽ� �(ֶ�Ol�=��z=�D�=
Q>�����<v6��CE�=6���&���LZ=����
���$���	��8[�qw�����ә������#=��<v�|���:<������=��;<�]<$ �2ɓ=I�5=g���(;9,>��=U9�<hp>�ļ,���7l�Y���z<k'X<ӵC= � �=��<+�N=����4
=�Zɽ���9B�=�֣=�_(��<���6�.����<���<�=� >2e�<8�|=�m�߿]��;?<A�S��V��D\f=-	="�<�V�=�r�>a��Y����<��=�����ZŽX����q=t�&=B'����%��
�=Ա���J�<ೋ<�����B=Tw���>{t��5̜��,M=������ּІ=�{�������駽4I	��#\�a�5�uS=y��Öܽ�E�<y��:��=���=��r�LὝ�R��_=&�;��=n
�ބ��Ø;�ΛL=��=��=!���Ô�=q��Q�>�A��?����S=Q�F��=���c^�c�Ȼ���,�<���m�<W��]K��>Mg���m��s��=�=>z��= ʵ��)*�ښ�;�6 �D�Խ�^���h=p����C��t���\���W6:ߣ=�^�=��/�>i�o<C�B��Mw�1���~ʁ<������Am��m�=��?>'��4�ʼ W�<:� !��D!�=l��=�����T|=I�0@�� k=��<�3=#&e��� �V9�Z>n�w�v���+>�?�=n�=_Į=t�y>&�`=A���9�3z�=�t��2�=2@��0�>:)>� �=��ȧv=�Q��A>�0��OMH>Ⱥ^;��� 3_=�
���>X�s=Z7���{��oC=�	=x�w�y_Y�u�=�Q��z�=�*��3��,=���=y��[7�<b�=�漹��<:�e="�9�ؿm<�=As�=8od=�;˽���xbv=��%=�袽q*�=���=j�8��.>��Ѽ�$>QL����I��<K����<0uT<���<�}�<����v��8,
�=�̴�;�>rԮ=�|�=��=0�彅6��.�v�!~q==��u
l�[�}�)j����h<�>���;�r{=��>s1�=9�=�Ш=Ҹ=�|[�[��=�G=|��<�wU=�����5��1�;9��=�?=��"=��=N��<O�Ͻ}�>2
���%��G��EP=�=02�=��o�婥=���~�D��=4e�N�
��(��4>9]S=8���c��<�ϼ&��3x彤�	>on�=V����y<9(�q�=[eʽ�=sQ�;�9�w�ȼ�,� ���v�=�sI=@��=.v%���t=c��a�P�Y�;����������JS>��ۯ�	�� »}�(�9C>`ٽ����l;�F=�A�=����y�<�b��)��=h]&=&&�=��='u��jĈ�Z�=�d+>ƶ���r�=8%���vp>��\�3p=lVa=cmH�I�Լ�7�=��r=&N�=\Ӽǳ���5>����A�9�s=뱑=|H������7�<A�*�Q��=)	�<�G|;��<��=�N?����<}O���=�_�=�̼=3c��;;���˦�=.��l;>3��=(����O=b#F����=2�=����ё=xТ=����l=O[�:o�==�f_���5=Or��D�[��ѯ=T�ؽ��h=̺O=������&���@�P�<>�>��<��ܼZ+�=�
h���>��;z�Ƽ�̽y�=X4 >ׄX�7�y=N�A�ݻ�<��"��>nK�=�6Z����>�<+���-P.��8ٽC�i=͓}<nR�=�{�<����B�=��U�# ��K`�F��=#J ��k�<g{���N��*"�=�&�<�K˽:�׼��Ž�6�=Oy�<��
��lU���o��C�<�'�A;���?ܽ��yj;�hR;K��<����~ƽ�h=��i=੃=��½��=��-����:=��?���*3b�)I�=�f�;�|L=�+�q�L>m0�-X�<T�Ļ�9мNlW<���;@����=7Խ}�K<��9W%#=x�=C(��!ٻ~!�;��A=~�=�a��j@Ӽ��G���~���;S��;a�꽭'�=�)	�D�>�� >\/=`�>-lb=e��=Mn=IT�=�3�=wڎ<��Žh/�<���=���>*��ie�=�e<��TX=�wi=z6��aj�8�=�����=��u�3궽�y�=���=��Ȼn��������㼫�ܼ1�+�6*�=�˫�������<���;���=M�+=���=��Z���ʽ�µ���ɼm��碽�-?;�ۖ�dh�:~>�נ����8d)���=̾>���R���uY=''�=��M=-x��_���~�=|'=�|���N�,=Y`¼��=�Լ��=�j����O<��߽:��<��=�L�;�{=b<�= �^�xɼ�-=t�1��cu���3���<�u��6穼��=������ݐQ>���=�H��	�ԼJ�=I�$>�=-t�=nM0>~L#<��I����;KJ�=��x�v����Z�;�'>��+���l<�����U=!�	��Z,w=p�f�.{�:R��;����{>�`=s�J��q����6��O� �?h=?���.�� ='��=�k�t`�b�/��wL�w��O��t�=���[�=�9�l���;#�WýS��<��� Y?����<o\���?�P�"�^O,��l�Q��=���<1� ;���=J=�>��w�g�<>�;J<�ʚ<��">m�;������=ػ��d>.8��x��=z���D�y�~赽����=`�!=gq4��f}�Q)=Z8>8>����Gs��Rν�筼6�=a�1��T���6=�����V<���ص�o����.�=��=y �=����T3�=Ֆ�<�W�=ڎ�<!w<>���<}�Y��J�c�N>Ҧ�=��������h�=�=d]�<(�̽8�<��Z���C�����CK� ��=���vg��'��{��<�s�;d�=�U�=�0N<k5 ��H?>^���S���lo��#o9��J�;���:G�=P�P:�7ǽit<]R+=�Y/��a\=��1=Z�!=��˼��~���K`�%}�=#6��\������=3�Ǽ�ّ���%��m:���<�m���<v�e<n2μD=	�������cb�B)�=-��<�nA=��S�Wh�=JQI==�抽�n,����=�6�����N=��>�	��O���@"��~�<cn&=��X=)�)~<<��>�j0>�x�<'���4/<]������=}?v� )G���>�v�����=p͓�E"����f; �T�<�-
��kM�����3=>���<d���4=�I½,��=�/g<)v���Oo=ܓc����<�uV�n�|;ᬲ��"���I��KO�=-�F=�ﰽ�#>C�=Mו<�����㱽	��:�2q�4=M�\;0��Ω(=|�<*ק=����Tݰ=�<� �r��:S���Ͻ���<���4�r=�˂=P��:�3��KO�`�U�v���	����}�<,��<b����9�v����6�=*��iLȽ◹��W�<��<$��M,�~
�=�Ń���N���&m<#����V����=��I=`��=ڡ6�l
��+ֻH+�=,���kS�%�><"�2�R7��=���=��Eb%=�<��>W~28��h=�!>���=�t ����=
LW��s�=����C[�v��=����j�;q�8�4ZD�!iC>��A��{c<��W>d�ƽ��'<��=Ξj=���=8ߩ=uP�<[v���mD=�c<h>)�='�����w=�t�=k��ay˽�g=yk���o=lb��=p&'=-(���;R?���=�����.���=���#YŽ�	�X�p�d�/��s�9�b���>�G$=���=i2G�-��8
(�W�����;ɢ��j�=��>=�=���;������5mҽ����˟=�9Q�>�;>�@ <�c�&1�=�9ټ��<�_7���0=���<Gjp�b�K���н�����|>�?7���>��@�@i=j��?�=�ۦ=Q0��	*=��6>mֽ���=U��<�H(=HU�� �;�R�<)�=��ؽ+��=7A]<�������9_4߼���<dV��JG�!vj=JE���=��<ŐW=�����uA���L�=yE�=�;�/$<�!���8�<	=*���IS���=�XT����<5+��YLD��%�=���=�,����aF��H>�F>p�?=�a=/e���=腄=<o=��=ip�=�/��C�����=j�myf���U<�L�=��>{{ ���X]�=�G�<�M�=M��	�0=^�;���=$d�=���=^d�=C�C!<=�	>��<2��;�%���eQ=�bF���׼�i5��E��0�?<_}�hy׼ރ���-ʼ������C>Y��Y�hte=�+���_���
�����FJ<�T=���;�|��7�=mP����=���=�Z;�������6��>\E4��!��W����r���.�=qc >8~&= �=5�I=<��'�p��a�=8����4j���A�n%=R�[="��\a=��<��L>�Փ�V;:Q����=?f=��R���2>�[�=&]�=p�� �E��=��=��6�	;��e3)>1�=��+�b�<D|��R�=y��<�%�<�ӱ< 8޽��z������=���%�=&�%���(�v8������O̷��ױ��X�<$�'��SY=d���-��Aڔ�����\�Ԃ/��tｗ|=(l޽��b=!�;�q���Y��6ں��üy��= ��=t`e������Z�܁(>��Ҽ����3����ȣ�������!�l<��ֽ�>y��=a[�=�����N>��=�=���=!> �x��p�<�?M����G��=<��=ḑ;H�"����<��<)Zf�};>F���CὝKn<{~N��o~�!1t=�y<��)=��@<�!���n�:��'=��Q>�M^�9	�=��%=$U��&���7T�O���W��󻡪!=©2���h=rJ�=i4�<`ϓ=$4V��:�9����=C�e��OS��Ž�͆=��P��2&�8�	�LRD�7Cd���<P>`M�=j=>�#��2�=���:Nx����=�Q�;s3<7'�=Hh/�o�K�<	�Ž�6�=1o�����`��&���e=�J��f9��Ή=�jp=���=,�P�L��=�����0,��d��Ϟ��o�%,n�h�=}M���<nЏ�Ix(�n�W=���=��5��ҽ�I⺉����==��t�O��=!��=�t�=����Ǟ<����P��=.�@>E�=�ِ=��<���=�؉��q:�7�|W�=�N`=P�	;�>�G+<�/��[i=Rb�<�h2<$�����<���<��!=E�=R>�˽�v�"}�<��<=)��=��D=�T.�0�$>d�$����,=��>U�=��~=Ķ�=ơ3�-+��.�=vѽ�'>*�� ����=`ȧ�{�(>��y=U�A=�=��"���=G�i�:3�4I������)>��1=���=�ʤ<�ƹ���7򖽫�����>`Ɉ�вA>�SL�� p��#����=b޽=#�t;CS��霯=SI�<��#�_�Ž�0Ͻ���=ͽ<t@.<���d��=j�=�h&=~������=8pZ�C�����=�:�=�1!��	����b��󼽈Լ��=��B>��=�[�=�I��ZM>�=>n�3�ɽOn�����vY�=W�4�+�=r+<@�Y=s&���XV��@��Y�z=����<�;=�g!>���HC#�?^�<+m���������j�;<�ؽ�P�:]������ӆ��%8<_P�<�/`�*Ï�2��=�q���]<�>���=A9�:��8�=����S߼x0%�:g;S�,�T[=#�</Q�<Ip=缼>��KV�=(2�M��<��g��V�c>�rV=���=�j=Q缳��.�8�.R>���@=B���?ȯ</��=��g�'=L�=:j=,V�jW�=gN�^<|(>�\�/����=�%�=Ro�=-���aaa�q�M����<+BK>1:��u�<��8<�޴=z�>�b�<uTT�N��=�T,���b>���=�.x��'=ಕ�g+0=�V���Q��N���R�>Uc=D�g=rpo�%�=F�C>ԂP<�4��"̇=��l=��"���<��G=h�=�'�;��㽓�=3�<=
�-`=��>q�`=�2_�_�@��.ν|q�sOV�g�'>c0����0�6c��
���vm|�� w=�Fr>�
>�������׵;�֙��Z=���=]���T�n��i$={�=f,0���m�����V�h�F���C����=H�B=R9�<�E=x�(=���=�"�<w�:<gl�@A=�a�	�u�iy�<8��=3$�^}]=���=Xڸ��V�=����2'=?�u��e�(߾=�w�=������=�N	�[0� ��/���
=��<Φt=�����j_=Ĵ�=���=�����1�=od<��r=6��gz�=oѯ=X���� ���������2F<��=�.�=�p8:�V����ýl2�����=��	>���<��ݽ���=1��;�e�.s�l�2<��=��껩�L�Ǫ��r�=ڬ�=�S�=�v��	��=�"=vnؽRV?���'�Ip����=�u.�Tt�=H�=�+#���:�g���O>y�Q���=u+�=��$���"�[-����,<]y��%=��q��lGA�Sҷ=|>�2���X�=)��#�=�hɼ�C�����cdM=�>h�<m({��=��ޮ�	�J=.�ۼ�z�<�7=If�=�b�=���Qwz��9���	�����=R���؝�?$�<���Qͻ׌�=���=K��bd\�p�-��x�=m�=�k�=+��=�'=Y��u@<�$a;=_Dd��-���>"����4�KQ.��=�=�G3=�UV����=��1�ٴ>�u�=���<i�ͽd7���l2=�� >�٦�^re�$}�����<ž�<}�>��׼u����vH�,yɽ<]�=j�/=�}\��#<�$��A=VT���⽌�=ŧJ�(��0c��0��}�;_�*�Z�#=-ɽ�C����Ž�Q�=[T��]#f���b���ʻ�'>�	="�i�G���5�=$��<��݋���}-= �ֽ��6=���<"i�=������7=���@��=vT3��伧�׼�H�*--=��u=&��n������<U��,��Ŷ�+�u�2�<"��q���H�vX��ȉ����]>��ܼ�C�=�S��*��Hv >���қ�<�����=R
">f���!>���}ɗ��v�<m2Z;D�W=tq���N��H�-�w�=�/���	�s�
=S�=��+�#���=�=�{˻��>��:��o���i�Q>G��=�qR<^r���J>_Y�&i�!~w��Z�=d^����޽���]�<�X��=�+=Ϟ�=W}M=n�`�G!�=����F��.u�=��B��ý{!�<����C�=|��=�F=L�=DE�&�
=����a��O�><����p��;����Q�=$�H��<@񙺭 �	�[���<Z?F>�h=����T�=���<�yX=
g���l��n�<2��cG�������N�z=񧄽���Ѱs��7%�qx]=�%�>MGB<c�5���:�Xe=Cb5�Z�=�>� �͏'<_��='U�=��;��=M�>��@�y�=��>ć=�
=Iə��l=7�=�+��a�<^�=����a�9��XO9�>)�@pV=���=Us<��B=�����9>Q><y��=��T<�:�;õ=-r�:��<`�4��Y>�u��6�ýqk<�x�<9=ฺ<�wX�^=�5�G导XM?�i�b=*�b=� >4�����<i�ϋ�� �;ykB=�Ǝ�|�4�JdԽ2X#����=�>V�8<�5��.���t<��<��
<\&>����:>c�g;ϵ_�B1W=^�<'�|=I�۽�=Y٬�`�t<O<�<e�0=XO>A��=���gY��K�9=�ޣ=o%�=�=����I;���l�<C�=�6�}6˻����W�|�[�x���{�<�ݸ�w�� 7<�/s�f+���e���=c�=<����lP��U1��?@�5��<�"���ɽI`=yX=���=��ȽR�T=�<���j��fܽ�W�=%tĽ&�(��6=|�c<� k='��=�33��{�;RCv��!�=[O<GJ��;j�ٟ�<�蛽d���7G��Oo>���<0@]<v�=�4=H����)=�U��{��_�=����5/��f6������3=�[>.����꼆K�:d��<���<c<G��<7�>&s>�R��z���Z=��2=)|���|=�	->P�[=��s=wM�;��;�S'���Z ����=���j<��1=�ʕ:n9x={ԟ�@~7�u:�s:>�'Ͻiڽ/Sw��	ڽm�%>��<�����<nXǽ_P9��<�<���T4��ʼv92=X~
�u�#=_��=�=�����#>�=]���=��=½�Sn��w=��%��'ɽ�N�<�ا=�U=5g�vi6=��ü"e�����n�]� ��<g:9>&�N�u,�4�����<�T�=���.�>{�,�΃7��9U�D�
>�<'�:8Q=��=�����9�0=�6=5N��g��<�sl�X�&\Z�E���M���=\��:�x+��g&=��
�(�=��m�=$�z��N_<w�=������=�zi=���=��-��)Q�Ad����=�	<h�������k�<0�ʽ��F<`s�䰽�w�={�>�<-�!=�I>E�<s)�'����	���<�D���}<!�%<͹<\O��F<0����*�Y�>��=��=yӺ<�#=&S=b�l�=Xd==a�=�_>%.�<�A�=��n=�q<��=�ݥ=4��=x"y=�,l���<l��Ɍ���=&
>�{v=��!�=�E=�Ð��к���J�=��;�$:=�v�=�m�=qg>XQ���l=�X�R=RZ�<�ѽh��=)?c=HѠ=�X���<�'�;kc�=FVb=IG�=����*o=�ƚC�IU=��{=��=hmL����=]�4>�U�<���|lO���=��-�ta�=k���TJ=k�L=����ZD��)�>f��=��<���=U�D��O�=*��b����d<��\��Y^=A>�=­���bb=�;+
�<<'>1�W���N�d(��]p=z\���wD<B!>O?j�zK-=9ș=���=�ý
�>ik�<�
Y<\���<����=���=D��T��" ��EY��K[�<��P�������=v�=	=%�=���<�L�=O�>�7�y#���2<->�=�F=��<�6�=�U=ze�=���v���2?k����
9�=�N�=�^�=��<8��=�5�=���<��$�
�|=Q�� t=?�=cg0��4�=
������=��o�_=)�>���=(�E��� �≀>�vl=X!>���%���O�-�>5z��WQ�,׺��H�C�=�O�=.��8���s�=*��zY�<
?;-,ݽ�V�=y�>��C��;��M�l7��'��<:��A�Ռ=!�\;^�N=�P��H3�>�NE�_�a=G;|���½0����]=`"R=����ڴ<���<*,���:=c�=�ǃ/=.j�<�0�f6��;n>�9-��=m�������9��=̼�ă=�37=�F=f$���^G�AQg�3z�(���=%]�<��w��p]�<>0@�QnŽP��=��
>;�=��<>��$<�=th>:�����T꽿�=��<�W>�0?<�FK�L����N������Q�=�=���Tb=�k>=�.�=��+������=!��|8���i=[��=�9�=o�.=�忼&�ԽCK=~����=�>Z�M<�@�1����|2>%�=�+B�4�7=xϮ=���h�=L�>q��:�p4=���<�9=�V�;|S��>�g8����=饳���<<s(�<$��=qֹ=�=�<༏��$�;�f�:/���%�B�ȼ�|<�`�*6<r0�Q������=^q�<`�4���f��d�=��<}v�=8/�A]����="�����q<(܉<���<�F>�N�;R�&��=�<=Wv��{=X���E%����=��6���=��2o�=��T�8�ӽƆ>���=�H�<A&��I�z=f'7��pG=Ċƽ1d=�o=���=��<���=��}��=��	�;�<�]A=xI��!�T=��߽�>��I�Z�l;��3��z{=�.^=�K�=x+�=��C�@\����<nҚ=�/>��o�����
��o��;��ս�z=�	�<�>��	��9��s���fh�c�м0t=Qɱ������̬=:R�����<�J=�z���->��P�^/�<��	�D�G�$<�=��żdg��\��=��=�fҼ�}��SU#�M��=��;���t��M;Ze��=��	>7q���ٯ��a=��>>l��q)=g��:ؚ��`������<��=�*�=[ʽ>N={�;�>��l: .�-7=��=�E8�~�)=�(/<�j=�pu<�z��pݽu��0Ň=ӯ���E-:�f<�~����b��y�
�2=Y�=��=�4�m<��=���4@;=���է�ͯ��>��>^�t��2�=:e��9L=?ۂ<dљ�\I>�
�	�x�o��=4"�<9�����<3S��3H�?��=2"�Q��0d����<n=���;���ߌ���	?;&�\=���=n'�=�_=,�=-�$�!�ܼ��꟧=;�C<F�>y��4�=W�v����<P��᫼�ν�ϼk��=�U=/�6�D�4<�<��= ��Kmf������k�\`�M}>@��=�ߠ�Ӊ
���Ƚ��<�#��G��q:ּ�����x>s�	>��=RH�=]@;�G���>�(�=r���C=���=�K�� =����M�=^Y�=]��jX=�S��	z���㣼W������=w�ļ�,��[��+S�=����I]��_U�o�#��M����A=�
��L�<=옠=�Ȳ�	Ȕ=��d<|g���S>x��eʽ0({<�A�;q^������������=��<��=^�c�[P�]ػ�r�=ǹ�=�������H,���?3�-�=n~���9�;�%>�>��j���9[�(=ݙҼ[܀�~Tƻ�vM=���.ր���=�wI=�u��#u���l�r�<B╽�p��NY���g>;n=�41=�U���&S�V�=�">��>����nq-<bT<��<�ܽ��<�O�=�	�����*)><��;�q���ֽ=�=�_y=`�	Ј������5�<G(=9��=)9�h��&�=��|���(>5��Ra��Yi�C�I=7ͱ��5�=�<�=R�8=�3 <�گ�k��9s1�pH��	_>)v�Y�N�B"=ԟ�w[�,O��E��x4>�L��R
�!��ȅ=ǣ	>5��ɷ��S���h5�^Ȁ=�Z,�܉�Da�ފ@��S>zg8=���=gњ<��P�yS�=�(,�X�<b�H���� �#��Yf��}=CsP=�HѸ.�H=����P[�=V��ۆu��﮽8a[<�d>�m=b�=L��;�%�������DuH=����I(~�#x�=�-U=��>6L��R��=���=�*T>*"��0I>[}��_ԑ=�����PX<��u��j�<�Tν��(�"�=�%">t�X�^X��a�=��F���<p׷���R�1���-6L��&��q�=�/��#�=������#� >�j�=L��=P�">�Pۼ�_ܽ��Ҽ�(9=eR����>�A[���w<�y<�н������=�Y�=X@��Aڽ���b�<�K-�꒲��
�=��<�G�=�f>B��=��0�[ם9K�{��=Aa�=�b=�"D�4�=�l���+9Ξ]=X��<&�=���/������=�
m�{���Ľ�Uҽ?A�=�>������)�i�����"�%�=����F� >�� ��+�Iy����=������<�?=�����?�=fǔ;�;�%�>�U�Mw=X�=U]��)=P����dZ=N��<#Ey=8u���?@��ݽ\,���h=�5)=y>���D;/R�Y�(�Z��=l�����=� ���<���;ą�=)�f��3���&��S=}c�=���Ğ�4Զ�1�r<��M�`�m4�=6�G�8di�Q}�����.��< NW=�G�:�T��Vś<�	C=�e�4׫����=���^��=���;� �<�;=J,�=��=����k=�?M=��Y��4<=�g�=��b=��$���l�S0;;NM ���~��#��y���Q2=�w=+���۱<P�=(�Z<�N��Ӿ ��<k>��<�s=��=QZ#������=�Ң=��<!#�=��=5�|=�w��4��=�9%>��=T �=Tlɽ�=jF�=���=�ۏ=k�d<>F�l�Ż������d=1�%>�b��U��<�p@�y�{=�C���볽eD�=��.�~���3��T=�~�=�J2��ռ5>u>\��=B�T����
=Sߧ�����⪽x��;k��;�<L�=��^=��a��=������R���
��?�=Eva���;�	�=lk>!�#3D=�>M�:��|u=v��=s[�=g��/�=uW<OX�=��ݽ�W�<-�> �ڼ�B�;�#=M*\<��<fu���ѽ��+= .�W�;F��i���K��bO�k�<bNO�)v�=��2<�����寽-&	>�7>������G<[ x=�Ƚ��C=*p�<&z�^������=E<���=�=����>�D�5�6=�j����P�"�hE>�@�<���=.�;�=vrT� �<~ӂ<KýH�*�����2=��+>]����W7=�6˽���=�(�<4�<�<m=Dc=y��0=�=���:z��<92�=%�=���
G��g�;�M���>6��=gǮ��(=/b��M�Cu�=�m���L�SI9��9��==!��=Oxl=` >X=�mO�@`���{=�߼��=nϘ�m漰D#=1��<]�=��=�e�= ������<D]�<�I�=z׽z���(�d����=R�>�65>{�V�o���� =��g�= 
��vS>Gq�<�Ԕ=��>g������iU��T�<o8�<<V�<��V;|釽�=�=qQ��R��= yh>vl����=�`ýne�=������L=6���ˎ��-^��q��I�z���/�<�S=N��=�f;� �F|�� �4<��7��;�Ի"�<��=%�o=]^/���=~�;�Ў=��R�=Ky��*����`='���'DŽ���=0��į��P.�_�6=����׎=��%>�Ĳ<�Dh����=���s粼P��=���:�!���;��>�=�M.�Rٵ����=��r;��;]|�=�D�=��%�ì�=$Q>�3�=�Y�F�<��P<���}
�<(���%���m�6���e>��=��M�h~�=%>`+�����<Q^�z��;��<<R�<:��w@��Bjs����� R�=��=��=��$��Z:�%�=�G;��ƽ��/=U��;��k�9�H=�׼����!�0������I�����=�.�<��|�2�o�Ƌ�;���U*q=Z�����<'o�<
0c=4�'<
=`n��3i=x��<xh�<���<ێS=�K���0�� �>�4	�ˍ�=:e{�z�P=H(��{��U�;̎.='������蜑���5=ZH>���Cx�:^�ʽEx��ٝ�=�]���SP�F|Z=�:|��<+�&��/:>+] =�Nݽ�ݖ� g��Dz���s
<	ʺ=��=.�ĸ�<����q�M��>1�R<�� =a�	=baD=B�ϼ��	=��<>,{="�ང����R��携�Cp�WF9=�@�������<Ό�=�﫼%��`o\=8�?=rR���0�<�w��_�=�����=��O�Ж�=~�=Rz�=r�V= r=��>���<<��1�9���"p�=�4��F�=��C=r�'�r3>ރ�=�;� ��e<�a��<�F=�1=8��<S�z���o��<))=0�����=��P<~�=��5�󝰽��h����>��)�oz�=r�+>�k7>��.����n���=��e�$�SZu����Z'�=|F�=+���5���r� -�>_5>�｡�>r��=r�+�5�ؽl}=�F+�کƻ*��<T~��J��?��<��1��(�Y��3���Š���.��d�<�Iv=���=�Dȼ!�����=�:@� �ɽ��#��=)�<CN���뎽y�=�v�;�ꑽ��]=��
��nY>!�=�e�;�D��LQ�����<��<Tmg�̪=�h#��f>�H��j����=D�۽`.�=�i��� ޽�Y��ld��o���U�Q��K=p�U;�y���`μ]=z;����֧=FT>�I>h-��܋�=W�z����=�3��,=����n�ͽ <����+S�=y�3>��M�5=�y>�u���A<W㘽�x�=9#A��x5�[v��Ͼ�=>�=D >��:<E��=6�ӽ��>6Ʋ=�蟽�P�+�<v��ެ=V��=�z�=-C��ټ��U���=��~�tƼ>EA���<j۹��鉽,H1<�w�>�&�Q8�=�㠽�H<�"����}�<D{	=�?�=�ǽD�>�ŗ�"�d�y ���~�;M>�=��s=Qu>�k=�3�=���<;�#=���=����X��n�����=,h�� ��86�=�)1�n��=,v�h�><n�=- >�y�=15��}ʚ=���=��.�p=S�<�P��*]�I��=�C���ʟ=��=I���<��=;ō=�=��_=�v�;����_X��#�=ea?=X;K�Ǻ3k'��43��L�=��A��"�=�&�Uyf�����2F�0�<T`'=Kd�Dӽ�]�=���1�>�ƽ��ý���:��x0���̽���;bf��J��A�G9>���ƽ�!��\��<�I=zvw���V��<�w`���><D�Ƚ�"��V�5D�<a�ҽ~玽�r	����=�OM=�i�+��=�=r����=���=���ܡ̽yC�=k)���=�=�C�=����D餽�/�<v��<kꟽ$���G�H�Y�_� ���=d��<���<���=���=�3��	�=M����׽�d;���;�ɹ��=^�RT?>$J�<R|���^<]��=�?I��(>�ؽ&�d����"J��L�=��_=����N��n��=5�>x�m<<�<A�=c��=��<G=ʚG�Lhs;<gj=�<2=�=Ny<�@)>�'G�N�J=;5>��J�!ƽdr���?�=����6
�����]z`�:�6��T �M��=�%�R��;h�=���%������y��=�0���>�����:��a�=�}Ľ��(����=��=��=��5�nyR<��=՛�dp������5�+p�<���=���=	]f�(�ν|{��>\�A�=����1�=o�X����=���=�H|����;8�<���s��< ��;[����m=�4u=q�}<R���݋o����=g6>Ek7���n=���Ϝ=�?�=m��-��=�2�Ws��Ab=��V�iQ�=���<�g�=�ڽC�%>ܽ�=� ߽��=��G��]>���=�Ă�k]�=a{:=�a8�&Jn=��^=�RN<}�P=%�P�`�JB�<I�J�NU����=��<�B��<�Y�T'�=0H=�g�=��=�~F;��p=�<W�E����<��ڽ�.�4��=2�B=�a���,><v�<�\==�'?<���af=ȁ��ļ�l%�l�l���>RY�<T�۽�7=���=F�4���@=?<��#���m�H��2���t=:�1>s?(<N_O�&����'=����#>զ�<�s���� ��<�/w��F,�Z-�=E�<'P ��`�� �=���=�8<r��=�=�rVF�*��<���=��<�� �,��=�<"<����ʣ<��
>�r������.c�|�<�W=z�=�[�=-�r=�]���<	b���
�<�5<��!�=���<���;W72�+��:�;�=y�=�j�=LC�<����yڑ<%G/=\[߽�$μ�FN<$w�=��=}���a�W�`�=�-�����"��:�o��=ߒ�=۽򐅻W�B����<�>m�G=����č�<C�㺞�=��Y=/a�8�r<V[=��:��*9�ƺ>q+=eM	�r��N��~;&��p�;��0=�qc��2&�a"%>������	�7<��н$h�=�b��M� �q��헋�"�)����=9a-=V����H���-=/���l<e}�AQ�<'_	;�üz���`�<�!뽜�>#��=/
=�u>�	��|�U���\�=Sԕ=,��;�7��9=�<��L=	*#�}�G<���}����1>g���겴�׶��"�>$�k=](=�p�x� ���߻7'�=Yu�Ȓ^��y$>�l�js>�<�f�<�誽桊=[צ=_p���鏽�B����>>�����S>��&����zb9='�����=�~�5��=[�E<�㱽Ms>;\�[��ð=�� ��1{���?�~Ȃ<�K���i=:�����]���=j=~��=\���7O>Grq=\`���(-��X>Cu�<��=؃��&�=�G�R�=뮽l��<�*���CZ=<g�����=ࢨ����;>5=A�=���������M��=��\��E¼-x�=��v=R�=�,<��<�95>Ɖ<xm����j��x�<9r���i�&"��l�������DGҼ�ż8Y<�k�<]��;�������=�S（�߃����<��=`PA=�N����=��)�K�q<��<"��=���<�$����<DΔ<��h��>B<�9>�z=��u<!F�=i=<���=+A��Q����3�풣���ڽ�%��Oݻ0�u=��=���W��'��j�=ƽ{���>^�9�$���6�<�����n$=�*��	]>
�Ž�̡=)圽�}�=SM�~˻�#��=�5�=l��Ú;<�n=���<a!1��R>�B$;r}�=!]��+���q�Y>��%�6�u=�Z�=��=���k�='��֕�=��{=�>���=��d������ˆ<�aM=A��|��=z�:�D��갽������Ž�"�y��;�T[���#><�%<�+{�ʍs��xJ>��X=�[=���*��j6.=�n�<����TN;�q>׳�����=E<6ܚ�t�3�)x,=������=�>�z$���=0%�=��=-�=�5�����~���ay�=�+x��
_<j�=�ʳ=tۜ���^�ĭ�=�ך�t��<j���#j׽��^=��{�l	[�)_����[��[<��=)�Z�3һ�D':��!=:'>�6A<��/�
��=W��<M9���=���<M�=���=��=�]�<�虼�:�9�=@�!=|�=�{�=ا;�ߥ=���=����?>���=֎Ȼy����>S1+>X>tX�=ט�<����E�l=��ϼi�=���=bA�=.e����닻48$;e_�=c�=����r��5����%���|��	;=��=C�����������T�=G�C�{v�=�ܼ��,��Y;��E!���~=��=6QT�%SX;�h �@=�^�%>R�=�_�,f|=Z�=c=y˽CS�=2�ֽS�4>�W=]���� �<�������=~t�j���� .=6�>P~��4�=��1�r%�����=2R��䣓�Ї<X�^<�>�%U��"�;%>���<0i��Ϻ�=q���ƍ��W���j�ʅ�<����w0@=#~ <,lO;���<Y�=���=�(=,��P���Go���C��Z�=�<�U=�i�<S�ôƽE��=��[�5�*<;~��Е�<��ѽ̃�=���=��ݽU��<�F�_��\R�=t䐽�ޕ���M�h�<�!��=�\?�en��W���uOb=9 >Ҏ*�y�J�f,�<n��+*=Z�!�Y�W>��R�3uֻJ	�~N���ة<M0��f� ��s�<x��4 �=����}mc=���=ꨰ<��½���o&s���=^AX�S��=������ɽ��Ž]>���/�=��2��0A��{�J� =�m�1�	>�s�=�w�=��]=� <J�@���/>/xt�k3[=���<Og�?O�<T �/���|3=������>�6<՟�<À>������½d�>)wB���}��)S='�"c�<Gf>RK:=Yظ;\ <�4�=cƽ�����J>�eP��Ӽ4+���f=.���/���Xw>��&�eA�=�a��w ��	ڜ�W�����#>��^e!<^N<�{<���=#��=X�L��]�=[����(���[�<�j�=!	Q=�\罂̞<�U=��=c8��%&�=�CT=�Y���H=����y�(��2$�Rj=	���m^����6%_<}H�;�z=c:�!���T��S�ϼ&��|�=���|�x=�Hu�۷<h�ý���=5!o��|�=D�"���ʽĥ8<s�>�o�<J���u�=���������=��=(	�<A8�=:د=}n�fEn>]3�<��7>�w���üc�0=�ˀ=E���u�x<\��<\� ��Յ���t�����5<�Y=c$��9L��ʀ=�<�<�d��fT+��ԩ<��Z=ZĪ<�!,<D&>�=�����S��<��= b��2n>�Б�P��<��=���=�=��;O�м���=ӯT����=���<C���X������>���=�p�Ds=�%�=%��ͦ�=m�ɽ���=�گ<�:=���<�+�Z���
�=󏻼��h�0�=�?�=��>��;ֆ�=�a��}�<��ʽH��=�oq���(<��=�~�=ni��Ǣ���=h&���O=w�ټ6�-=�f<}轤�>3�(��"Ž��H�F�>���������;���<����ٜ¼T#(�8N��M�<��=�k�=�[�=@l_��!a�I:�<�Pp�j^=�G$�WC�=PK�=�>e�ʼm�;=��=s1�!�=e&�<!�>>�Zi:��T=������J=�I��=彅����; <��=CZ�=d`��%�=k{;h��[�����6��Y�=���қ�����{�BϿ�v� =�0���D=�
=���&3�.�<%'ٽt��%ȼ�]����<9R�=՛@=��;C�;�o>�	�=
ѻ��#^�<3�=sYy<��l:�#����<Q��%�����7=s,��W>1]�=,g=1gʽ�N��ܽF�n�W=1G����*t<Uhý!��ߨ��U�=��U>��!(�=]���"�e�&,"=�?��7�?9�<S$�A�W=4�<O��=\`s� �!��@�<��$� �Z�[=�=���=��=������=��%>	��o!��[. =z��*l������.>b*>���=ҙ<� ��&�>h�;m�f���>��w�'1��z����=��>�0��4�7=�`�=~&2=��N�`�>n�,�F��b1�<G�4���g=���*b�;)K�<:���=y��=� w==]�<F���N�Av�=kkO�<E_�����`}�?��<F_9�&y�k~q���5����������=DmW���<`�c�[����='U�-:�=�i=��;#���н=���C�=",�<Z��O{�D0<,<=�7ս�QC=֌����z��=�����$��8?T�3���q���>�#=?LؽvC[>���<iA~<��>��>5���eg���>�@k�.��=Rю�o�*�0WM<O��<t�<�`��E�<0z|�Qi:>u�@�*�=�<������=SS����<,]��=o-o=숐=�1�n�Ǽ���=���;0�=�=��0/3=j�\=F
彸��=
�ڼ۹�:@��;���<�ڔ=v<OT�=�$��P���G�V=�&�=�Dк2�<�f����<���< \>T��=Lf�=�^L�#��_$>#��=e��v�e=�|A=M��ƔȽ�$��>�.����<骿���<�
=P��<�o9=���='�2=��p=��=S��=�N��ڽ��=��=�'��`�=]{�����ȹ���`Ľ9tn��GK��=ս<�3�l;v;>A��n�<g��=� �=��R�=�=�y�y�3<�ز��l���o=۪=g">zޠ��;<�)>�M�=��;�U���]>��_�U����8���F=&�%6� �=�4T���W��L<�r�b%��.���<��1IX������<2=<H�rhv<K���!A�2�0�ќS<ê��]4�:{ Ƚ�|�I_�=���<n�>�[�H��s.>�<_nн$ߨ�_�D�:VȽ3	�{��=ĺq<&�;BR�=�Aa<��/=O��=�#=���<{��U�1=3o.=S��`䴽���q<�=�� =�O��1߽6�>��~�bmQ��g>u��Mcս*�(�f,)�!f>`�U��AW��P�=����|�}՘�;��=ǫ>ڠ=��R=��<�숽��ڧ�=K��5�E��"�=;���=J笽�V<�c�=E���7=��<ZB���ƽ��=x�<]��:/=z:&�U�=Q�6�����뮼��6='�\�O�x<�0>�b½��e��<�Pݽ��>T(�=�ZJ�G+=��D=;)��4><A�=&]
��%½�һ<3���نG<X�6�F2�ͼG=)2����~jR=6�=\h��Qh7�i�3�ʈ8��#�Q:�=՜�����<����J���?>5�`�eW��\&>�T>��0=��&��j��BU��>�aϽ��W=R���֏���F=0�����׽�u��V3V�}�g����=��t��=� w���`=%�m=Lt'������4=�Dἷ�߽V�=|��<7D��#}���&<�_λ�-< f!<0H;�_=7<�1�<S>l�>q�
��; �+M<=�1���.��<+���*�=�,i=1���e��p{��ԽB��e��T�=@���F9=�����\�K��=>1����=LM=0Z����=�F����'�::ּ�;�
��<�<�|�Q���j�������<�݊=�<"=�����,Ƚ�g�C=\g����vi�q6=x�=��<R�(���:����A.�<�w����;�V��F�`�j+=��=�H=�&`;i��>Q�=6E�����=��=�z3���<���;RF�<x>�q�h��=|�r=ׅ����HT.=u4=L���`���5���2H=���=3H�R.��k�=��Ƽ��#>��l�A�=|�g��S���U>�F0�h�=�0=c��=�L,>��=�_�=$Y��Lܽ��*<P?�<V+�=��!<u����5=�J��o����:>��#<C��<��`���=��0�`wf=3�=l�I����fY����=U
B=G�>���=y�F�< �	>];�Ka=po5=d��6��������t9O#�<$�ƻo%=S׌=)Ui��=4> V����H�=��9>غ;�+=;е�=`6�<_>2�6=]z�=���=[�н�f�=M�d��E� >� =���=�N`�\����&���/�r����׽�T=�%�=�v6����=��j��p�&�1��DV�=e�<��7<tnD< 9j�	��=c�=�8u=��=���5�=��J��f���=��'>���=���=��¼�v�=�c�=�ߝ��T=!�<=#4�Sم=F�����mw= �}= '�<X%���=s�<c�/�&�����`= �t������n�����E��H��=����J(=ӊ�����k�
�����'���6�qG�=����[>vFQ�"R��O#��dI�<�[<۔�=Im�n��} Խ��=ғ�DYG=>L�=��>Ĵ�=�i�=w޽�G�=�ۼ}�ƽ���~nb=<�K=���G��=i��kh�=��=�b��,�<��>��h�� �9@�`��,�'�Ľ8ݽ	�*=s3T�n`�=�Fμ�ٽ�̬=��<�T=~A=c<�ܴ�=g�̼NiZ�B�D=FU�<���=Z�����<�+A=l?��O`���=0u�yL6�/9�a8����wǂ�G��<��z���T�=_����_�lPY�
V�=ph�������>ݟ�=��ѽ���{��=��=StQ�8��=IlB=F��=CS>���� ��=էw=S�-��μ8��=q�N=]K<��災��#���d�]= N�=�!	� 9=��/<���7%�ި��<�Ga�=�9��ǿl�F4�<�z�<�E��`����=���ꋳ�si�����<+�)�{Z���<���=G�g�G�Q=>�T=������=p>�=*��=\�H���U�:o.>_�0=���|�>g@�=�vD=z�r�F� � _�<�
�W�A=�(�6�_>��=i��<�+z=�*���]=PQԽ���=o�&���8yqO<�ʭ�mg��	 ����$0ܽ���=/��Q� ���)�� )>+]=����hޫ<2�
;~J�<u"�}k	>��;���=#��j=�=�����9A>g�=�=Esy�U#��E�<�=*Ҧ=}�ۼ��<��=^[*<։t�MJ
=��h�/��=j@ܽʓ=$>���=�߽���=�y<Eg¼� ��ly=5�>����%��v��X����������5>ɹ?���V�`��=_M�<c�a=(�nz �5�2<23?<���=fxʽ4�̻:ӓ���=I@��`<\��fL=��{aR=��<M	H:��0�{:>��c�>#��=�(�=�=�=K)�<���<�e<+t�_
 >9��r ���0�<Àb�^l�=f�ƽ
����w�:�7\C��c8=/�*��텼�(��3�3=O�:���=\e�?੽,�=^@W�Şk���=�5�=�2�;��=�7��i�=P�p=��u�eS=��,:5@:?�����<�O�=\�>��=��;�	=�7��!�=��=ئ+=�2 =l�n<���=(=����6׼}ܖ���x�"Lۼ@����c==��/��ʻ�WD�e������V���	��+��=$���ؼ���?�>&��=&�c>� =xh��w۵��a�=��:��=^9J� �>=D�޽�V(��{ >���=��<+��=Iqq�BB��l������֏q<~��=�W�`e<<� >���=�J�'P�<A=<�������;�h���K �3��\��=�*�;y���%�R=#����׼H�H<�%=o��=Q������~'�p�A=;�M>���J]���_$>��+���<.���p� >���=�;D�ļlg��JP<r���QX��0�/�U�v�p>o��<7�/>@eX�r�a=Ɋ���A�<���="���K)=t�=R�K��G߽�q$<��$>#�=�]�=	��Oc�����E=�Ӎ<d�Y<@(.���c<I��W9��<!�>�"]"=�(�F,=L�-=���=0i�<ܨ����#=�&P<R� >J�ʼ�ʮ<�P|=$lA=��4���(m��P�=��;�Sx�������=^L�=����V�=��>����A�� e�<v�'=��н^� >��<!��=���<��=${��T��u�ύ���	��]
�>h=*~�����<,����l߃=�9<�5=1e8��R*=�Jg=s{�.����=�罺�xL>�4�<y�=~~A�sR)<�|n=0�⽨����"�6̽��=>G
�=!<>u��Gs<�E���D�j=w2�<[�~=��=#=i�Խ�96�f�R=�?�?/ٽt��=3�=dȮ<�\�s�;ฦ=�">��'=���=�ѡ�	O�=��7=��"=h��<|}9=��<�/�<��Z�yR�a��=��=i?����c�l�\��=��=$�==�-=�FP��@<g7�/Xý���3�ļN&>h҄<�H�'�E>S��<K�:���<���=��f<9�=�)`=���s�=��ὺ��<�>��8�^my�*�=�̼���˿Լ��E9�;;kƉ�*�`�v���!�%q>�Qϼ��еG=u���=�q����=�O��oe�;V�׽�9$�g�=���<B$���IK>O�_��ϼ��<��`���0<�����D���;j�<�0t>���p������<�K+=jr��UJ8>.�_>���<"�"=c���Z(�=㈤<L�}=ˠ=�Ψ=b&��,U��D��g暽p��<�%�>ǀj=�)��U=H��<ɻV-̽g}�����<y�=��<Ot >���VS��Ր=�ZH��G�=��Υ�[Wƽ��h��Q���o�;���=�~ҽ��������;2����=�}x���T=C�:]�ͽ�� �f\�="t�=6`p>���<�N=��q=�ѼW�-VB<	�X��;҆=T�<r��=j34;^z��A�=�h�=�\�{���ݽw=�v��	��=S�;h徽�e���魼�`	�# Z�y=��=�,<�-=mu1=�@=0c+=�h�h�n=V�ٽ�i=rci=�2$>�&�t�C<��B�~���b�=�w>���=���%+�:f���'�=����,��<̅k��(O���e!C���ӽ�t����-���<�r�y���S?=˒
���듁��ȇ�������d��>�z�;��==:��������F<���=�;S=?30��e=�ݼ�c�q�6�z'">���;hGǽ��9=��hmT�]$ ��˄=�Db>?7�<;O�=�a>���dI�= ��=z��`
������D<R	_�{��<���=I�Ȼ�R�<���<���=�q�<��=`{=���9~=��*>ި�<�ӽ�״�Sۡ����<�˽������3���+��ZսkW���5����Ut�=�ݙ<m�F=����l+=x�½�Yn=�Ն=���iu>���<|i=|1�z�ýJ9�ZI��]+���k=z�"<�O��H8= J�<g��<��7����=g}���>Q�}I���(�����<�� =x��=�">�qg<(ŽiR%=ɕ������ �=�ێ=�=#>QS>� Y=�Ԗ�'�Ƚi��=�A�:��3��=���3i�<���u�����<6#�=]5�,��=�C��>��/@<hB���Ƽ�n<��=p�<�����.�� T1�Y+0<:�7=�B��`[�'"������-������B�dsp=UI��	¸���=�ݼ��w=P��<�N�����Z����i�� =�=b"C���)<����J�*��=�5U��9=B*�������m<�D��<��=��S=�}�o�!���ͽͫؼv+�=�ٽ=��=	N��k}R>���8W�ʜ��	�¼^��=�䍺2uƽ{/ �q;F�������<3IA=�l��,㩽�(>h�6��O>���?��6��;�n/�|$��)��b;J+�=y>h�u�A�;'݄��2�=���=��$=�-��P>b=OA��=<��&>k��=-m�F?=jȔ=@��=��f=l�h�;l���"�xC��>�>=Q�����L����=s�I������Z<���=�S-�A�>�^�KL��9�9��=�G���%�=W�;��N>�	J���&�����>����R�=�|�<qm��ݎ���ý������`2>�>��^�YJU���=�Q,�ਢ=:ǳ<}��;��9�o��tm"=����Z	1��v =Bm�=e6�<O�a��뫼�. ���>�`��f=Q^�=�Պ��$�;K�p���S�bN�<a{�<����}�׈�{��;�$>=(���D��<.>C^%>���F�8���r��L0��k��GŽƘ%;.˾;am/=�\N��x������l�i<��>ڎ<��d<���=�|�V��4k=q٬=����/�$�>�nU=�3=p��>L%�ю6����=d	>��&�F�>V�=+�a=�>�A�5�A<���3����=��H�=wP��:+>���=��=Z��<Ι��n1����.�<T�~�߽�@>���<V��G�&;�=�=S7��)ڼ�W0��7ݽ�HͽWc>k��GĒ=�m�9�4�O�/�o���k3�;1\{�A��;#2i=����De�=�{�R)��tr=�&��D�Ū>Z:�=��;���V�=bP=ޜ%�6��=�g�SƤ<� w<[=Ny�W
>w�z��8v��^ƽ�W<u�=��<1�;k~�=ĉȽ{8�=?z.>�0Լ�����9=>J᛽�����0=�=������q�MԼ����*�=1۷��=	��&�ڻ�rS�*��=�<��{�>Qz"=y�=Խ^��H_�=Y�=����5�=���=�M>oj��R�W�;�>Գ5��Y(>q������=_7>�t*=_�<<��;�6*���=���=מ7=�����z��`�K�ོ����滯i<s�(���ӻ��߼c�g�[#�H�>��|= �컑��=84�������� >�;4��)>GVp=6̆=�w齼���P�ν���=���.��� �&=n�;��55=)]��i�v;t��=U��=JVԽ�s�=n�4=9�=�ڷ��Ņ��!;��I=Վ6�-�={��/�>j'>OĪ<�*�<i\����=�8<eZټk�a�`A�=�*ҽ*���b����Y�!Ἧ��;F���$`�S竽�E=�V�=O�=�8�<�RP������5��\���7��OV�<�+T=NXY=�;�=X�z�����՘���d�<xhؽ�<7=$%<Zu
��7	��=E��<��XjǼ܀=
g�8�<m�U<��2>y�ڼ�T<��̽���=Jǻs��wɼ����聽�ꮽ㖟�i��=D	��U�=1x��>ٶ���a<I��=�Z�����ɽ�;��q�3��r�3'i�ê}�
@I�r�q�L8ٽ\M=T:�=�E�Ϧ%�ݷ9�|��=p~�=_e��7!�=������r� =CJ�;�R�5��=j�M=��]=�]e�mF�=�� �<ؽ_�=H��=C`;p���ýy菼�_'���-��Q%<�s�dLh=�Z�=:�>�l������Y�>�X�=��@=�G����<��F<�"�=��w������<J�=����=T�=�r�_�=@���o�<UK-=��X=
���aD<�p>H�������\A<b�M=��^/H�	B���=���<W齽E�X�_9r��>z����<��;�W<�En>����PC������0=X���[�=\E߽w�&>�Ѥ�PTV>�%����S=m����?��\$��S��E)����7=�����������ڽ�|Լo�;l�w�p��;E����ڽ�i<�����=�ٽ��=\J���V�;����<7��n��ؠ(=�S�=�\=��C=�Cq��Ȭ������$�=H��n�������������ω=�h�<��=/�¼��>k=YxT= ����T����<���J�p<xC���e����^=�3�=/SȽ�.�X���� �=�$<VW��֗�����o�<R�==��'��ٿ=jE�9�3�:�����v4>Q=���=��[�^܁<�Jo=��a�܎I=�I�< ���Z�����d�����->Ɓ���Ѽ����w2�Ký���=~�=��#��h�����d�c=6ϰ�2mĽ�2_<��y���<���<e��R����L�=�½���=ߊ�=v�=�py�0D��CY���W>����
��;��Y��=dO�ᤝ���B=_m�����=���=�þ�ہ>��h<'l����< o�<�=�=�=J��%���-���>���<7�;<d��=�x;�0���lh�=�a/���=h1�;덌�F�׼�c!=��-��~o���=a��=8�d<68=@>	>��v=ښ༪�#=RQ+<mx�=P�<�琽�W�wB=vd����P��_r;�V�#�l>ٔ&>B6?���V=L�ƽIuϽ5�;��(�|Ά=�����h<�tL=�z�[�8�g��p���!<wٽġj�n}Z�G�C=B�;SL����<�=aN�����Mֽ�lμ�l�=id7=eB�=7X�=�=>�*�=���;=ڟC=S������=
�/��SW��J=�'��p����=%>�:��;2B���	��l�2�߽��=r�I>��=�5��K���[(�{nI��"�<4FT;�A>�=���=�˲��e!�
��;�=z�+=�|v=}ك��=�$��/�<�7׼򃪽�<�_�=YT=���.9>=�:=;D[g=��j<��<"���>
*b<��< Z>�F�����=yՄ=#��<騠=����=H��wD�S��@�=�=]��`�<��=��ʽ���;�<��>A�=��|Y��Lֆ=�����֨:C���o�<�R=��=��o����=2�=M�1���׽M��<'_=4z2��~=��*�����.�<O��;�!^�
��<�Jͽr%Z=�Q㽶;~��=��q��������>qM��������m�U<�a����<�A_��߆�d����)>>�'5��n=����)�;~��=c	�;�M����;��Ӽx\�=~�d�O;���cf<i�y�4���b�=9Fg���<S�4<���!�����=�x=F	>������<��=�ϽX:|��$V�/��lj�i(����&>;x=?[�=tt�=gM�=�� �J�Ѕ��(�I�=�{5=���<�ƻw�D��
��B����9�eS���P�'=�<��<��<�1ܰ=a��<ܱ��Z�ܻ
�f�w�=� �nǌ=O�$��=-��g�-�T�=se��HH>�F�='�-=���=~��=�ˑ���˼��#�u�=n����eIt��-<� =�:ٽ^2>=1�H���<�F=Xyl>��b=�S�:?߆=��;���;�x�=��=�ʏ=���=ݡ���H�;L֍�XV=&$��[�Ի`�`�ZD�=�(=���<�]���Խ%y28��=�O>$)J>�,'�]�=��|�=jZ��6�
>���^z�=ژ��䝽����(�q>��	�n��=~h<���<�8=��U<3��<vln=�Z�=�8׽�ef>j��3ش��.2��Ǌ���G=���>����=���<���<��=���@�>u6�=�>90�;�	�:��<�v=-�4��=�>�=�̄�q'*�/�J���Y�=ߎ��$;���e6��;���>�=ڙS=V/���l�=�Ɗ=X�2���w;����[u��y�=Fd�>Bz׽�`N�M��'�y=}�=t�=�D=Yq=�Lý��'��q���*>/��=�f >l{���>h�{�A>��(>���s={�\=�&>`g'>}d�>!�`���J>��>k܌���(<�>��;�r=��>�v����$M>��=1\=gĈ<���=���q =ԣ�=C�i=�&�=>�r��i(>1B�=�<)����<='!�c!<�U����=��ɹ���=���= �=fռ�����2��-��<�. �@A޽�vu<��޿;��]<�5
>O|�=��)����<c����y�<+�;^։=5��;�B=߳=JA�=�Pe�ɻ���y>�=��=�=����=i������N��wA��ԗ��v�Y���w�<w���\l��W���^j��7�=-����%�=�L��D�C� ;>"�>X<�n����X=3����<c��<a\q�Fd��>S@4��ν�Lq����=��7�d=·Z�qh=X�&>���� =�Z��9�êԽ?H�<��=,ĽY�<O)=��=;��S&f=�g�XH�<�c�<�����<�*�=������:��y뽣�<�1!<��D�!h<��4�2�����ڼ�M$=�2�<Ы��^��=��<%��=�a�=.���8���^;L�=� �<�l�=���=��p��=�W<�rM����<�ߣ=���=�=�*��kI�<�O#�����T�1�K=�i�F��i�>o��ڇ�=��=����D�o���8=��"��&�<8U�=\4��Y�>W�{d�;0�J��5��a�=�d,>��	��R���y~��zd��
^�=�M�=q"�H~ս[��=7�`��(y�kL-=��=ܔ|��q=<A]����=͓\=���;d�;@Q!>ɭ?="�&��7���o����9�{�<I�&��i��/�@��FE=f=�[�<��==r�=���R�z� >��<'X����>����=��]��J~���=�	�=l���q���r�<��
>\���QC�=
�;�½2��<ᩃ�g.�z3=�,w<|�s=�Z<��*��E��>J��=�c��=��ǽ��;�6罆��>����HH�M�=��+���=a�[=�=�%��z#���6�)8��=��>}[\=��=�R�;��>�*�ےg=���<�3���>׏��-���j<��e�����Ѥ<
����7�;s>I�7�W�t=�έ=�í��f<�v-�hF�<0G��$��=��L<\^�<�� =~�	�EЕ=�;�=�ט�Z�t=`��=���M�;���=�r�]2H����<��0���t�;���=�2r�j
�=��#>Wk>b�<K���9ݽ��N=�0��X�� ͽ�z	��誼=�&<����S��1�<�=Vl���=����X�`=���?2/��[�kk�<S����"��=#�%�טڼ��y� =Q���$���}�<7�Ҽ�>r��O�=�e�=����o�<�	��3��s����3=?vν0���('�=8���Kv8�/0a�
!�k]S�ˇ���2=u��x�	�Ho������}{�;%%=�ꔽ����P>�q���=���=[���۽.���f�=�_���^���~�T�Ǽ��=w%>����Cʐ=�(��W�\=x揼��=�>k�K��:�<�m->��=J\�=;i$>�l#�����՘�����"�w�R�d����<��C��E����;fb>�%>a,����/��<4X�=�S��=r/�;+rȼ��}�3W�/���Q�=V>Y�,�T8H���e<��*��v���=0�<׊�wZ=�@)�O�=�C<%�=��5= ��=��=����k=���(��<�%�<�z�����*��"g=.�>L@��)�=3�P=W����<x��=�"�+�=� o=56�<��=�ގ��V��ݽ��t�A�+>D47� �=-�ؽ=�>;ޚ��?M�=%�=7�}<����1�����=�	�<�/=D�>�m	�Y��=}}=�xJ=:��<е;�F<�'=��+�;�M�W�=�e���[��8I���=�b��3�4>�>r8S=�%>�����'>�r������ݤg=�p�����=&ǈ�p�S�%�<��\'S<�⤼ZI}=_4�VZ���~�9`3�=�g���=�=��=�t�o��}�����=�$̽�3ٽY��<y8��xʽ�4�З�lf�<���<cc<��� ='���=�S�=O����R�;*3�=�T;�:>J5üxJ�<#�л�}�<����h�8����[˃=~ͼs0F=��O�y~L��ݭ��bW=��:�%6?=�G@����=�l�;f˽<��;����=q��"�=q� �`�=��Z���=)=��=�
(<d��<�5νً�<�S�[˻=�-:���>�'e�������9< i��R=S��=���;Q�=\����=���;D�̼.	(>:�<(��Z{)=?�=��3=��=�D�?^�<WӼ�,=����o*=���=�w�=Vw<��=�<>��G��::=ֈY=�E�.ٽ���={#=vzV�м]�/���yϽ��s�^�<���"��<at=|D=7(�;��<��}:n���K��=��'>�o�!{׽�%�=}��=��@:��1>�|6=(�=8>����M<\=��=�ϳ�
�,����<�}�<������=���<i��<L�>Q䶽���</�3����=�Ľ�ᄼ�=�pŽ�0�j��%���><D�=�X>�2��=��Ƽ'�ѽ��14�<M&��#_���=�(��_^�\Q=�kY�V���:\�>`2.��eL=ꑦ=�~E�(������=7Ao�u�8=~OJ>��	<�,b�$�>7��<gu��1�="�>��=���=����%�7<�Ͻ_�i�k+<+0�=M�>�5>!���]@�=h��=�P��.?<G.>�d(>:<�d�=D����=۴�yLM��,ڽ��w=g4�=�`�=�Ȉ==y��#��=M@�;<�{="<��]>ߠ����;��==�z=��x�1A�=�p�d�(���=VY�-�>��0=�9�a�B��FR=�~g�f�=[{c=q׊<s�����_=�Rm<�����Y�&=��&�Z��<�J6=���;�M>�XD>øo=�J���*f�d}x��Ӽ�zŽ���=2���.�`�%�!�?���-;���<�C�����{;L�z�=z��=h�=cb3=�p���C��w��={��={���.b�A���%>�c���X����<��Xv�=[�!� ��=���9�==ő<ຉ�v�K<=鏺jj�=@og�:9q;R����=�H�<�6+��O�;��=x������=���>����2��&|=3��=CN��/���Ķ��M^�<8��;b�^=彭=��k=��=����0�l�A�ܽLY�"<��=̞�p�>ජ���=�	��00Ӽk~�<7R�=gۛ���=;�������j��y��=6� =yKv=�<h=k�3<ǿ;c�>7��ƃ»Ч��*�y�b.o�n�m�1;>�.u�X�ӻ��=��$=���>ְV�A>>L&$=�����<$��s�>���=!�:G�=�U�6t.>�U<4�����=��
>����0��
��:�O����;s6E� ��=ʓ�=�,�;:�p��F���B�<#����8>N�;�b�=%�
�k�=��3��=�&c� Z)=���I�O=W�@���6��0�=�8�7@>��_����!<�|��I��O6����#=& ����6<`�ȼ��d�q+=o�E<��x���r�:.!�h=��'���R�|
7�07�A���I
>٢y���C�X��>>�87=;�Cཆ݈=�񽑥9=;��=
ev���<Ң
�����1�S=(m��<Ӟ�<�f=�0#=3��Z>��:>����7��EFٽ���=�1
��GA<��r=)a|>a��=�,>s<:�K���O!>�J�=����q���a�=�E�iy��ee��
�޽�_�<:��	3<����=�3�=w(>k��%�Ju-�ޛ�3g�ꋿ�s��=�B
�Q�Q�Q���΀�=�P��2��[
=�A-<�(�X0� t����=.~f=Ae1=��=�k<���B��Eܕ�c�A=M٫�1:�=s~=9�3<���!$Ͻw3"���@z:�(q�O�<k����"=ծ2��@+=
�4��*�<=��=��9N=�����ϼk����}=�ݫ=�R���=i7=�tҽ�j@�~o%=s���	��<��ù���<�
����=g>=��H=K���ɠ�=�!��
�=}<�=X�c=���=Q��i�=���==�<U���1;�b=�谽�yM������9���Fa�9Й=R3�<N =�*���[U�wD^��=Gd�<�(�<��<���곽�m��e������.1=q��=h����`�ؽ��#<ΰ=�Y��
�8��=��a��K�<�\�.%�L�>=�ͨ=��Y�ٜ��BĽ�e�<�����D�<2=�����Iּt!3�,��=��+=��]
e�X����<b��"3�=�>F=N;��ԟ�=�;���ɡ=M
�I����!><��=�>�̲���;}S���V�=W]=�=XW,<�_����=��޽�=�0����=0���g���)����<� �<�Ȃ�������h�}C����k�4@>,�<͠�F��<���=l���*aI>Y��=�=b��=��:��t4���-<���=�+���V@=��=PΘ������%>#���*�ʼo��y�;ߒ'=!���"�E>����=�=���<{8=G>��ʜ2�[������=z�|=�#J=�'�<#��=�|=]#�ų<G�<��d�B���6��U����E���~�=���Y�u��ļ�]�=�k��{->i�*�ʹT= ��3H->��ؼB�\���>��=1���큽�0s<D��=V	���hd=�X�E�ɽ/�&=w�=��ܺj�> ����d0>��$���e���*>��ɰ=���ޡ�=*��=��*<�����㼖o�<'�>�\�=�M���0=���=uX=�>>fQ���"��ʀ�����;���=A߼FY�q���q�8��=c����c�=�9�{ �<]J=��=[��m~�����*�=|�<R�G������=��7=�;��|~_�����=�����	>�Q�=��O>�굼C>���� �ڇ���Ep�=���h�ğ��d�߽�-��$�=쵎� A�=[��=+����5��¨��������<Q��=�<���g�=���=~ p����<�w>6=�u�=M�=C�=t&��S�̽c�U�>��d��C�=�	 =��Լq���I2���!�����N*�"�Ƚ����)3��=������Eg�<G�������^��=;!>����kǒ��ù=�į��-��<�=�>H�ܼx�;w�>-���[�[�>i�=�
[�n�=�8���>���0�W�m�g��;Z$d�\����sN������+Z��b�����=�E=�|=T�`k�=��<�%�=�ˤ=��=#%<��=\�=T5>G��<�(>i�<M.���ȸ�%Hн�pX>�w�� �=��W=�OνK�|<:�<o+Ͻ �<�����C�"qk�Q^����=�<��Yk���1>���<��3=����ɽ=&><< |ܼmO�;mr���Y:���/�������= p=��:��H='�Ͻ�&Z>���<��n<:o��)�{(��*���d���$>Տ��}= (��`�����<��N�@a�%)`=d;�
ls>����t��V5=ԙ�i��n���v߾<���='j�=J謷�|�=1=�$Q��wi�z0>�	�=w�x=D��=L�����Q�j^">U$.�����|G��O4;�慾*�=��۽��ӽTlb=ݦ���oԻA"
��i�<��9�)��z���ʻ&գ;x�y�ν�;~�=V$=t�������?lg=�[ٽ�{�=��3>/,>Gmǽ<6�4N����wx;2��=��=I9�=���MC����<y$������H��W9w�
���=>۽��b?�<���e��#�;��F�R�ؽ�Dh�O�׽m�A���[���J=�dI�ѕn=�2�����#0��:�B����Z�=#�޻�bX�#��=ַż;�<�ڊ=���
�>x�>N=�L=�=�� �����\A�0�Q>^Y=��y�>p��T%�j%�=GW:>��Pl�`�����	5��)�=���=A�l<�,��B����>?� =ӽ�"$�����۽u{=������p��;$�=7u�=��������E�=}?������<�;7�Ὁp���=a��=g�T>;
=�ּ��=0�⼘ֈ=C����Ѫ�o0 =k��=�{��ݻн�(�g���50���w�K�i��|�V��|�=��=e+ü�;LgY��L=���y�~='c���=���&|= ɽ��伮�0����)D<͇�f�W�X,=Ѽ�>�J��f�O={�������ى����<o<�e���'��=����	��>d=ε�<N�'��-V��:=�=J�a�n��s����;��2=���=�w��t	��6l<|�>Li=d�ŋ�hK1����<T��<�ڷ;;o=�@=�&o=��=% �=5B���1@��g�/��;�W�=��K�n����h:3y�<n[����M� �0��;�=�/�<Q�0���;mL�����=��=׮=��<g�=*�Խ��> EU=��=��ڽ_��<Wo�=�"E=aԽތS<��
���,�V��<����.h�=N>�=tM-����& `=&<?a��=���Y<��E>'&ӽD�=Y_r���"��D�=�<N�K>�ID��?�<'���B&ӽ�GG<xt|��>k[<�4����=M���=>�y�=�	>��h(K=��c=�s�=Q����2>�E��sѻ���&�S=��Ž=I6���`�=�<m�D=m�.�j+S�Fԡ�?�ͼ�����ͻ|*=J <ԫL=;��=���twm=285�3���4��+>s��d�>Ƌ�=������=��;=�mg��\���t���,=2���*���p���`n'�rk��k��;g�Q>'*�1���[O=j��0P$��3=��->�ŗ��O���e<}E�<w=�=��I��+�=�3ʽ��6=�e����I�= ���D;.��=�'����<#�=���=�<�S��.>�C���P=���� =sM>�C�aǦ�h�=}6;ۊZ=�c�=�K���M��s=������+;I�
�ӕ�="���&��"�=�y�=9h"=Sֱ�F��;���=1�=;պ<��Ҽ|�>�x�c�޼P�<�μrC9�2�T�>
G��'�g�̶l:�8�=���k����
��A�}��W�=�M <��Ż��=9=ƽ�7=�HH=´?=me�=�����e�����x�P<઀=r���)<���<����<LR*����<5j@>�wཱ�=F�����>��̽�3G����=��=����=ܥ�=��^��R@��A'��d}<��Ǽ�L=�+۽��A��oR=��&=�F˽�ҙ�:�^���v�P�=��f�y1��=���>+�&a)=��U=3��/=�ټ��)=]}!�X��=�nG<�L��
騽�%~=��z�̢8>J���i�<�{>G}ؽ���@!��[�<]5U��"��O
��(�ɻ'�r�W��=�&�^�m=���J����=�qJ��V=?�~=�WA=�a�=��"�ƴ-=*�=C�0>�L��쥽�����=>��<�)A�s�#>�G�<ܺ�Z�D<�K'�\-��~�����)���@=�!>�(t=(�<@��^	w=�@�==U�A�i>�Q�J<�=fػ<� K>�cl=ԧ1=�-%��/k��:���>]n���T=<7Ƚ���=٘=�s��<�<��8�1<Ch��ˊ>HO�=���<+d��Ŏ�W�8��F�=h���N�r�=�˽�c<j�ǽ��ټ�ټ��ν�~����e���;=�@�������b�<)3x=��!��:�&��<�0�<I�=C�a<���;wuȽR}����<���>����=���x�=e�X>k>��y��<&f�=���;�b,�EƂ=�%,=����b��g�6=�����=8?�sV=jg>G����C=Z���-߽?���r��{L�=��M�9ﹽ�߼>�3�V�?r=�l��|�{�=h�=��=�������c>���=z�;Q0/��D��0vy�O����� ��n�
J��i,<^0�;T/]���NU���<e��<'���K,��{���=#��5�����<xX���>hY>�����<��<.1�ƨ�=q�ͽ�p�=~�뽐���=�J��d�<q?u���>X� ���X�>�p�=�v�=���;��%<�H�;ɂ>#�c�;=I<��.�:�-���Ƽ��=j9��0&����h;1�='N�=<@ڽ���k{�;#��(�=�j=D�=N�伇&����`=ް��\]-=N��9)�=܄��V��������¼֢����3=p��<WH�=~F�=h�=Eڎ��P	��퍽�'=�����ܪ���=dM=9�=�z�=��6���:= K4���2=`��=��.��>�ݷ=�#��H�=�|�;ֿD�}���ޕ��J~=Oƛ=����F�Z=~�W�����|�hн@�k=���="�=)�%>,�/����=���*��=�P�6LU<;��:G0���u�.f=�`	�ۼD���%����=R�=;�S=%�����E=�R�w�2�ё�<�#��L�=ձ�=5�<s�м��[��̀=,��<Xc8���<jjo;/�'��TB=���<��=��;�����˂=
q��)=c(�¡=��"��H*=�F<O��=K�>�-==�Ѫ�kԯ=�"���@���P�u�������}��D8���K=��Ҽ8�>��=>F�=D��=BU<�c��韲<��<U��=�B=���)R2�%`�<)�K��W=�S����۽ �r���H��ܻ��޽���sҠ�?�=A=35��}탽�K��p���߯�g�����/�=�%�l0==݈����=����;���=D��<Ռ���=���zν�=�۔;�^?��=�>����%= �<Ѣ�� �o�(�y9
���/G�=��-����=V����=�#�<�=��͇="P9�
=;&=�<2�*=(q�=�؊���<7e@�ŷ��n�=���<�i�wk�]��=ƪ=7��={�)���B�������+�ཱུWO����<ބ>�(>��ټ�����=j��=�[�zB�=�(�<��J;��_�V[�;��<�3��� �=/ v�T�=D=^T���W?=@��n9�=�sZ��-=V=�)�<���=�F������>��=��U=R1���0���kC�Ks#>����4���#�<[>��aм�q�񘄽�3��������ވӺ�L>!��;}�	�&�e�yW�ϫ/��Y=�`缌�ʽA����jE�C�W�ͽ?����!�;c�>a�!=eL���$�<q�����N�#����;�'$����=Ȼ>�"�<B��=�"�<���<f�=n��d,�)�;�B2>��	>�C�=t��':ȼ�ޭ<h�ϼ���<rV��
毼�X�;��ν���=�܁�?���d�`=1gE=����:ؽ��%=�7ҽ�)�hr>�?a;_ս�ܽ���=O�=N��<���R�b�4a�<�*��m�T=:<�^~=��ӽ��;��;v��m�#>��)����=�'㽔��='�;��۷��!�=�������=�	j�g��������k��U���l�<��=$X��]�����[)컑;C>G���=�W껔+=����+�Q�>DB�w���>���zZݽld@=���j[h�c��=ӂ��
a�=ʭ�u��=��1��k��U>���[������P�;�����.ν ��=�y�BM!>4�޽�r�<Is�6��<�ۺ���@�95=!��2�>ܓ=�)Խ�&}��4�=u	<�(���ڼ��=���=Y�$<��B�{�
����<ٝ)=�ۍ<���l�>-�?<�qh=���%�w�{ޭ=�������=��<L�I<�`$�F�>�|��<�@� �>̢����漄�:�z������� /�<��Ѽ
ĸ�������%.8��M�=��	�k�x�z
�<�,ļ�H���O�=����ؼ�}>�G"=�D=J?��q�=^����f�=�&k������5A�����w� Y���҄��쵽'PO;�~6=8??�R�X>Ǹ̻��f> {>�l�=�;e�Z:�<v��=\�����z۽�刽�<	����<�^�G�_<@�.�2�d���e��A~>8�4=�l=���=
�E;�+�=�2>��=Q+Ž�F4<><�R�={��<2��=	M�= �ϼZ2��	����=
�f=�SS=-x��UH��۽��E����ɋ=m���-O>���y�;�߂=���<C�+<J�k=a{�=�`ʽdž��>�L =��'����~�[��l�=��1�5�='	���F��`���KB�y��;CQ;Z����u=�ֽ:�׽N�2=���=	>��T��<^ۉ<X\�%�=�F`=8��=��=�Z=��<zXj�@�=I�
�,���\%�3ʋ<r��p�H�^ ���;>�"��bN<+����Ѽ=M p=��>`�F>$�B�-չ�<7��`?">�B�= W8>����ׇ�<5�#�B�=�.���K��~�=�n���~�;���=�l<}
g=�n�.|A<$ּ�g�ަɼ-�*>f׏=��'�~޿=D�=�F?=ٲ�����=@���5t=ɨ�=�#���>:z�l>?��ъ=�_P��=��r�=i�%�/�>���=N��+YQ�VN�=���(�8��M�=e?�<����2a=b�`<X�ν*�;�b�=��ź<8�u=����DD�=�i����<��>�A�=<:��������=��X<�`�i�B�[�=G=%�[�0#)<'�z"���X���C��]�:
����=v�=[g>(>���.=��x����=��E<���;,ܸ���1���*�,2��<�L�{�C=$�6> =7�ͼ��Q����:�ȕ�[�̹"ld=�Q���߾�ֹ<
�a=΋I���>�`꽌�ڼMN�H�V��=*Y>��f�=���H�=�-�=3;� ֽȱ�=Qj	�v�=�����~<�4��u�ƽ�&*;İ3���=�W"�Ý�=l ��l
�=�����3���{��C�=T'ӺS�����b���<{"$=�e��=�<��yu�<��=ڽ�HF=Z�X��=&bd�g�>=G�0�S�$< ��ر�=��ڽ��$=�
+=�C/�<����򣄼j�����ʼ�i�&��t�=�s��<'P�<qY̼�������o_����7=[�
=4��=���H�=����-uٽ�J�<��=��=5���v�=��G=،��S�sc�<�=l<�=���<#��:���=�V�=je�=~����$<�=�O=�l��P���%��;U�z��=_Z�p>�4��,�
>�_����H�>4=�iؽ�!�E}��M<��7���<8�:�׽�HB��5=�S���� ��u2�c(�=R\�<"D=���:��/�
<��X<TY�����I-=�<����l�=#gm�.у���(��Z<V�=VA�<t��>�9#�-ǽ�i?�=�5���L>��A={č<�M�=� �=�7�����jj'>��d���+��N<��#�a��=�����g8���q=ud���`=x�%2>�P�=іC�ⴧ��I>B(>�|�=��;��O�|� =�nl�ޛ���_꽬�>�E׼� ��<��!���=Z�m=�F��>��< 1 ����=�?�=k,�<��˽���< ]=\>���ӽ����`Et=B��=}F!�l�<�r�j)��w��
={�=O���Nr<�G�=�1)�kҽ��+�4M1�mD=蛇=�s�)��y,G>1���8)�`���=���5=6>�=t��	��<�`<2�f=Z�G=aTd=��i;k��=S�=���:�dͼ�F(��x=���=n��%`��z�p��=�a<����JcI�3)C>Kн����+�ڽ��]�%�e��C��=���= �=���=%��� >�=��մ<*�e��Λ=��=�Ե=U.r=T<>���<[���S%�s�����=��`��Ǽ<٫�q��=���=��#>�"�;8"�����Ar�p����=.Ư���A<�����Ͻ)�=�
=�x�F�<��>@(�=2�<2��=hs�o���؇=!�	>�;[�m=.Q��3:׼_��8�X=`���͈���ڽ).ɻS���)�	=�,8�El`>w�s��̜=�b�=4=������=���]R|<X7x=��<5����<�=��R��l	>�痽�պ7�������=I���-�X;Nԫ=�H�=7�F�?�&>�5ؽ�Ϟ<�FԽ�5�� �=zW#=�S�<�G��:�=�'+>9&����=oR�=�h�A�&;�渽ֆ���]�=3X>+憽w�;�q8=ie�=��2<��|��Hz=����.^�d�Z,=<�4��!��a�>5f`����;Nϐ��L5��S�<�@�<��ν5�=����j�=����p�<�Ͷ�3����g��BL�q�?=�o�=~�%HM=.�@����H�o�8G�f=<�U���j=V
��:I����V�=>�-�=����(������F=7l��Lwu�(I�=Ӹ}=�S�=��=ڏ�=���=;7>4[�<��T��^>��=C睽��F<�_�&% >�HN=4�ol<q�*��a=�୽K]켍���i�S��������=��x<��;=:pC=ǆ=��<�>K��//>r#�W|�=���=-�w�=���<#�ѓ׻��=mV������ٲ�ǾX=S��<��=���;����e���d=�41=��1��%ڽ;�K>��=�������-<���<˂����EҼ�XD=T�%���<H��=��=0%���*��?%�ۢ�������m�=N+��h}�:�S4�y�߼(OɼdYh=�6<��B=��@��A)�N{�=����-��LMq=��>��J�<��=~lR=�[>=)�Y�ve�="���l�<C=��5мo�K��u��"Q���<�<��,���ҽ���=l����=�<�pм
��=�v���B� >Nټ���=�A^>D��=6ힽΣ���+�����8�)��� �M�=i.a��c�tx�=�_	������WT
=� >���󧤽I�q=��&�f.�<�gۼ�q=�v�=$�=��I�i&=�oB=E)<ؓc=J�޽�������=�����(=Νݼ4h<��̽��;b�н��<�
ۼd;> >>T�;��������<;(���=�P���=�4�<�Gg�{��= ���d1=��E�[��=���_f�;�l�=���!�<]������>�[�a"=�{�=c���ZT��M
��Af<p��=�S�=���XG>�|>���A{=*�㻠��=k��l�=�x0=aԥ<��=�f�<=�5�AŽn�>Q0d<��>���<�ɽNS�=dZ���ŽNI=p�^����M >������=1L�(D��#�)�=��� Q�=�\���zE��}����=�1�ݪ>3\�<"�S=��}>�3�=!�-�=��������=������>�3�X$���<)m��eUd�2�S>��G<��>�Q���H������<�=�J�<�j=��Hf��<�s>�+>>X��oo�8);i�;����\�[Jg����=[ܽj��=KG=<ǅ�
 �<q�������c�=/?�<�k�=vo�<�5ϼ�t*=	����@�;[�==c?�ȐX��g��qӻ~xp�~�9>&@���Ƽ;���=I�=�E=��ֽ�<��R=�_E=���<yV@;�?E={ʘ=t��<�@O�=@�@0�;���=cm9>��=s�6���=���=׆��!ؽ�0�;&W�Okؽ*V�pt �A��=?��<�8�����O���\��k�Jb���Ğ����<~�(>EWݼ/aP�t����>�;��x���4=�Y���<�W�;g�>�L���L>߶�=�K�i�y<$�<q���`Η=�M��=F2=Ѥ��\�=�"��u�0��ͽ2"�=5���5=�'5�����>�Uܽ\D�ⴟ=��&��J��F�>.�=�!������K�< ��=26׽�B=�w���}>U���?k��nA=">��k<1n��r�;2��=�i���^9h���N�u<���<��<�5>wC�i߼<�@���{�[/�<0gq���Ľ
"(��^a�:�1�kA�;��3=�ǽ2�<<�½�ļ o���������<�v�P�P��׼��+�{�f�ͣ�;�����?������z�;�>>�P0>��p���� Ľ�.P=���=aI�*��5%�=D��=�a����>�k=4u�=G��=#�=p��=���<��p@z�l������zڼ�Y����=���.�8>{y3�o@ ������
�='��W1.<xT2>ҫ�=k!�>4���;��y���Z=���=r�"�ҁ�<@�y������9$�N���F�/>��=����ی�<�$<B�;G-t�k��=�TZ�ƅ�����2��f��lм���<W��u�ҽBhV<�����=���=0��=�=x!��fۨ�<�=���`*����(��<�<>G�o=�=�ؽ����B>�\x���;�(�<� [� �)��8�=���=؇�s�=�C�=�ͱ��4���;�/����T>��;ʓν<�=�f=Y�?��bƽ��?�Q����G=x�H��|�<��qַ=��'�8b>��<�!���M=���w��F��a��=�Ⱦ�3-��*<�n5=T�����<�C<��v_�0���l�!<�����3�H"=�i&<�������fS!��r��!�!���V�s��<?�u=��<�ae���4�)���]=ZP�=C�2>�Ƅ�L��vc	���+= ��:7�<.�=��!�p5�=k�\�=��q=	�j=�&G����<���;;�=MR��Β =P�z�dE=�k��[�<�h�=|n/;+��}�p<9�)=$C�<BY��c�T�j�҇��ƽ�Cz<_�#=���<$�=h=؀��$���<+�=����5cu=��>'(f9���=�!��l4=n4Լ<�ͽ�&��3P<J��;� ?��p<����`o��L�=Qχ=��J=Xw�<�b���.ܽg/ �Q���V��=�ߴ;�6��%>\]�ҏ��>��L<'E>��0=ϱ�<�J��� =��=�=�<���I�<鐦<��=�ϼC�$�̂�;���<M=�>==L_�w�G�O@��]�� ��=~�z���g=��<K����ʽs?>���=��-��)�=�i�=��ԽW��=�=$t�=V�=��ĽJ-�=�
=��A���H��I�v>h�����@lD�ЭU�����"Cy=뛊;�_u= e�����<�i�<_:�����=
N�=Dc��7�=��*>��'<�L=c�u=���>O=Ж�^����z=��>p����n:[=�S�=���<�>�<��8�;Jq>��=Y$$��|'>
e�= �<K*�=m	>��<�9�=�6,��H�=�j�=O� >�9ü�u����c=����A�>�q8=��=,jʽM�&�wm�=��G���ݼ��k������uG=i�˽�㌽�0�����fF�|c�=���B�=x����B<><�V>�!��9"��(�<���6��~"���]=5a4=,�t�������Q�%=�Ѧ��┼�� �Gj4��Z�/�g=��=Ű�=-w�=�lD����=E�S=E�$>ض�=�cQ>�&�<.I >N�e=�ה�o��m�R�µ�=/�8=�B��z���d:��]�6��=�!����H�J �=V���9��<"�������+3=����y������7�B�J��g��"=�)��Է<�9=��/>8
�<
��<0=�ýU�D��n���=��>�=_���`=h0��ʎ�<�}�����><�n�=i�Q�=�@>��N=o9��2׺=����C�=4�����=�=��鹪Ԅ=s�_���=[��%3��x��h��;s�=1�=��h=�`�<1���]�=�B=Χ�=d`9=ua��DؽkEO��h;-@��Ϛ=��=��>�)M=5>F'�^�=_ñ���><%4���'�3�G�=�,>�=|wS�w���^�=I��^Z#;x�t=���W��=%��=o�q��&C��"�<���V�=��*����&=�
>l�-�I�Xǃ=�V�(�VjX���&��98��R�=�IS=��|�'>~n0��p���Bl=8A=ٟ��)�V�K=ǫ��O����9���I=��Y=�N=p]�2�Y�䂤��ʰ=C���H$�O	C���=�[�=�_�JC�;A=j�~��>z?��^e�=��B�_&�����5��<c|>(F=��=A�L�^�D>�����x��n�{'#�"2�<�OR��7	���ӽ7�=*=z�9K��O�;��
�vw�w<O���N=q��=<~G��=-X�����=P;��-]ս�R�=O2߽VTr�*��D��=��=�w�;I�Ͻ۴X���E�o�G>�3D��5��
B=l�W���ս��<[��{*=+��=�݈>�D�:��"�ƽ���=1�E>􇡽?�=M�<4��=ɞv��};{sA�u��;��R�9��;]S��̭�>żi�>�ͼ�"���ז=����R��9�9�9����=��;�Z=�_�<�p=xA7= ٬<��=�Е<�u�=ڸe=��I=�=}�.=[G_<����A=q\н�սR����<��g�9���[�����������=��=�f�����-a%��Ӽ�~8>a��kV�1��d��;u��<ۆc��z?=K]
>7��<�l�=A�P�9�"���F:=iݽ0�I��y��EB�;~TνA3y��%�����
9>�D ��m�<'l��J�9>��H=���=�Y�ڞɽ���9l+���5;�1�_3�=y�ɽU٩��d���ɠ�p��<��ѹ��=�� N}�G>��@>V�<�x��TX��u8�L��<����#�ǚݼji<�5ؽ���=%���|I���*);�ߘ=�9���ӽ�����ֻ��<&
��Ӡ=j��=J�ņ��>F�9*�;_l{=C�3>��r1s��콉	��_M<��Ox�<��P�� [;�Z:�ZdĻ��=K��=T��=�޽x�)=У=PC��e��&���Mln�M �>� ��]����<�pa�q@=X����`�mO�]�{=r#8�8/��1>��=C|��2b=ïv�!��=�3I�f��@��=M]��"�{>�<;=n(����=P������?	;��<K���㽉c~�">�S=��;-c�=9x�<�խ=/�=�=s<�
ѽ ��=��:,��7��d�@�6���G=�!��۹�=�u/��W���= 
>�Ͻ��=N�>���=7�>R�=E��;k��fW�<�U4>^-���9��V"��+�Z�s�6 ��o�=9��<5S<MsD=�o��Ej=�A>���$��<��
;�o=q�q=ji��m��/�<�ڤ=�#>�?.��k�;O*>J3 =?='@1����= ��=y7�=�蟽�����xܼ ���|�;��>���=�&<<��Hn�<	�V=�&���n�������J�H�<��<��޼���A�=1��̍�������=kA_�Q�ͼ/S�H[��S!�=o��=��꼸�Խ1�B�K�>�m=/�+�+9
�i��=��ߗ?;�Y6>���\u�����+�������üP��<_E;I׼C����<�\o��ν1ä�C��=��P���ݽ/��<��$��@|<|m�:4�[=�N�=]�<�S=Y���g�T)�=��=�܅<%5�����=�9<Bk>/��p���z���v��Ș;u�;M�н�;>K�D����;龻�P>�Ww���֦�l�g>�kM��b�<��>c(2�0���5�K��:��f@ս1L<���;�<ȽK-�O2x��73�3�R�R^ս.j*���<ah=��݅�:-��=&��<�.�=�������I��=�=i]T=/F�J�=T���[!��0�"����=d�n�~m�<��=\D�<^
��D���Ǽ���
>9'�<�G<��⼝�#�T>��(=n���C=2�轖)�9�� r�'%}�D��<��>�|�<�y`���<C�=�A���'}<-��s����Ž���k���W���Y=�x���K���b>��>ǻX��	�;����ֽ���=)�j=�YO�ᫍ=`҆=�ɶ�`>�ϡ=�8>�7�#f\=�(2��U<Ȍ<i�<�X�=�@����<9��1��z��=�&�� v�˱w��G�=�И=4���8=�=�U3=���@�S<7*���؆=�1$�D�>=XS�<f*O=N56�7��=K�>U��=���=d���K/;'G�=�]-=:��=���=�H���7+=�$>Ȫ�=[�
�m�;>�3�	d;=HX�=�M�=2_=�2=�|�<��Y��dM����<]�<�;ۼ�\�<h&=+���ae���Ͻ];[=iE:=ᮩ=�s=����L>6��&�"��=خ���vG�0��{21��2>>�?뽶b��[��<������L���	>��3=��O���<�W�<���om�=�;����VA=w�����=�ƅ��^=>�*<�R���u>�<3=�RE�*���i�=�Й=�>5d�����ؽ�=b��;>�0� �G�7a��6��� d�=]}�<�$�����<ξ�=���=�!�����=6��=��=��ؼ���1A���ɗ=
)������0��-��U���!�ju�;�p���`�=�y�=�{=���/�=��<��;�C�=2YN� ((>r���Ž��-�3�X�� �}1N�K$+�{��<�w�=�\���b��n�%ν:�����z�=퀥=6�=��E<��=>�\�;�5޻i��=��<������򽮎0=�	>�;��ýr}ý	�z=�#Ľ��=z��w�<�$=��1>I��=�49��q�=r^ڽi����$ͼ�ǣ;�^�=��6�T�� ��C�Ǽ}�YxM=�b�=��8=�0���~��8;��@���"=�=���><E����?��@<-�<K�+=fd�Q�<p#:<)`q=�=�;�xu,��J���y�;ߪ��S��\�1��"�=uc>�.�=t����;�i9���r����=q��P<�����5=�	Ͻ��J>�-�<yV�;O&��4�=���=�.�)1�<(W�=��彆����J�[��=3����v�=�(�=;�=�ޑ������!>w.�T�S���0>he\���>�E��O>�!����5>�q�-�=ś>�����<����`�=�=D����ܴ<���<7 )=6��^<'��=F�%�A^>�^�=��?=�A�=/�<�� ����=qL�G��<���JR��q}`=��j=~U*=��>����i+��"=��T=�>��D����_&=�9!>���=LV>ry�=B�y=9�	��'ѽ˲�����'>��S�6�� ل=�F=�@�=��;$½��2=�$y;ߪ_=�� 5=��;j���@���=g/=�����������=$-�=�⬼�1�<!ʽ޺���q=i4��+R=�-�=4"9=[>��6=׀=�W�=��=i3t=���Li��j7o�nC`���<v��p�=OW��O0�Aܼ���=���=��ռ��(=�B��,�=ˣ�<���<p�=��,��=�6�< Q��T*w=��;%@�=�/6� x;N_�0��=�ۼV�������;��h�D�=�C�b=P��<���=&�˳��'Z=��>+��=��;�[@���:~7��kɫ=��=�ݣ=��,�$P9>{���d�`�=�*>����`<1�>��@>��*;>ᮼj��>Y5�;�-=���<�Yؽ#=�
�=�a,�Eݽ=p����ʼ�:�<G[��x�>��
����'=�/f< ���>�=�=;�=6֜���<B�OLq���<޼D�M�0�=����=�3��z�L�ڻ�~ >&�'�m�=�vԽPU���*ǽ�񎼺_=��<P��� ��=I���!���uzS���=���6q��pѽ��1>��=�%����O<\�Q䃽�`C��y�<$��8Z��r�k�|[H�r�o���˽v���ǳ=�T
�΢�=��?����04=�����Y�#Z��Ƣ������7���=ԤӽYLC�᪂���\<�&<c,��SB�r�>f�{���޻�+V��V�-��=KԽ�#�\�� 76=�#+=<^r<�5�>�>��\=�Y���<=�[h=m���0[d�D�S;��=5�ɽ|��P>���m�=�u�<���=u�t=��;��=��=�������姽�*ؼ�Uo=�ߧ����=��ܼ=;�����I������=�C>0�w�[�x��e
>;��=~�=�El=��J=��0==Ǯ�y>�ȽԭA���ӽ5Z�=�H<Ӕ:���#�e�X>d��$�ýO7����w����#=D�9�V^><W���=���$���z��ؠ=e��m>тR<f=~8X��|��6���δ�<���/����$�A�= "<��=���9"P=�D���:�<�7��q�<s�o;�&�=�k��ԼL���J��6�4�_?ͽl��=� >EL�<9���k=�ڼ3>ڐ�<�:�=�B�=AA��̽`����z=r����ɼ|E�O��;3�W;O�ͽ���������=��!=a���7I�<��<Us�=zG�=e ����Q>�ʜ��ܽn =8:��}e�1��<	(S�B��J:��>��O_A��F=F[�=�Y�= ��Q`���z�=�A�=�'>�}��7^;��i>5��=������L<D!=�yC=�T�=N�=IG@��$�=}��=44�����<�:��@�>Y*>=�A�<=���������=�ϼ��X=��
>�e�����/�s<�������ص��ZмǶ�=�Ž����+����,�f����+=g8��e3��{w�;���D���Y��çf=T�`>�T�� ���f}�x;�<5O/�*`��0���<s�A=�<��
�-W/�^ӽ��<�������x=��#��������'>�2�x�)�J￼/�6�E���?=H�aY��	G�=�k�$���8=E㌼#W�=Q�d=Q��=�����"�p��[>�A���R=f���|�����)�\T;�C'����=)Eϼ�`@�T!>�!ǽ�s�=�+�=Ɂ�Q��=��=�l�ZO���&���黲RZ>�U��$���<���Нټ���=L��=P">7^�=@d�=�hg=�e=���Q��=fdC��)=�ҽx�d#B��K=�^�=��<�ˤ�!��=�oֽ��M<��v=5�=�k�=6Zs��޵=3s,���hF<p`�=f��=*�9>ew\=�xO���c���=W4->4�>{^F>T-���T�;�޽F^=δS=��2�炼=`o��.=F6ʼT]�o�B��)l=5&���;��/�aZ�=6떼Y���ּ��R=T��=��h=V*l=
��<*�=��=��C=/Q��&1����r��=.ɶ<�Fk<?�.>��n�A���,|> ���
�=3�=���=��d��=T�	��:� �<���=���n�6=e�L�!�������S�=[<Au�=X>�έ�_�:c�ټB�0�I��}Z�$H={ƻ;�E��ղ�U��+�=�l��~�<tD�9l,�=r ]<�,�zS�=Ձ�=u����!ûU�����B=r�M=�x�V���~��yCs=�)>��=dF'<�k�=��=2o=�P�=?Yf�Wqr=itڽ�ꑽgIg=�ǚ���>#��<!"�� ���顽�����=�Ӿ=�*ٽ7bӼ�{�<���=��9>V�Ӽ6ϙ�*Jd�Q�l=&(�<>ӽ7g>�%='V>��q�=1�����=�(�=N������=fQ���`=d���6!��
&��R��;dP�/�r���=?�����=���<IY¼���� �=�󿼹s�G��=�^���;&=�+_=�C/>���H�O��p��2W��N"��N��3=\G�=N���9g=�X�����kRS�碀�}?�}�=4!.=���9f����R;�fz�<��=�p=T��=����ø��j�=a���t�=��C=B��=��.������ü�򆼄��=諅=��<Ґμ��	�* �J�w=�;=򀴽X�=��<�.�Rq���e�=M)V�[����W���:w=��<���<�҂=�=����<�?L�uF�=����`>���H
���㮶=`i�=ѿ�=u~���>���������R�B�z�h?��/��=y�=P7�=�/�=� ���i����<�� <��
����逜<Gh?�O�Q��ʙ<��I�'�v����fV��/�<"Z���~]>[��=04!��u�=�p=8���^�<TS�w���<�-x���g<��-��9�<K�ӼL��=��[=$����z�=)<�A�7��z=q��<������ɽU�νi�Vp�8v���{Շ��憽@{x�$�<k6�=I�ӽ!Z�=���1�<�Q��[B��d:���6���0=��U���;U����Ƌ=H�^���K�?R��z�.=T{v=O�,�"Tn�9k�O>nh�<yT�<����-m�s��<;�=�v�=�[�<�}-=�=a�ӻ!O�����x�.<%��L�;NL��rc<%7���19I
>��d�,�$��+`<��=�v<yE[��j��}4>T�����{,=�����=�����ý!.����<���=9(�����~�"�L���MҽIDS=5<�=>e^��@���g���r&=`��=��>�S�=+�ڽ`F���h>�x�[������*�ͼ�ٽɽ{>R�ý*CI=��w�}_� ǀ<�#;�s��<|�i�7��=������<�����`=��Y=�(�����>��Σ2>+s=D��;���;@Va=�H"�/|����(>nz���D�;�.==܀�q����A�,��Zk@<@>��Q���>�~��������6��=�#�����&<���;mآ=X��;{p�JW�=��^6�=�o~�΁>T����=+qs��o�����D �5ݔ�1y��J��-f���ڽk���"�=�=�b�l�ػg.ݽ�|E<���bd�~�<�=>��<˥�9J����=��u�#�����L=�s7>?�ϻS�	|�=Gu~<�,�=��<Î�=i�b���=���ˈ��H�=`��`��=&!���%
>!���ｘ��=�"�=�C����=B�V�T����G=��<�|=L����|�������=0pj=�d���=����Y��K$>k���e=�re�R��<Jp�<Dr��_ڽ:�O��Q�D�<��x;���Ģ���{>�R��#���F�F�
�����X��t>�I#�/��<r
L>�i�S@�=ȭ={�+���=�����h;§۽��=]D �Y��� B�=ʷ�ҷ	=X���Ӽ땶<㕍��|:>:x;=�x.�f���]�=Vp+=u�<���ML��Ņ���>� �=�2>�H��Ҡ�<]�*=Ęӻ+=I�WV�<v���޲"����=�v�<�ὸ����� �*=W0����Cǡ�s�0<�{�;?!�<4rC<��=;{Ҽ��a���X�AL��eL�=
���!�-=[��;z�.��>H?>&n��<>�rн�߉��3%���V���T����7�;^��3����%�<����1~=t'�<.�=�g�=f���r�=��p�n�(�˽����z��:��3���E��;��M��U���ǽ�<w F=F0<��8>�V���*�=�S��ܼ0�*=����W于rܻ�
.���=v��=!{=��}=l����%#>�%�OI{:%	�Lk�<9s ==�󽕂&<y�>�X>]�1=U�=^A�=��e7<7�S�{Y=��5��C߽4q��_�n�����e=�]L=O�Ͻ���=5ڜ=�b�=o9Ľ��{�x�l����=���<���=ߒ�=�.�����=�"=�)@�]�d�j��F2R�!W�ʐ�[��ĉ���&=ꜩ;;@Z=��?>6�1�f���ۗ��4�������]>�O��ܽ��˼7��=�Lo�P����ڱ=͸�=��ܼRȥ�l �����?�R��<��
�H��nN$�c��=�ǽ�`="�������$�,��s|<�����ݱ��g��������= �,;�+�r�/>Y� >�>�a=��'<I�<dl
>�%>f����S���|�<o¼���=y=�q=`8q=p8���a�u��1�>�����=#}�==��:[�p���(�
z+=s��:��*=8���+ު�E8&>��������=�$q��X=�̠���v����R>�w=,���h(��,�A1<-(��8�ʼ�!ؼ.!׽�@=�.�fX�Uۺ�|=B�J<��Ľ�Z�{y=�j������Ə��}'��MH>o�:<�e�<P �<���+�������=!��mֵ=b=e�/=o��#ȥ�cZ<2��p����$�)� �<�����d=<S�뵽��>�i�������>ث�<n���R=�?ʽX8<*]�m����a��Zҽ�׺rOb�J*�;؞�=�ZP:S�	�I󼽸�|=�ҽ�=J��p�F��� �=߄�<�*=QIe=��=M��<˾��ߘ*=��{=�4��3�&<V=��_V�4��R���!�J=��p�(�	G�=��0=�_;�>�2�;7q������fĺoV=�5�=ku=�d���S=�����oً<"3�O��f-�=3�%>����_�k=u ��L1=�l =���=r��[+�<��<�｣�$<�4���ά��=�䜼��^<�>B�����[ڼ��޽F9���U?�_�<�j��KȽ^��=+��=��=v� >u���7e����m=�j=憯����=LY�=�S��E9�:*��<6[���1�= P�<(!��	����~<����E��=�Ƚ��;u[W>�9�=<)�2 J>�5�<�7>b8�5k��i-�<���<�����T�a"�<q��<�F9�k@��n��=x��AO�<W�����s;Y<��^<�G��
�i=�~�����bJ�We>�)�<<��F<1O��i�{=9T>|����H�F��=ǴL�����O[�x�=��>c�>��׽7��;��=g� ��Y"=��8<��!>�b�;�v��Li>��=�\I=n����+=��=P��=T S>*��=�H>4W�=Ϊ�=+��=����2�+���u=�Y�<:s�<&�>�y��ע��^�Խ%|��>��=W܏<^�*=�n <Vb>N=n׼;rM{>���<F+>Xm�<�d��ȴ�=QP�=`��\;!>�[G�s%>�{��_����>Lme��ҥ��ǽ�}��l�=}7轗��=6�Ƚ��ҽ&�7_��J	=ᚊ���l=�w=���=�B��p��]¦=^}�<�@=�f+��~b=ͽ��)- =u�=���2�=�a�z�]=����=��R=9�>�	=%��Ƴ=�dg=኿=�)n��@����+=/,�r憽��<��>�N�H��=(|b=��ټ�9����=&���-�=��ӽ�*��,=K}=/��L�ؽk�p��q���.>��=!���z)<y�*>��ƽ��ҽK>+=i���]M=����H�=��=Xb=�G=d�=�ka�<�Vu�7��<��R��g�=_�=qx#���=��<��=����.d>�3�=�{�<�y�=��=f�M���Q�}J>|`ý�}������0'=�����0=�G��2&(:��<���̎=�vĻ�+>�QA�X�1�~o����z��VJ�u�4=L%j�r���꣺��N�� ��A�=+@=��½Ý��(X<RJͻ�=ޗ�=��|=��:�?q�����^k\���%�j�!���;�N�qu��_�� so<=V��8�k=�y�<9�R�b����N�=�����y�$G���D=o_]�U&�R��<��<�%=�w#>3ߑ=�[~��>}��97�%�a�<���$*0=�F���`���G�.�ݽX���>!*.=]@�w�����bt�+��_�<���=��i<��ϼn,I���;�
�=�ݳ��[���L=��=,N�=ݽ�#���a`��#���f+_=�X	>�f=�� =p}�=N�I��sE����=ގ��R2�<��<
��=�ة�/C���:��+��b,>YP��.�;�v|<�T���"=��=��Y�+ֽ{��;��=�<�7�=*�{=~�L���½�8>�ν��ݽMv���cM��XE�5�/�1o�<a�dX�<��=�,���q�ؽ>��=�)=S�<P+����=��(=p�?���>��E�"�6�u���νlQ�=��<+׆�g4ƽ�6�=D�>=�=}���K�=	׊���@��i=�yC����==�=��ǽ��O����=�j���a=���=Q�\=a�r<�K4=kB�a�=���:��y���=��̽�-Ƚb�2�u=Pa= �����O�<3�b�9�U=��?;̄X�����(˽׎Y��ũ=}��1��$%P=H�4�͎=���3�<�q�=�� >�\�<V��=�J��;Z��c7�2 D��>��B=��>y�<R�>�&�xgk�z��=(��;����b����i=�u=��M�����q�O�8�˽�&5����=$1�������S�W�R(�;=��X�d��=E��H\q���<H䈽����x
8=Z�K=_bQ����=@	�6��<���;/3p<mS#;�����=�f��Z� � �1\l=t<	=V:X�);=��= �=�o��cᠽD�Ӽ�3�;-�r����2���z�����F��<0ڽ��ҽ�|<z7�<�K^���;��<�M�= <>E7����>>b7!��+(�\�ü,���n�鼗�;>��l=O�^�=ľ=���=�	>�P�=*����~$>:1>NKͽ��H=� �����=�"%��n��Z>x�<���<�|ӽ�Ż� �=j{=�=ֵb<h��r�M�������:-�>�_���Ag>y/>g��;�;�����<nH�ы;-V(�U"*���>��'�>�Jd���<;�M=�9�=P{0<���L����=���$�n�E��=�M ��rK����;an��4>�G��4S=���<$��=[�<�o��dw޽��=��>���ټľ*�[F>}ǃ=�Q"=М�n�ʽ���9!�>�Тx�REq=�붽[��7+>��=�Z>��/�a����սr�=��ݽ��=��콥��=vҼ9�>�cýkh>v�=�����fJ���*>�x�;��=�.>��i>c�>^)E���=��k<q �p�v�Ř
>g]���+=?�Y��8��+<�su=eȽ�9�=���=���<`���ǘ�Yn*�)R�= �"�~�<ф���7置lڼF���4=j��<j���1E�;P�=Ũ���2>d��2��z��ȥ��浽A�7�_%��9�$�=�=+3�HL��A@(�\\u=v��<��=/:���������Ӝ<k��=��=>�y=V�ۼ-�d=��Ѽ;��=��:�&=[+D����kٽ�v<��D={==�.��R����n=F;O=4�h<��7���b=�7=^r�<�=h/�=��U�����=��Y��w�QO=�=G�>@2���Ȼ��q��w];��;�߼��ѽ:�=P/ܼ��>_�
>�mx�bj��'�z�,�F��c�<Ns����#�鈛<�^�=gbP=��oKм2���-��v�A�%c�k�伅\�<��s����=���<�u+>���B�l�5>gت�r)>Q"�<�<Tf+=�0��P,?��n��Km=��<=��̽��=v;=Fr��Tt=C�^=�<q=��N=��4<���<�f{��W�q�J=ֹ<�Z��f�8�<YF�<�瑽
����1Ļ|Y�=^�:;�cf��^�=ϲ�kΓ=%�s�͡I��*>{��=�<�3���:?5�<h��=�9�<ƹ�=|υ�7�=���<�$1<:�P>��S�j��=��<������=uG���=�n$>"@<�M仧�w�1X���T>�u-=�җ�0Y���_�����q+=�e�|�̽U��=ͪJ�b�=���ߺ<��<�A�>J����=-��<�U��~I<���侸��w�d���ZZ�Vfj=F��<^���N��X��),&�d�,>�����z<w\8>"��[k= �f����\�&�ԟཤJ#��8>�e�>
��	�=����i��f�=182>$R򽇼�=A!<>~�>����P=��	�T[�=�h%�
�t=�?='<�=���=
<x�(=�O�=*�H=�
���c%>c�>����;v=�K�{��@�>ڕ���b�~.����=a]�<����S=��="r�=�ن���ȼ��=��<�X���u<vw=0e���O_����=�~��(+�;6�=c�u=����X6��0м>�Q���o��yS��z���u0�fA�=�#�=�Pǽ<�!�=z�=�M�%8��'=u�;X����&`��|�=RSv;\#���==�pk=�{<A=���=�:	�oԼT��H�iN����=�J������_��н=0�=3 �=e�c��}=���<��$�%�E=�ib��5O<�x˼�|=�4½��ڽ�8�=�q�=,#=3L=�4�=�[>1����J>��>�<a��<���=/5�=&w���[m�����J2����=��彩��:��	��� �$�����
I[����X�g�7=�W6�3 =�ᑽ��4����Df=NH�=�d= /������{��'e�=60�<>��~1�=�X�<��>>5:=<0<'kG=�f;�yD��ݶ;�{�=PGS��ϻ��[C=�c�<o����Ǹ}JE>�O���$M=w�K=���ο<鴭=oX����9��3
X<�� �"�=���<˽C*�=�����O=��#���m���C<�f=Ƅ἗�>j�u=^�8d����[��<"�a��>ס�=��=� 3<8��<�qѽ�6=���d��I?=�>��M=x�=�~���=���;}E�=�w=�ѽ�iI����=F�=\K�J�>=��g<�xm=/8��=�>��=�&��Ɣ�<�G>��ʽh�泮�y~P�E�ٻi�s�M�=ߞн�]�=���=�m�=� A>�j?<�����>��<���=��5��ʡ����r�	>N���,Y�<��>\.�x��<[�>̚J>q �=�� <~�>�:û�����"L����׼��<�*�=b�=��w;j	�L%��߽��$<��=ùк�%p���p=xW=m�=���=��$=�&�=�o���^9���=��w��ٽ��R<)��=���=�8��)	�+�߻Q�(�uX�;��k�<�)�<�J)��f�<搯�_@>�K==���<)�=d<5�yy ��B��]��%�C=�!��Y�+�;g=|K�>�Rg����<;#}=��V;�sO=����Đ��S�%=0ͯ��}=g<�<B77<)��<�L=�_�~o�\px�v��;5N�U��=�.����*>��=)��b(���w����<���۶�#�R�9��<IK�<�x���= r�<�&�=J���5o�����=�4̺���=�|z�Ѥn�����~8T����W�1�[ ��
=>>�ߎ={�����<�a*>#�W�}�d=K�|��t>�t���7���2=z�{����<���=���;2	e���	�n�����R���<���kY
<�������(>V@��9�C�A"���!�:PkW�&C�=S =~Y���<	9�=Q#=QD�x_E:�Ё=�=.��+A��%u�<B�=+T���U=,k��)���u�<hy�=�Fx��������=)½�7�<K�=�]��B�=�=���=�s3=Ħ�=�>x=2�=,9���Hk<~��=�j�<*=�rǽ
ݠ���:�� C����Ka ��/�=�=�<��=�$��f$�=���<��1=N\�=>�=�h�=Z��0�I�P����E�b@�F?�=�<u��x'>'W����>I�Y�t��;�'���Rk=EuY=���q� ��[=��|=V5��(S�=�;u��<>%����۔=�U��ƽ:U�; ��=k�ۻ�	��Ɠ4��(=�%�<w��<o��=[��<M�s����ݽq�K<4�����'���:l�)<�
S��㬽+�"=|��ꁼdw����ܣ�;��#=q>�i�aS�<!Z��v�J����=��>�=���_O>/o.>�^<�>4=���=B��ZvO���8=2�(<�"=�ִ<.�ټ�1�=l����=�����������=p� (�<,F=�p�=t��,U�<�]0��x
�"���璽2��=�F��	��+�c���=b�h�j;Dw��ظ=v
R=���=����_=���=.XR>��>���l�^<�q�<r�ӽ���<��=ɸx���x=�Z���=��<�g�;�t��)>�Dн�u�����j �! �04�=���=Мj=_8�=g�->8�2��¯��L7�ދQ�	��Tȹ�'�u=��u�:�cü��;亁=q=]:o�����ӗ���=�N>\m�=�}&=	����o��S=���;u���M��V���G��=�}e=�1�����|½�;X��5P<���=Q������=���=���ɽyN���� ;NE�<?{=3�i=�=�OU=M�ܼj���'㟽��n=�9�=i)�<Y��=�ǭ�z� >P4d<5�
��-=��=X�1=�^	>�S;�����y&=׾>-���V�<�2T=����<D)�D��6}	��h+�KC����%H!=�q��].;=y]=h\�=��>����;�^��;{�(<��<�=����>?��=�R����<����9AK<�Rl=&ã��K<-�1���=eR<�Q!6�P���r�=�r�
g\=�c>7Y&=O�&�n��= ,�;����x$>��V=a(�<��<�����\@>�(�<k����,Q=mE����7>,ax�`,Q���=��l=e�
�#���4>�<�gH=�p=��Ѽ���<��<���=�R.=<�'���½�����>2�����&>~�c�S����&^==��=#-���N$� Z�<�ż��H=�5����u/>n)>�W��|�ԽDo=��;FtA=fFY���>R��=��>S.�<������<�+ཛྷG�=+y�=^燼�_��h1��h�=��*��p|�K������<[�T�wnv���=�A>sė���=�_�=�:��״=mRS=�;B�`�$>3u!=�>��
�cO�;$r�k���ޣ=�"=��0��(2=�}�����SO=A����H�)QK<���+*=㼰��<��<�$�L���)���$=-ڼu O=�I)<�D=6���<��<>'>���U4�<�����R��=�q=ֽ>��j;�u�<tRN=�8=t�.��aX=���=���;�N�ٶ���M>��=M%���<���=,���<����:�^��<�S���<Mߥ�]
;E�����>1�=�0Y��~�=!j��i���=V�=�ڻ�+>޽�� ��j=$���Ѵ>��R=���+(q����=�V���F={Ņ��a>�	��3<�>޻�4��/kk;�_��L=��=T�K�61<(�j<��ߕ;�����N�4�l�s�� ��= v�<�!�= �=�~��/?=݇���=�l=`�$������9���6=�\�<*����#(={���+���<@�=*����<p>�]�=JH�zb��P�ｳ��=G7�;�X8>�4G�{ػgpn����=b�->�� ��~q�T=#�b�,�a=P�G�	�1��C�=�&h<h˛���Ѽ��u����pN���	�=Q#2�@��<ܡ˼�=Րx�;�Z�]�<��M�<f��<<�>�\���Z</A-��Y��w4�>c���v�Ph%��rP<�����	��v�=!�>1W�=��=zZ�<�V�=.��=��=<xp<��q�Ă�=�3���n�?�>D�=�ܽ��H��T�=�<7~˽;>~�꽥[�=w)�pf�<͉=�OC���|=�k��~>���u�ݺ<�#=�ǻz��ꌴ=��~��Q=�/r�����-(���D>�;j�9=��=�^(>����$��H������'�I=���=5��=&L#=��=������=onE��<�<_n�=��>b��<I\�����d�2�;}>�00=�M�=7/=�R;=V�{><��W>!���)�Fw�=�ܼMֽ8��)����Ľ��=�4�<����j~<�x=���<N�ý��'>��Q=��+= %�C�'=I�׽c��=+��;c%ܼ�ʶ=�5z���=�I���>��霼c��=�0(��;=��F=E�=���)ö<�'-�#�/=Mk��i�����a=��J��A"�Y�O��J����<�ᨼ�I�MS
<�=8滽,�=��Ź>kP�=����W�<\�#>F��<Y�߻n�<h&�=�ۖ=7M=W�.>LP�=4�O��z��f�����;T���{� X$=�(�f�>�Ca����W��M=�iI��6p���3>L��<�]�����X|�<-�=o~U=��k����nB;�-=�B˼,O�=�f�=��=�BC��u�=m���������<��)����v>���5H�V�ȽҠ"�[i">�'�i�����V=�/^���ͽ��&=�ɽ�Ŕ�Z�;�f>�ɾ=�n&��������8h<����� �=c� ��_��r�k;*j����=��<���/�0=�_'��O"��v}=A���鼼k��Hש�׌�=��8=�����X�=1煽����\=eR}=S�i�&��=k��=i���zP������VԼ���<8���}�q=��<�>�P���>���=c4(=�X���}=Yp>��=�4��M�<r�w>r�Ԭ(���ȼ^��<VWA�&���7����H�=�J�������.{=��A>�;�=�"|=DVJ��{=b%�=�0��O��=�� ���U�q����L��H�J=�@��=�ѽW���D�%�旞=�G>�2�=�h��!�=�G�����=��?�%��O��<&=�R�=u��u��=4��l)�����)�"��<�\���,>#E�;�k��=���L�
���=.P�=�2�=)=Y��'O~;wq�k�j�n�萓��?�>�>��ý��X�{�>�~l=�>g�g�Xw;�����X=�X�=���<g�ؽHt�;�Q�<�M�=��'>#>��<y� �y�=��6=�z~=Yf��6��S#>!�O=O'�4=��q�=�0F� ,2�\�=�p׽õ���1�)WG��2�=/���W�ż�X��=���<il�������l�<���0-	��) ��y�<��,=���X��=%m�=��=�Z<�,>��m=�Z���u�=ޮ==rp=}���#""�_"=�4=��<E�=F�<V��&��Tu<�����D��HD��C�"��R{P=�᳽�Z߼'���.�=_� ��$����;3��=���<�����G=>"��kc=޼�=r2=MJ�t��ꏡ=����L��:�{o<���<��<��=��)��E�=�V�=��>!qW=R �=dfi�_Gx=5��=|ۻ��M�������)�=/<ݽ!,׽�%=[�:�;�<C�$��/9��SK=�V@=9���݋=�_>+$<���N>����(i5=5۱�� �w�𼻫Ͻ�W�Ie)=��=Q8 �C���Ƚ9d�<Au��ͫe=�l�=��>=C�O=;� =wb�=�H�F�=p$��1���<4Ǵ�w�������xB=�0��h~=U9�c�g�a��=�C�<0f>C�G=X�v��v�<T�=�u��7<>�k���;{^*�Wz�X��=32���=��>���͎�)�D�>����<.���Q�;Г��u��(2u=�Ь�M�Ž���:���;����|��=h����E=H6�=q��=��N�EiX�Yeмܨe����=��D<ͨ7�H�>^-̽�=�:�=Y�=&Y=�>��:d��|b��h��=Ѵ�<�_V�s<B�l�<�|��X���1�=�7�-|��Py=��a���&=<C��wP�<��=�
�~���u���&�=&�g=:���<n�f1�=
� =V ����=%�=��=�T��e��&�<B��=�e�=]n:=e>㇎��T�����:1��=(���š:=�B]��,�y��C;�==�i<|��y�<�И�;�۽w��i&��C#>S����=|�y=q�;m���?��;B?�Rʎ�f�>կl=�6��<$ �;�ӽ;=r�<����e���=�ӹ<";5;�O��=0`�<5�<t�@=��1=VtC=�=�jo��t�=�s�����a� ����:6I�<,�O���<���=W�^���=e=pw�<�����0�=��.��R<`vf�B�*�[Լ��1��O|����=s�=�=�>k���ݼ��>�*��=�D�F[ʽ+��=�g�:��><�����Z�<>��,�ýka;S*t=;��ٟ���]�=S��<��'=5�j=�&�̞<�д<����}N��L��<>/���N���,=�=0��;e�>>i��<��<.�<j[�:�j=�~x��@6�ѹ��0=i;=�����=̽<=4\8��9�=�r5����������"=zp��3��:`9���~���=j�>�'�d��=S�[��Z�=[�q1��g��d&��f�;�ʹ=Q��Z5(�g$<E�e=�p�;s�g�Yz8��n
�S�2��Ϣ=��D>�r�<�
̻��1�z#>�%���:&=k���B�E�c=�	��ɾ�ï?�pa��&��=�.�=E|��i >�뎼��%=9F�<B��<�o�Z2�=�8%�!9�=�y�_z\����=ӽ���=]�I=p"k=�W&<~�D9[���,k=�	=��y=��>׎>����S���Z-�!�:�+��� .<��P<�6U��^�=�""=�J��6zn�]Z.=�,�=9,<������g���l�J����k�ȅ�=?��<�y��B���F��\F�g���^&���䩼dL�&�ѽ�>g^v=�����3��|>���=�\�=�N�'<�=��ʽ� >�S>�˃��ض<:��=˨�"��U���<,�y=� ���>i���T="��=$A�=%�:��O=��=e���uB�Y�>�t9�}꯽��e��}==]M�=I"B=�#�𗋼��D=8��_	>�sL��-��d�=:>�>	�ҷ�=�C=�
z=���>=���2�=���=�A��ɼ,=<'�=�'n����=:av���ר��C�늮=G͟�R�:N%%���+>(V���7������ >IF3��������0��=��>owX���ҽi.=vY��xڼ �m=����O�9=��>@��=_��;�#�<�	���(�HU<��>=3�*=<��p�+?߼#�N�lyX����<|=��&��b��Sl�*#>��=V�=w�ȼV�;Kf��$^=H3޼.�=N�=�ł;��<��j;
P3�x+��֛=��=�������<M��;�W�=c8�="N=!mt��P�a��=��>�D�g����Q�r�=�B'=z���Rj�=��I>"_���Y<�^=���37�����T��=��E�`�	=�w�+R�=C�����=)>z=�4�����. ;���<���;V�I�,F�=���=����2�=��#>�=^T�=�s����C�kT�=
�0��`�</���Oֽ;����ץ����>������ֿ�$eW;���;|,"<MC�;|�]=)Yo=XD߽�3�<:����=�G9>���=�<=cݹ����9v9��l]�5M��`�8�����P����~��㎽b����/
9O4ü���%�/��=��<���=�i�=�*׽�x�=w٘<9��=�e2�;�*��>R�+=���=� �=W/�;
���	���xu=�	��[�X��]X=C��9[�e=j����=�<��~=l10=�o@=��=\����ټ�3?=����;"���=�e���(s�������=9R:<���<�d�=�v(<�_s���W?���=t�>��|��P��P+>�Ȥ�e�h>��ܻ�m���,'<oWǽ�#��je�l�м�~�=�A!��=t#g�/���.Տ�@X�<R�!>���<^��tӣ= /�<�F���Z����=b�=F&�t�:��_Ƽ�n=�K%=$�ֽ8�=�<�=kռ##׽��#=����j�N���;vI\��Tu=Z�=� <ڟ�=l��=J#�=�%����/==��<)���Xm�<�c=�0c>����o��������r=�\(=�̼���<S	L=���<q�j=@�ٽ��	>����[^�<A�Ǽm�Gd�����=��#��9><��=���E�=�NE��������(V<�,��ƴ���(Q=�X�p�W=��鼲�<X\�	�1=h3u�Z�<*��iM>{��;l�=l3�ںr�u�$�3�,�=����-��=�<�=<ϓ���z<��=	=}�z�A)¼g���eR�ʒ)��==��ǥl<�ؚ�qU:�v�z�@���W��<�'�=e�\;ꗠ��ב����;d'м��ѽ�1�<�;����}�!:U�$U�=D�u�V��= Y�=��¼�0i<����i�;i�>=�=�K�=���<���[��=)��=|�7�8�/\������<>����={��=7���q}�y6��G�z=����q`;{�P��*���ֳ����W߯<c�g=����Y��È=$6X<�Cz�C#��������<��7=�h0>��D=s[:���>�7��0���2����F=�lu��+b���6�ڪ��8)<O0�=e�{�֭D=��W�5�=���<�d�=5��=�L�=2�=�O�'��=��@=�x�< =�	n=�~�=(|8��b�;/oR>4~W�f�O�3ߒ���I���<�J���3 �X9���=�5����<_�=�f��F��ɼf����F�=�'�qͽ9��<y�V=cY;A��=����%��	�+=f����!<=V%;�i6��W)��l���{H�Ɔ=zo�<`��=.gJ>��=P�<�T�<��ǻ�=<	{-�O��=�m�D)�=��q����=��w��o�<� �<�)��?���>=�-1Լ3Y���8�=�����ߡ�ý�k&>����*�=�Ь�G�>�hX�d%���L>�*���
�=�:���R�=�B�j�<;�={�=�<٢��*�<�=�������l�R=�)�;.	v<Ƴ:I�=� 潋̽t>�~��$˽���񻼽�E�h�[;�� >���?㖻�Z���z=3�_=�jp�|q'�{�;�@=Ŕ��91�<ʹ���X�<���GU=O"
���v�T�T�2�3#>�O;�K�=z�ޖ���t=�F�=!8���YT��̼ޭν�4��t�,��\��ls1���>0e�<ϓy=tE�<�#ɽ� n=����#ZK:��x��輌`+=岗� �?����M����l�������3 ��.>�M���h#=^.<���;/#.>�(�=������H�󄽌�);2���d�=V{=���=&P�|��=�
��LP������<gg�3P>�"����5����T��!'g>��J>̘���
=Yj��Ŧ�1�u�Z�=��.>f����x>��=�M;��"<�
>w�r=�M�^����!��"��]��9ha����<���ɳ6�Dp0��lb����1��䶞<e>{4<kj_��+�=uI����=�]�;�;���0y=�7N<C`�=9� ���|<l;�=�'$�hoo��;=�藽��<��=��=��<P������h/>Zw�<���=�G�=��̽��<4 =�y=�N�;�Ž���B�$<�5��t�qѓ�ں����=Ń�<-u>_fx���]�w>�=�=�1>�?���������<�oS<�_>73���ܢ=VE���ļ}]�] ���ջ�����<�G>�>�=�P>��D��Yʼ�M��H	_=��ɼ{A��/#>�6�=��=�o軚� �A�T>_�����ؽ�	�=������C<�=�3[=B�w<Yp���;��^=q~>�^���E=����=X�=���<^�3���w=UY���@��"�>ʽ6��=-�L� ��<H�5<G�C�9���R��	p�&�|�#c�=2�=��=$��Z�;=d�=���Ҧ��':���=",;���=�Y�JϽ�%>>e����경,.�<wH�;~[ļ�|<�"�>0��g��*
�=�$W��r�<���=<�~��=N��= ���(�P�����'~=NO��]A=��;=�p=g?7=�V=٨ɽ�ؽՀ�=b%ü)�H=�)��AFǼ�)�*�<����b=K��� ��=C��:ֶ�=nz_=o�����O��=?�F+�={�k�����1��<�=ێ����<Uz�<M9=5.�F]�=��<R��_��k�Wא��-2�/E¼=��=l��=�_>�����F=��Q��-�@��<:�$>Y�=� ���U�<�x2=Y%��H��<��3=�g�;��=RL����=6E�����IP��a���^�=�k��#����>ɼ/�n=]����<nq=�l�;�^��ˢ����<~��=7�	����=O�Z�0��=��C��/H<e�߽�\��C�u���=�W�<��;;xY�=����'�X<��
eh=)�_��7��t <Lj�<dW�=_��A{���c=���hS�=�m��G�=d�J=�b�=�r�3K�u����?����=;��=$�>\��<?�����<8�>�6�<n/ͻK\}��*=��<2��<��=��;�>�ا<��(<��=���=I�W��x�<.H�� >��	�z>��W�=k�k=��޼����k`<������3�fa����`���ؼ���`Qk�Q=9�˽?�۹�L���=�ܫ=��(�ﺋ9,&�����x���&�;�X�=@�������>s��<$^����=�/>���Q�པEs;ͩ`=��e> R.�AJŽ�B�=Ȳ�;o�D��Խѩ�a\!���v��:�!��=�S#��=�1�=.����<f岼^>p�r=��i=r!�=D�z���<�Z�b�A�Y��=3G =4䰽GoJ=�>'��>�<u ����;[�x=���=�=U7�=����~c������~b�B�T�",�����=�X:<:	�;��O����=��;�=Bܽr�Ժ;����#Z�!7h<uH��vG�=�1�<is���GX�1ů={]2�\���f�=�8�=��a=�~�=�����>j��={�=Ĳ_<�V»��>	z7=�����������q� �|���~=���<p����=��j��kм�'�=y`,����=�)(��(�<(�<٥�=ņ3���𻟧�=�7ļ"�f�:��<"W��#���=�Z*���<��C<���e=g��=���=��/��VƼ�'
=��=Qxi=P��o/�z�=���<_�=�!��둽�@��>��:�o�< ��===���=����S	��O?:���;ѼS�V��νT���X(;=�
��h��/�0�%��=z�� �`q<#�-��+E=�^7=YV(>�O���0��&K���ɽ�&=�r��d�<�'u��=�㼁1��Ѳ!�S�����̽(��<�;A��ì��ڽ�'>@L9;�2���;:z=��
�)���9�=��P��=��"�ƫ=a�^�!�=���<�՟��=�>��<�=�g<�˽f�����JN��^���5��KW���!z����<"�3��c<$|�=������<A?���� >�l��Z(>����M#��r+=�=:)ѽ�T����)=ݻ�A�z��H���U$=���t�=/B>��B� �<�����p�����9�:=[��=ԕ$<��?��?�=�ڪ=< �Xx�[:>>M!��ܻ*��M��p�<��ѽ
�?�_ ����Q�L��J&>.>�6x�=����2�j�:���%�#-|��4>��%>�b�2< >io=p?���>VNY=C����l��<�!;���<`�����:=s�?�.[�=��:��x=���<u	�=���=`�<�g	=#��<K�=<�b=��\�����q=��=�Vr�3�<��)�x��<��n���=�?������W�=�^��O�]<�1ݽS�;���<��M�]�%>�^�C�8=<y=�C�ͭ<%�=sg4�C?�={ң<�ܞ���O��Խt��u韽v�=C�>���<�]�=@L6�vU~�ˇF�]|��o�=�iD��(�!Y��鰋<������=��j���S=ٟ����>�}��0��6]�R���A�<��5�@��=b9���1T=�sO=*�1��
�=:�=�;�f箼�Ƕ��i�=�����!=r%I�q�?�j�;>04��ɹ;�r=��<���3���<��'��%=莗��a!=�փ<9��|�e��*�DuU���=|,�
��~=�#�O<�½q�=�¿=DǗ�',���t<�'���p<�ѻ�N�G��`*���=����xս�B���e��E�1>�'>ڴ!>��g�	k�=R���`=-��<�=>�97�;��9��SW<��=��=Ԛ��Os�>��ؽ݅���b>3<u?��f��=�a�=Jc��=�� ����=�{�<V��<��>o�@�����<l�Q�c�6;���<��c�;&�=��l=TP�a1�=�¼"T=+��=��Z=3[�<��h=��=����OL�=R%����H��AἙ��<��=^�h���ؽ`&��L��hY�y��w�&>F���$�=��]=���R�=4�9&>��>���<�hӼk�C��:��B�<ܸ����%�H>��	���=��=b�*=�Mo=o�
=H�2�o*�=��
>�.���ͽbŽ.��=��=B�����<��< ��<�$������=��=�#��CY��� ��Q���+|=��2=k�����=�#)>%^����=��;>�un��T�<?��B��>���>�D���6D=��y��2=��=9����j��E=��G�><p:Ә�=ڽ�8<�	�m	Խ���6I��8ь� B>T=ʽ�ȍ�{��� �@=�F��$gn�D�Z�hZR<���Ex�t����<=��M=�~���n=��潬����1>���;��r=��Լ�xW�Ğ�=ՍN���t� �=��=��=ad��T�=cc�����/�=E�8��.����1LH��=�r(=�͑<���<XK���<��<C>�=m�����>8�ջb�S�8M���9P;�?_=��=My3=/9�<C*��c�<3�=Y�):kQɼ���=��ͽ�:Ҕ5;7�>�㈽�~� W&��٪<!s����<[Ӫ=�5)���<�=��5��:���į<iR=��<��ޗ<�k�<��<ק5=0<<�MF=ȝ��p�84��:0½T|=�\"���=���<��h=z}���;�@�'�����8�4�=-�=G�=�]E���
=X��e������Z2��T=-��.l<|g���B=�`�<��.=L��<���jn�F$½ј齒�y=b�Z=�+���E�=��3�Lq�=*\)>1�`�҄콢˙�#�f���üg-���. ����<G�n=�N�9�ā�`c�<R�;���<Sۥ�)�(�P����ɽ���=͒���N=��,>[v�=���S��=0�1=���<+�;�9[=g��<ܙ��(�=�#G=o^:���9>����l��Ǩ=z�����?=��(1>�H�V�<=�T.<@I��%FF�@�V��������T>k��<X/)>!��;�����н�ک=��&�l�����޽N��M��0=!(�=��=��;�'�s������<�f<�65>�]=�C=�����M>�.�ր��P��OI>G5�=7�=�,�껻���+0ɽ�nO>O]�*o��g�=��T�<�Nl�0�=2R����='����<>��>�3�=��ڼ�
O>Xe�����ۙ���*=�n���<��;�3=�a'=><�<$@�Rum=�	�����:\��	Z=�	-���̼��>5�=Ε�<t����<=؋�=��q>]s�<y�<�f�=Q2�<�0?���*��� �u�+='=>��9����=��N�O�=ʍ����=��=�����мU��CF2����<*�����;���=�(=q����=����yӽ?}<�:J=���<�=��>��=�F�����WȠ��y�=OɁ��n�=��#���e����<\*;Q&)��2����<�L]>I�g��dT=&��=iԟ<�+��h���.=|�*>�+Ӻ%h߻��=�$=�E����z=f���`Ľxƕ<ZJ�=ؽ����g;(<�W��Mw
�&�=�1�Ťj���򼐁F=zH�=�W<�=�̽���=-��=)Þ��5żT�s�Kک�	�'�|
�%Y�ۑ�l~�=��>��=�H=�!�p͞��N2=�\�]~��fx+����=��_=�*<���N��=�<֖�w(�=3u�<�O�<�Ҿ=��=B��Xs仺B�<�_�������F=U�@������>��m0�=Wҽ,����#f<LD����<9�p�E��==�ƽ��_;���=�>�-��=��g��=x���ܽm��\�=��<��y��<�H=��S;A���O��d�ǽ)𓼫Fp>�x�;*�|�\`�<�=� ���_����3=��N�=��<砼Za�=���~�<��ϽZ�
�e�<���=M(��� >Ȝ��m���M�=T�\<!��$P
>�D�=8|��*��9|o�*?�:�>�`�=�ƀ=2i����==�I=�`=')�+�R���u>|@��`���>J	�<¨�=��_=�4���l�=�e�<]�M=Q½��=dօ>����J�=־==�0>�|��C$�b>$=�a�oђ<<#�����=��(�����?>g\�o&�지=ю<�Ȝ=oQ=}Ft;�߽�F���"�;D-����`�=ӽ��=��߼󣎽�x�=yL<]��Q�(�U;
=�;>	�sˁ�2S�=Të=k{�"���6�=*.�<�>��=���=Y������^Y��.B=�=ڽ�VZ��Ͱ=�V:��D�;�Ѝ��v=W�bf�6W%��:���=���=�٭����S?�<�Lq���=�d]=�֜;�+�<���<���=�'��5+<��=Le@>J�I:���}���n�=�$>�`K�=�W����=�Ì=7���0Dp;�'�=��<�U�=������<䑼
���W����=�5����p�7V��S�!��g�v=����w�����
=Eν�O�'�`'��k�;���=B�E>8�b=����T���Ž)g�~u =�Ƒ=����~=��*�� G=^W��Q*<���=��*<���<�/|��1=s��=ݎ��b� =���=�X<�O=�!B��<i=E�=1�y�IIf��"�sh�=�~==��l=m��=:	1;bң�E�	>H�=�#��. ��ٝ�W ������K�=� }���=���X;>ۜ.=^�n=�G��a	>��<4�����9������6+=m�>y==e劽
�<�.Q>�>ټ��-�� ���<��n��4O�����g���^��=�����*�=��3�H��=
��O$ĻU�K<�,�=O/Z=<e�+?f=���!��:�J=����6^y=�=�=���=�R�t߾���1��hz�Ž��3/=�;<*e�=�z={�=�ׯ�LU�=׶�=V=�->�`����$��Qrd����<6�*>%ڪ�-�<9��)t��o]��2��=N�>�B��_��>����b=�9=��=gEa=n��=oT�=�j>�d7�qC>A�<�p�=Oʭ����@f�I��=�y =)�I���/����=�=��s=�:�=Ҳ��נ�=��=�*2�� >fDɽ��=�=�'�Ƞ��a�:���-	>�3�=1vݽ.�\�K�=.�̽J�=$=�Z�{=une<V��=4+ ���>��q�l�+�L~=���=N�Ƽ���=v�<(9���=�{>�=�.o����2�=��Q=tҶ=h����^��`�<2�ʽ�r���1g�������A�3>���=�e=u>�y�<4���f*���)���<<���=0}<�H&���<�r�<]֕���=��ݼ�ő=��m=���/�f�5�!�f���<�C>�=�ᙽ^��=z�R@=6�q=�b��s>��T��^�%tԽ@�׽�1>���������x�=[Q���=@>̼�<�(�=r%ۼ��=� �k5���x=�>Q���{�������1��\'=������=Pg>�m�<	|�<e��f�=�u=�4�=b
���a=޴��D���>̏��G�A��<7j�=���n>��^=?�����-��d<���=Cz�<b�S��mݽ��<s�=4/��l	=�yX����ܠ�����=��h;��= �<j�ؽ7 u��<��*���>��L��i�<�hZ=���c�ob�4��;������� ���V����:#L=m�|=�qY�/a�����!>���;-c�U�<_1㽍J�<7���l����<F��B�=�?�=3�=M��=�X-�_�<�I˨=M�����>X��;B�<�/�<_�	=�̰�%_ν�1�=U���w�=��л o����=Sj�;�z�<u6����n�z=
p=I/6=&�I�z�<"�d����=kQ���==餽�s=G����� >�K���x<���=�J>>�=@Qٻ��%���e>Y>5:�,�=�*��8$;>�q��^��
��^�;�-=��<��d>=S�=��K>�@�=ŦM�۝W;�r�:.�;�=��ֹ*=. R=$�,=ӝ����=�o�=O��P�;�.e�=���=_�ټ4�C>�Y�����iA6<Z�=��zt�;6�v=i���g�=��P��J`=��x��Ŝ=Ĩ���:��H�aъ=�y?<MȎ�ʡ�<��d�;��=eg��&~���л5�꽝 S=�G��%:��J�<���=5
�<�L=A�=�<EЖ=Pm ����=b��m8��w�<�7=����μ�O=��=��=������ջ ����<
9��4����:�Ž^���Z�=T�=/�Ƽ�Tz=e����U?<��)= ��<���ޥ`���<i��nI)��Z=�l$��@7��"<����U�X=�[���N�)Hm=�=�=�>�<>�=��=30�<'M=�u�;E>�xJ=��<-ƃ=�0��Q�<�������4��<p�9�܈�<�)�=��p�Q�<�N^��<��`�=X�|9h`<�+>��q��=����J�Ը���;���=�>=�fݽ�u�=|
K=�QX�iw�=�&�U�= t�c�ݽA�缰���Ӌ�=��:�+����Y;<J0���2a���|���I���@��&�=,�!>���4�=ռ17���8=�v�;f�"=��8�b_�=Ƀn���x��J���ٱ;���=�Ee<�����=q�=^���]/�<`#ԺR�>��0>,j��d�)�3.�=Iȑ�L9E�p�ҽ҈>;�����uO��.��<�DJ���[=�%ҽy��=+=<pW���-=�k�.�k��=+�b<�j��y=1��,_Ѽ����ӹ8�=���8P��&<12�<�sL�zԒ=�����L�7���9,�<	-��+�<�3�\��<[�=h�n�׺��I�Լ!%��D���a����=�b��L��:t���o>���1ս=�$=lCR=�{�)/�<���=�>�=6�W=z\d�|	�<�;Hsc>�g�}��=q�����u��x=3���Љ	�Z2�;�B�����=I��_J�<�2[>E[>�ὢ��={5>��U=���G����H-������>ܽ�9d�� ���=@>�3G�e�?��%=�̪�Y�1>�1�����=��=-8ֽ5�o��5B�ab:��������<OH���=��X�(�|U
=w��������Z=p;YR�=Ll��I<��>�.��u">��o����8�<>��L=��<���=�y��p�뽼���?�=���<.z+>��=�����6�=�ps=�V=�:V�ö!=��%=�I�=vQ�=x<��Pf��ƈ=q�սT�g�R �ZX>e����>]�۴��	�ѼW"G�B���&�=����5�=�vƽ>d<�hw�KG��j�J�>V�<pf �0�<Z��=�{}����=Z3�����Ƚ���<��^<�F��<�Y=��>�}˃=h��YЅ=o�3<���;Yi�=�=���SL�ò�<>��o�<�m�=���R����#���nV=��X�])C���<A�<bI������$oS=LC�<��ǽ���Q����R�=�4s��!=�F�<�7��v>��[��`q��HP�� �o��=[(g�	W=�9��P�<�l��î��a=���<S�=UF�=U-=�ܹ���t��㸽�yi9��=.Gj���F=�d��:;#�(�ڠb�6ø�Fh���ʼy�;�aq�B#�������$=D"==��u�f�Ͻ���>���;�K���~;>s�<p[\��|R=�U��>ں�˿�A�u�}���E[�M�=8��V��;��=���=Ti�<����9G>��<Zƞ�a�ּv������<�T�l������=��켎kݽ1���)[(�m��;������=��<��V��ݼ;lN��R�	� �X���p<k����_�`i�=r�=}�p>"��� �d=�=�νw~�=�$=n�=�=d=!�=�� ��i���=&�=ӳ<<c\�<VP=�8��;ؗ�WRZ���z�7���=�$j�+�F���UR���S��<k���8�/�^���cD�=��=���<�V��*=(�Z�Ś=�|��Y��=@
���� ;��:=?�\>�G�����H��\���;<}�=Yl=�CR=yDZ=�>n=�阻���=3;�<	S�=�ܢ;ǜ������1=�0=J>�.E>�=c<N�<	s	�'�w=� 9� T�B��Q7�<1_�
ˀ�<R�=0½�l]�,������F,=ګ�ZoG�?=���Z��ګ����F�t;��Q�Fd�.kӻ��J��MF<PS�=]�*=~).��{�=.�����=�M�=]��K�<<��<�:k��̪=t����[���ѽ����|��>����J޽]}�;8�|=���<�B7>Q	>�4�VO��8�t��d��/�~���L>̡�<�����?=�l��=��;꧙�?E~�ii�%#��������6��m�=���<v��=`�'=���A��<���.�=1��<s�:����ӽH�=,z�<���=	��=;8H���F�w��=�]�<<�>e�e���o���=y��=bI�b�ƽ4�)�d�=3g���X�1 w�FC�:^ �=<d{��`�<�6�=;�=N���zmC=��=���6��=�N\�/�Ľ��'>�:#;Rd>�zI�/�ڽ�a�=�V5=���螼;s�=�ұ�^�;�>u�=�j=�s��U">��=�={7�=`�!=�=D��=���:�=���S`</���ʼX:=ӎ�=��ɼ$V>A�����=Vi�=LQ �!�=��=]�ѼQϷ��&A��Y�n	��?=�=�u�=���pώ��E�=X;���I=�s��^#>�dE�PK�I��=�mB>���=.�R��"�=�4��l����n�=O���Q��jJ�=CB������qT�D�%��a>���1�>ո�=m��=�=�ʗ=�
�i�>��f�)�=F��_�܇�<MM=K㒽j�ٻ��<�G�=ay�;=k}��_\>�?�w�;�fN> ��<ڦ;�����C!<+��>kr��!�=�6���;��=e�:���=�Qڽ�B������v)��1��/m����<�����'����;
A�<�c��	��=����;e�����*>Ө�=���=x'>g�y;�/��o�=�0=Yn6��d&>�*�=}w���
<�U$��6M���>�7;E�f=4TB�{ʎ=a	|�AؼY����Wk�;�L�=���=��;�� �v$��>= ��:���=�|>�����=!��|)�;�O;=v>����:�=
*��o��r7��e�'>i�	>K �=�q�	����u��������=������Ӽ�2���$=�����;���=q��<�����U=�g��y�������J�=�`g<񢍽^���H���� =؅�=��׽_=Q�G=��g��D\���/>�����~B���z�\�	7g]���{=v�=%N����_=7
��m�=Hl;����<��{<�E�=ϭ���0>�%����=�3�<(׉�X!��+����}�|=:o�����=N��<��b=@@V�ِռR�(�#ҍ=���<O^E<�7�1<ս�zM�}c<P�=Sa=_C4=Ͷ.��*��=�=4)a��^�=a�=i��=�3�=^���>��<f޽���;�﫽g��+Ɉ���=��ƽ��{<��'���;�2~�W�%�x/�;¬�=��ɼ.η�E��<���=�[=+�������1�n=�	�<B��Z��<���<=�����=V ��=��<Q��;=���'����@��	�����\=��⽰�>b�<g�s= g�;Ͻ�����=���=���	w�<�۸;�|z�G�=)>|�#����?�b��b����\5����$<{�]�e�0��t�yJ�=�<��=�oe=���w�R��,��=^�<�􉼢Q���^<Un>��=�+��Y�>9�=_��<0�����=�<4��Cڼ��=�b ��)>��=M��l����&� 	�=��=�����}d��fʽ��'�V=E��(<Y@=Zɒ��{[��^=�t�=� �1yB=U<��p��Y`u=]I�f��=)܅<]����	����<�����ϼ=��8�4�8'�<=!�<[`}�����M�.�����=��M;k{&:�
F=�R�"�=h��:�<�C��9�S��<mS<m����k�I(=�.�=��<X�o��^<��# >Q��g�C�o�=�Պ=q�۽fg>y�H��>9<�st=OW=65��Q��<�q��|#��_=.��<@��;i�=�U����4<nB�e��;U��=0��7h=T?�5�='!�<}<='�a��� ����<�1<>�<�=��<���=�G��]-<XWp����ɖ\��<���=�ռ�$½���=�f�T`)�O+�*�>���!w>Y��=y�&=�7�e�:=�k�=n�>.�Z���˽q��=Kn>�u�'�Xe�=��u"=������
���[��7*���h=�E�=Qg�<C��-h�;��>>[�=�� >j�\��2=�56>� ;���= G;ru<˼�<���=�,���;m G��=l<[����д=�  >��=p��莽���=�=S@�=+J=�����������U�C�Ǯ���$=�
=�a= �=�K�� ��=\U&��#���@��wR�ri�<�|=A��=x�C<��|=�m>ġ�=���ܢ=0a<1�<g�j%�9�B<�ʳ=�-=㵬=�vZ��:���]*>��3%=}���D����:^=��@=�`b����:��?=h>��=�k��唽2�T=�%�=�Ez=cx=��e��=���; ���gqI>���J =^�>okE�)
�R��Ǉ�H|1��j�h���2=Зa�"��<�=��ͽV�����<Q�O;�w'>@@�<j�E=�Pݽs��<� =���=�#�e�=��p�"�>�'<��x��	��qҺ�C�e��#p��> �U���J���B>���=oU>��Ľ���<a�=�
��:�<6=O=*�B;�=<C����F<��!��=|Z��|���*=�%���.=����0��=�=2�<-����%���臽��l=��5�?6x��o�6N#<�P�<�,�<s�yª��m�<�i]>ю���G�����8f-�Q�-�q)ʽ�7��c��{tM=w�˻X�����<p���rᄽ�D���Ɔ=�e >�lY��r��=�g�Pl�<r>|��F4�=���=ҕ�⏃���L�����*�=�놼���uU=:�>�z�y�c=R�4=�G��	�� ��<���;�>(�=�=�|�<�1ۼ�Y�=���<�i��X"K����=k؍�θ�=��U��w/=�>7��<+QZ���)����=qÒ=���{~�n��=;I�=^��]�@<.;�=;�ܽ��5=sF��ߙ<�O�;���'�
=(b������e�=f�=��w��4=�8U=�]罽u=Ь,�QT!�l�=!�_��k<��<Y�
�<�4�<:��!8�=$V=���=j�#=��1=Fd��j.>�:<�q2��Q�<���<��ѽZ�=�h4<8�|��dλ��=�s1� ��<�B��\lf>�~h���=!&�=5����#=�I�{��E��<��a=
s=ȼ&<G@O���m���������e�= F�=	���ѽ���=ߡ&���>=�h�����<o��<��=�Zw��c'=�>����;�	���M;)'(=A��?���ܽ�i�=��P��pE��q�=�y����f��������h=\���;�
��A)��ҷ=\��=Z�0�h�Q<&�~�����*�<��_���j=Ga=,x=�R����=�Y=Ʀ<��>-��=��Y�@q�=��=
�S=�<%�C�h�g��=DR=zd��><ws>A�ż���;���ч=_��=[Ӕ��@n�$㌽��H>��<羽6R=�L�;��\< 못퟽�u�=��t��;�����<�Hr�諽�R��o>��>��w�i΁���d>��_�S��TA=nI��"��=�ս][�<�1�=c��n�>�A�<#�&���>�<&l�;�#�]��4����=A���*7�= �>�Ҽ;Օ�i`>��<����,�Z��<:�O=9�=���%��=Bས���j����}������=F҇�7μ�eL<�Zx���=8�=>����� >��b��0�"�>��=�\���m�=�`$=t�P=R��<Oս��zn>R|7�o,=�}�,�=���=�Le=ލ<f���j!˼$s���*j=�J>O�=tjݼ�f�=�I<>��;��=��<��T=ڃ=�z`�<g94�s$��P�<KѽM�׽M�x;�G�u4 �s	�;�� =��=ed�<��W=0㽹BF<�������<���נ=�~-��=��}Ž��z�=�A�:�����S<�`�=aF>*��=E�S��m�<�~R����;�|=�/N��~�=w�����q�/�5$�o]<pt���f=�ܑ��WB�7�
>�̛�z����s�����u�;[��f5=��'��>���c>���=���=��4���+>u1�;�D=�c�<ȾH��O��8�:����c��$e����=a���%b=݃I>(�="�%��=�p�:�ܷ=�ע�y��=�<���KO{=�@W=���=�y������S<��Y=�85���=��བྷt=���< �
��䒽�3����<De�G�r<�z��޼�ђ�{�U<L��<.)4=�Q���=��ڽ^x���#�=З�=��=R��<��~����=d8�=��νb�>�`���_D��Խ.r=��=4{�=G��=������=T�K�6p�@�`C���p'=XM��%$�`��Me=���<��a>'׹=]w>dͼY��� ���C*�=��=-�����>F�.���9�/�s>��=���y�����<��'�Ǻ���<i>��˽e�>�2�S=��ļ><�k�OT)=�ה<�V�=]�=/�����>�=X�h>����>���>%G�=��=�F�<�W&>Jن=��Ӓ8;Ky��4=�$�=�d�>��Z=�$B=�et�9*�=�+ �oOͽ��ƽ�$��:���=�����Ӫ����<V����_;���%��=��]���ۼ�G5�[	�=�<f`Ȼ+s+>:b�O">J.c=V���M��->�=�9�<*HN;`�[�Sj���q��}��;NڽS5F=��=��F=K0��̵�=��Ͻ�e�=�9>Q�?=!��<c���7���έ=�柼a+�=\e�<\�<&ם�og<��r��_���>t���s=�q<Z�3���9�o=Q�~�qL9� ��� >�.=���<#��;���<��ٽ
us��]�K�'�t�f����= ����<�K��0<�.M��{y�PP=;���+�=h��=�ʽu��7���~5����=�y.=q�P�6�> �P>鯉>kٽw�?� �ҽx��F��n�����,Q��z��̱�z��J²�ߜ�=$۵�J"g=y�>��g>�݄���L�x�=����7ý	��/��<��ٽ܂�b���9�B=:�=���R�=Q=F��=.��=��y�[��<��>�/N�+�*<%�&<���p��<~��<��=��<6$��ҽF� ����=�!�=F2�<�"�=�h�</A!<�[e<�F콦�yeb>zu���C�;��߽؆�=z���r�<�p�0�>�Ւ��7Q=�{)>!F����~�Z��F&=X������V���w��u<˗�?��T����d�==��=o�����Q�g=ѝ�=��=y͙����=s��<��=�*�;)� ���]�=}w1<��%�ҝ��o�9Ѿ2�f�E>�#=�B=9τ=�����=�~M�h���]��฼�o�g��X
����=��ٽg$���{=Q�>��>�k=�*>B!½�q��lݼ�L:�����D�=E��Ϳ�<B�f&�;�m�=����;H�����=}Jʼ�E�^��<����=<��!>�'�=��o����=Ȑ�<qü�W��g>aK�=�t��I+>z ��<��}�����=H�X��'i=;�=��K==���a�%>�n���>�rg=6D?�U��=zr��0=��!�.a�=+�~��J�<&����'�d��=;���d�l=��w<3�������G���=$ >���<F�;f·��F�<�?%=2����/��=wݽ��9�R���'�<n�&>���9��\������;��%>.��9Ž1�:<��g��e�=,��<P�^J5�;f��GD<���z��e��_>e�=�G ��L�����K�%=�/��x@��tЩ����=��=1j���������=���= �I<�ؾ=W��=��%�et>���sc=�GȽUm�� /G:`N׽6�B<�@�TA�=PWP���c��?%���=�fn=��;��> F\=Q`4��P����F=�´���'>�۔=�=�_����%���=�D��D�1<r��= ,��Cmջ�����=GZT��S1���=����8iu<�0=�g����=��>��=��t��H�U�Ѽ
��yI=�_�=Ġ6���ռ�ټ<-,��$�������=���;�|=j�e�^�'�Y�c�>cH�-Y>�H�����=�g��ѽ��<Y�����i=T�=�s�;Y����i=h��Wȴ=7#<=�Ɛ=�>��܇�=��|<D���t�;=�?���"�'�>����l�Q=��9�.:���)7�=�̄���<\�'����3T<7z�<�}|�����7��<�W>�	�=|,>Z)+>���q���=�}7<|�=���<�"=��L<m���~7)=w��=@�ռe8l=��r�����I�½��k�j����>�D=���6G6���
>���=�Ի�I����=�=��*>����N<�:�����
�K�;ƽ�)��[�����=��|=A�=�衼��>���=]��=7�K=@���9>;|ŽUI�<Ž��w�=��m��4=*_��P�,��˭=�q�yP;��5=��ụu>?V�<��=�L��P��<���='=��	O<U؄��n�a��V�M<_�Z=z:�=�w�:�� =)��=���=w�?�aSϻ�G >�❼#:�=x��<1��Z`ּ��Ƚi�C;*�C=y$ּ��t�z�W=�2�)�=�ڄ���=����r� =y�:=�[=G}	=]�����w���6��G�<����ܒ�%u�=s2��q<mK=N䷽����K (>���<��"�_CY�[>��x=��˽Uɪ;7�H�s���{��<���=��ʽcu������|8=Ť����<Q�E� ~=v����=F޽&
���#�D"��ف�=����/�S��U����uu���c�=�핼�m2<���[E��w��K�	����=`��=5�->�= +¼��h=,�=�������d��q5Q�󀞽�� >�8=�G�=�CQ�֯�=�`Z�6C�<H��3����u��Ĥ����=�Pݼ(����4��`0��)��9�>�
�=�P޻'3�u=\7��7dg;��໭b���Z�����SV=w���f��Ș�<�X��O��2 >���=�x�����=�T��LkŽ|H	>¼н�3�{�=Π�<<�=(�N���Ӽ�@�=�u�; �e���>F�~���=F�\��m�=5���缩_�<��=�#�=�JѽX���\2˽�?>�¼�μ�W��X�c�	V]=����<]���9k=&fy�y��<f��:�=�Sc=m_����`�<���;Z�<�8��ƽ�>��N�V1�1��=L�=a����6:* ۼ�L~=M1���7�,E�=�e��L��=a�A��J>�kw=���"u���=@ӄ>'�>[]s=`�ӼN�1��9=#ue=�p��ژ5<�ߗ���<��=���=i�T��)�
�༨B�=G˒��g�=�ܶ�r a<0fR=�θ;�먽ȫ"���=GL�Q��;�T��#ͽ&�<�(�<�>�d���yG���
�����k����K�F��=Dj=݂��=���V�7=d6J=��;|�=훡�QK�=�ʼ��#���8=�i�=
Y:��ͤ=�
>�d��{��P$�V�=q��<�`��꿜�$s�L:��^Q]�s�=�O=oj=]��F���ݡ�nǽc=a���P%><J1�(x�����=��K=D&(=7�(�]"�=�b>�0ӽ��O=Ri~�+1�f��<LN��6����=E��=���;ߵ��YFӽ�I��n�P;k*��o�<X~�=���*꽧˛��ݼ�Ef�����T?<I�=D=�O=�e�=��O���S��9;aM���Q�=�>r���=9����f��i���ʞ�<!���\#�f�=e�=󶀻�V'���5�:�k�=�ِ=�C�=���$�X��<��=�o�^ܠ=�9�N�P�{��_V��"f��~_�g
�=jX��`JH=� ��o�=X!׽�rW�{;>�Ĺ=��3=��L>�o�������<B�Ҽ_�b<�]���J𵼟$>�q��=-(�<��<4�<���=�S���=��1�f=�$��3:���<u�����?>��S=A`�˛a��oU<��=���� - �~9��-���=`RR����;�^Ի��ɽs���ʑ<�9�=��E<�2<�3�=~��;�ֽ��>��h<�ܥ="�'� i(>[l=&Z/�..V=���D��=a]=��=Ia=�-�<}�:���<�{>�� ����z�է��}���B�����; =4E7�B:�=<��=�aຽ9Y���k=E���Б=i��<��	��=���%>��=���=��=MZ��+��n�����->.	��)!ػ��>�U�}^5>㓓�{��<!���HJ���=8�<�A�=k<
=X&?�eS=A��=�Y6> �4���_i=G9��{�Y=`8R�X]>�#����=:"	���_�����ʶ}�,ۊ��ܿ����K�⍽_�G��=���=D�<=�`=�\;��|:����2�<f�Ͻ��>�ݫ<�;C�>1�=W!D�+�[��I<���K2;��7��<��̲T��Z��VH�=�����?=�y�=:��<%��([=��=�F�tL�=���=��=�+>O��L�H��sl���=ly<����㯽�7�=���=���!���5��ٻ�T��`N�aT��RV�<�<�p��>���#A�GB������M.½�"7��S=�:=O��=)�=\��!&4�6��=@���fBp=b�=r$ =`j��2�	׵�7w�=��_�-�>�DA�P�;��%=��F= ��޵=��<};��=�?��Z��>;���=x���d�:!�o�zʄ=�w�=l���$��<J�!�<����i��; �=`��=�M�<#��=m�<�QG��j�='Rf��S⽋51��%�:U,�<�:H���T=l��<A�=�͉�_,�=C�����Ｉ�=�B�`��<�5�=ஒ<x�=�/m�2&��^�L=H�<�(S=�e��xe=ﵼ���=&�]=��<!�d>9�\�^$��DI�W��a�R�	��<��<��n��">��= �;^�����	>�ʵ�j ��y$���2�=����1�=Tt=<�={�N����=I�<L��<�=kq�Në��Ð;н�ɸ�o7�X�мF�6>�֚=�C�=����=�7=�۱��0=/Hf=\,����>ǩL�ʉ�<?�x�I�	>r��v^����>i'ݼ��/���!>%쪽��:"��<����+��=F��KM�(,���Zļ���v����=�L�=�DϽ�g�=��*>��=ן��\,>��s=41���zu<9H<���D�a�>��]<��>-
=ou8�X�Y�*�'��K)�E(�=}��T�d>�>�=��a���\�|�w�fǄ=
��=jලE*�=$��=d1��Z,�=�8۽�ݽ���=��r�3N=��O��	<���=F"�=�Ƚ8�"=$�I��֞9<D�;��=�=�%�;���;9`=`T=�,@��s�:{t��M��cyn������=�<G����O�ݗ%<��%�q����4���a�L��=H�#>x��<:�h��={ĉ�^��������1=�)�<{��=�}�&#=��=��ǽ��J<�Q��܃!>��;�OA�UĀ=M%�=��<b����L�<3=
n�N��=R+��]�=O2>�Vս�T��j��0
A;����f=�_�:��[���<Q�A�/=�!=�=gb~<��=�D��T�%=F��=gU=V�"=\w)����00e=��=�ż��,��/�a(ད������Ft<�_<��m�R�0<�����!?��V�=V�ӻ�~y��#��}/�<�{<~S:=)D�<h��<o�u�%�=�/˼�>��=X�C=����T{���=.b �
��=�1� ��<{#�<�3�j=p�]��>��[����<�A��B���ڗ�g!��=�:��ȼ0���|����=}�=��?�$�Z�Z��HY6>QE��
���"���\g��D��fU=
���QSU�^6h�ฎ<�ƽ�������=�G�L(�=��8���h=�G���">���;2@����<�a�=�=;�槽���=��;Bڽ���4=,w}=m�[�����]�=���=l���'� 9�<D�(��4>DB�1K꼦7�=�E(��^?>��=��໎Ah=��=��B�[\�=���������=��!~G=o/=)=wm�E��]G�=Ӕ>��	;��=�>>���=�Ga���=M5�=�t���U�=	|�=���=�4x<]<�+M�;��s��ͽR0���j�<A�n=7`�=.rM<%�=��9=nF'����=�z��,�>�����8&=�7>#̓��FϽ���=r=?;(�ھ�=S�v=��|=�U�=�.�<J�.�5�%�@2f�K�������	���<�T4=�}=B���!#���=�"�=j��<dbV<x��=�{�<Ĥ=S^����=&(�=������:=r@����=�����f7=���=LL.���<���=�@�����<f[��5>#����5=����g���[{=��>P�y��<���=?ꢼWx����+��)B���z��7�=�\>��=��<���=3 Y��d��F@=C���{���*�<��H�2�ͽ��4=Ё���ӽ�m�<hRo=���<�%<D8>��>��L�=�g�=����G�����h�:*C��Uu�_�><���ħ�<��#��H�<�L���R�b������:�"/��#>��= ]�;������;媿��dL=b�<�l5�:%�~'�<��ƽ�\%�X2�=��l���
>����2���wK�� G>�N(�ƾ�=q|h=SV��Ȃ��l=�/=�08>��<�-���]�LٽP�ҽ��Gι��N�q�̼�k�C�<�c:�C���=�=<e�W=ThJ��A=h3���'���<X!�����?4�G'���i�  �<B̽�x���{�=z8��"�������<��
�����ۑ;n��=x�=�w���ڽo��� �-*�.��=M�=U?a>����t�ۼ�_��ie���½�m���� ��v���T>��<۫��D|�H�#��R����=�Ľ�a�ӟ��޲=�d�<J=<ȑ]�V>/�}���
=t�n=���᥽�-�E�3@5���<���f��"��<��>��$���G<;{}�[/�3����aE=�v���E<��J����<��I��:�/�������̼�R���'�Rc<es<���=q17�����>��KS:�.����&���m>�]�=F=|�Ӽ�&���9�x=���<"�"��>��O��m=a�;=)A)�c����%�=�s��<J�ܼ�0׼*Y,��F���w���t�v�o�]��<W��<�A=���v�->�����0���I����lz�ϲ<�RG�fױ=���<u���#�=��(���8�����L@����ܺ���@��<pt<≽�%����%�N�>�Bj���=��ռ	�e=7�%�uMb;��g��+k����Q-𽞔�<�I��p䚽5(<>��,�N<��<a�=gÕ��>�=a�<\ >�s�=.�o�
C(=QM&>���<�U�=�y���C;���< Q>&�	>Ǆ=�:�=��7�ѻ���S���ǡE�2(½��7�s^�CG�<��)��v[=&�{�&�'�z=	T˺	��	=��:�u���<:)�=����i���%;?ْ�ߖ>�����ҹ㲌��0�	K½i��+�5��G>)��=��N�-�W�e�����՟+���=���Y��=oa��}�=�{Խ	 >������=���,���C������^�3��4�=�X#��A��O���t���Q���н��=���;b��?�=gIý��=U�0��<�����=����,��M<˕ͻf[�=b�׻o��=_�;�A���\�<���|>:��9�m8���1�=H� >�P.���J�=)�J>E=����D�<,�0=]�=y��=��$=H9<���Լ�=�����!=�0��z�|�m<ih轴Y�����
��R*=t���Ό�9�Q=���=�i��K=��,=(F�<���=t&�=ց�<��'=���=�,<?�>�������i�\��%=��ؽ����!�<�P�:aý��N��"�M�m=^��<� ǽ�Ͳ�$"�=�{"�� &� ic�P�6<F �<&�f>7��<�x	��?7>1�2��gX=���X>��@=.�NF=�������Xֆ= 
���E��t��<���=�;{=��G�um�U�ۼ@P�=@��=w��<�gY=妽��ȼ�8��G����f:���=}��<;-��;_���x�v����_���q�#>"�U��½ ����P=�챻[�=-|<���;���7�{>�+Y:ɂ�L|�<$���s��J?C�f�=�=�M޺i��>Vw<�+���;&~���L���=b@A��'=���*
�A��=J#���:�\L��U��1Y>[��L���7(=w9��1�齜	3>M5E=k��:aq�< �9� Oq�9�W�n�R<�G�<��|=��=d>�U�<Y��<��E�=�(��JVI>�;ü`	Ҽe�>)M[>���< \ü��A�U���4��4�=Oeֽ�ٯ�n�?���@��� =7k=lD޽���H=��=��Ƽ`�v<8Ǟ=("Y��@���׽���ݰ`=])y;�>���=��.=̧�������<�=�I>w�,=��R����<����'�Ѽ�Ѝ��#M<~b>��=�-<J�0��XI�Z�=󚽍⧼4�<0��=���=)�=-�<E	ͼz��CԳ9�v��;����=����W�;���<k�&=ए���/�h|���'���<]=�<=u��=~����(=;�=U���-�@�Vr��0������:Q>QLŻ��==�s�=���=����h���H ��>�D�=N�(�Զ
>�=r=�p=o�^=�Օ��U=�C~�ͅԽ9һ��=a�>���=>j�<־9�B_������<w�
F�<q���`�=�8�Ī�=id�=�X����<2��Y�=�м	;��8�����=�����u=��½�8c��2�3���x�;p�j=�ٓ��ǽ��)�l鼵u���Z�3�½�s~��
>�����7\��{�= �߽L0�=���<���>�o�=u5u=x��5�=�M�<ՆS=����Z�;|ʴ�<��<7�>��j�=��]���A�q��0=0�R��`�����PEP=��<G��=�� >%Կ��r�<9��λ��,J����S=3G\�H��=���=�#��q�=��d<&.=�l�����H)[�0:�4����!>F�-��9_=(�v=�8���T[�=A��=P(�=n�.=�����E��o�<�"=�mD!=����.�0��n��<=v���t�ǽ�ϩ�.S�dZ>�1���?Ľ�D~���=h��?<Y���4=��H=��������2�<˥��Q�����<ۂ�=.p�=���;%@x=���;dH��)�=H�?�|��\����=y&�
�=�+����>��G<�:�w\$=��$=2rS=٦��==��>�gƼ(_��',�;}U=��=ȼ-���=��=�^n�� )�����=L�>Eꇽ��=�E�=ǣR�6�<�@}=k�=@�x=(5>׊�=X���2Q=EA�̓<�=���
A��F�m�>�aD=��p==>G�Խ�_��[T�<RR�������<��<n���뇽c9:�F!��>��=6�=���¬�<���DI><��=�9@�2��:��6�ڠ��ǽ|�=/�[=\���)�P�8��[�G3=�c{=�*Y�7���>f�=�w�05=�Ct3=N'q�L0��}�=|fU��;��D�~����<{x�=e�Q�`#!<Et�=�(�<�>�=i��6>ӽ��<�1�=(�<b�=9�=��=/!�sA��K�=�=�%;=����2=8s�ļ�-=>��N�jE�<�g�Q�e�*@�}��aA��G�}��ֽ&���F	?=��=����#�=��<=8{=8�ѽ=��<&Sؽ<�=��>W:l�Zm=c�U�LX��F��=��H��XD�ɗ�=�����>�?��
/��U)>j�N��˽2� ��l"�:�����*�b�=3>��cq����E�"�+=�6U=��=4M�=4p=��q=b-	�~����+�-�(��n>�#=���=�~�<����= �wVټ�]�='��=<�O<v�> ms��A�=��߽�]=ٿy��ʌ�O�:�G&���Ny=Q1󼸜�=�h�����~��zb%�m�<�B�;6�Ӽ���(>>��=
'�=Ԗ�<����=��=�w�=Ѓ˽��>�V;=Z6��m��;> s=���<�Q�<4��ۊ�����K1>
m�=ŽX׽1\�E/��ړ�><۽��=�0(�s��\��~�S=y�����IS���M�=8���S=r0�;PW<m�=�A >um=��T=��<�ޡ�X�����(Q%�S��Q��Ҽ�x�=�H�<FB���	=����7�����U=!� <Sy��ȼ���������<����+>��+��=�d�����v�>-�<m���N����=M���~ѽ�<+C/>��	�Y�:}K���e=��'=`>�]3=e��<.�=��ĺZq�)�ͽ%�<�8�;�AM=� A="����L;�is=i"��ڲ<�J$�9?�<!`;Hď��@S<rI=��"=��ͽ�?��A=P$�<jМ����:Lf��:�b��EW�<$l(��6n=<i�=+U�<��=�h�ֿ�=v$]�͡�=�FO)��z�����$����B�/���..�!�U��To<��=���<;�����>�V;�g���=0\��'Iv�̊X>���_����ݽ��:(Pa��	=@n<=k�<�wa�Zu=�]��$�=#�=b'=�# >Sx�<-�C��Q(�(k;�hd��� �<�#�����<&�=��)�v��=�x�=��~�[�=���S�l�󚄼h���T
�=�)��*�;S�@>1.�����<m��e�nwS��R=㨼���=i�)=c��Up>��i��8����ٶ=O������m��={Â��@��X��ŽU`�=QT�<����%��<�(`=�l��y���t8=�(������S�Aw�=�� ���=W��T�:�u��=��=��5:����;s�<��6=ܛ���h����<u��<<S�� N����=�h]��	�=QCܽ?��<�ѽ�|�=B[�<�Y���y�ļz��;i��:>�&=Ot@���K=�h���@�=�"+��<4qx�+3�<j��=����Ō<H꼄��-�ܼ�F���<��W�"v=Q��=�྽	sw�RJ=�-(=�9r=���^�˽��V��^�=C�=�׻S7�=�&6=�f�
='ez9'��=��ڽX7ѽ��2=��ܼ�Œ=�����=��e=d5�<\��g8��`�<��>.0]�1�I=�|���0=&�ۼ�!>���6�;���=ސ��%�=�gJ;C�=����\ ��x.��L�H��D*E�{���7�W=��z��>7����q�n2=�X;�c�=_;���*�<>{{���=�}*�ߐ�<�j�=�Z=be+�9)��2֢����^�X=�u�=�#�=Nw���ƃ�R�W�Ж�;��D=g>S=�a�S���i�=l7���ͬ����=��<ưs=I�o�,ͫ=͈������5>�w�=et�;���=3���ct<O�=^t�{��;>%=*x�	{ܼ����X��<ﻕ<�{����Z=���[�#<�%�=��<%��Mi�5S=7���A�C���>=�x�o��b�=2��^FY��ҷ<�3g>sR��@�<ך��.��y}=�̽�?����c�!>��[����<��<)�+=`�	��!=M=(�;��N�=��=�,���HS����<-�=�c�=:���?�=�t���	޺�R��<���*���(����:�AY߽!a1�@>���T]>C�3>O��>���=���<q��={%>�z��bW�7>)�=+�+=����C�=䶵��і��[=�%Z7=u��;��A=6���@i>5���ra�V���Rt�P�>sH����<ʰ\���\|�<�\�=W��$v5=�в=8!>󛾼�mK=����=�D�=3�5<^��͘g�..e=1����t�<.9��]��a���v�e<�lj<(� =��6<�L�=H�E���ڼv��T���p*>�iҽ��lr9=)Ef=�V�=�,���# ��[>y��n*��g�9�L�;|������<}�s�X�L���,����&_�䧼���b�f:��b�=t�=�臽�D�=T��=Z�Y=L'�� X=��_<ƫڼrl�=�ｻ3>=�R=��e<���<k����;B:��^���>7��=wS�����=֓>>�r�<�ڼ~�=�<]�u!�=U�=��0=��;Q<��6=�̓��<{=Yf�;��=:b�;��P=7Iͼ�^F=�=�i.�����[�Gb�<H�=���<��,��:=S���=�(�<.��;ԗ,=[W�=��e� `)��N=]=��M��o�-Mc�z�>F�IV��M�m=��=�VA=[ >Գ�=�k�����=J�Y�\G��<3=B#>w��TMg��>Z�U �9G<��WG������}��-Z�Ss�뻽��)���[�����=Dm���we=���FD�79�=��<qԤ��Vy=-]��D��7d��H��ĻW�\=?#v�4�Ʋm�䭩<X$�=������Yh��i(�D:�=���=���=�֎=$xz��������
<��=��W�-�(���X��(!=���=��������_�ܳ�=�j<�ü�۟m�~�� qH�� ��<~!��Q��=����vb�<#{
>���<f�^>9�S� =�P�v�ܺ��?���ӽ=Q�cX�[J;M���u�#w >v�t;1	���Kܽ�٦<ҩ>��н@q�fmI�L�={��;�v
=7��=�<<�k���/>xq����=oŽ����h����
%>0�N=%��%�B=�h�<�����ҽ��;'�D�"3�<�{F�ez;��S�N>���&�p2�=�)��W`Y��(��	�=��=�h"�4��=�暽�;��i2�<	��=ZBg<0Hc>ԛ��D5���
>�1+;/��@�=e`�=
l��h�����;͵����a�sޓ=��:�ռ��T;�L�<x�W��(�<ݿ=x���=�[n=�y>���$?>��<9��=v���ȹ�<���=6�@��s�pe����=��=�/3��S�=�����Ƚp(-��F<�Ͻ��<�L�<��� ;q��� ��
��%5<1�W�6���c=S�ݽ��;����p<�u�<K���*4={M(�Q�=ZQ7��f=��R=k��;x�ƽ;�%��+��E���I���'0)�qi��C�<Mܼ���<Ң��O�]>v�=ȢýX��=�q�<�1=1x�;�ٽV�=.A_>� ;��=��<D{���O�<0�!���)���e�0�	���1��vz=jQ��.���B�=w��=�{��;��C�=�P�=�I;=�^&����=4��<���m���1= ��;���=�������R �#�=�Â<�S�<�ʤ���'<��z=��[�`R�<j�09�0V˽@k����D;"$�=1��<>��+-�$
�Y��U�t<�=]t=5�ؼf=�=}D;n�;�����)W=���j`k���𼡺��Zq=��=�E�=_�ӭ�;gVĽ� �g+�J	>���=���э�<��:�;>�E^���2>�p<v��=p���j�=i�����p�>����=6pս��,���Q=��<�<x�~����=7rμ�lŽ���:uo�����X���y���=<�H^�'�#>KΎ�NMu=�i�=�$G�E��Gޝ<"��=���;q,�S����a>�o�=H�=x��<�3X�D��=ͥ;Ϩ�<��Ú�~t�'4�;@�=�'%>������=���=���S����&=���=��=���=�b��A�=ua�;7��=㶯=�O�=�Qe=�$�=l⁽� j��WN=��{�WI�HOn<�Ո=TP=�V��n��=�=� ���=�*��X�<uM=�nx<�����9	=�<���=�C��Z>v�=�ü��)�n���G�=w����#��Ű�/=T����9=�4w��c�<�/��j��}�D��=��,��~�Q��=.A�=�2�Aee=7O��^��7]8=�5=Ĉ����C;�)��~�ýO�=���=SEt�ɽ^>���»�*� ̝=��$�ԅ�=Z,#��+�< ���w�">A�W��5=H�!��=�b���ν���=E���w=��w�+������I�b��=��<������n=�=^��x;�!I=���CZ&���4�uQ��L[��3�5 M���G�s�J=!��d��=� ��W�<L��
[<x��=b=(���;�9Y�B���ԛ=l�������o������>,N==U��nc=qw�= ����=-9>/_r=="�ɻ" �=7��=�K=�����=�5��Ɏ��%�v�μ#��#�Իy�<��n�yڽ�̽�A=�I��P�:��
��8<v�9<1�S�@��=Gd�=��>
�7>"���A�0W�o��}�=�.=���;'��:�0�uA�<oku���>h͔<l�K>�U�=z�*=Q��Ʃ��&��=}2�=�Au��˔<���;���xR��Ew=�<R�E<��|�XϽ�:�<}l�<%e�9`;Z�<
hb=����+5��gB=�ֽ;;�ν�ٸ�*�/>D������=�(= ��={�/=&Ƚt�(=�!`��-{�*�
>���RF>�'��Hy���P���=v�����=K�򽻩ͽ��/>�a��d>hn�<z�2>����F�<i7E��E��ɐO�?��=��2=Z�0=M��=�O�=�m�<┽gw=�4�=~F��߅���#8��A<>g��=��&>=l�Z��>����M>��c=_U!=w��<0@�<&y����N=�=��<��ར�q���=�r.���8 c�
`*�G-=sĽD�����8=����>-��=w��y�=�I[���c>`Ε���a���<�Տ=��}�)��;��\=�� ����=�ռ��=��=h7>�o���=z0���V޽�4�<�?˼6oY>�5E=�?K�'�=����;�o��=���h�%�V��̭�g�=�ڇ�߱�6����F������¾��=b�^;��������=>���e>d=濋�F��{�>yϮ=l����=)�>U=���i������T=��2>��e��n
E=��> ���=e�=ںO��l��p+>��1��i�����?'d=�W�=�Q��V��<��!�=_!}��5<��:�Yw�=U�U;��G>�#ӽGc2<�p0<��)�g=�ܦ�נ>:�W��j�\���ƽ?��<���m�=L��=d��b��I�5=���J,�=e��<L1���#�;�����i=��3��=�>v=g �=gՏ=��y�+4���/>�̼̽�CW	�F��������<��m��>~٢<l�c�R��W4>�I�v��=-�{=pV=j�=x�h�8�Ľ�(;=�Q�=	E�=�l=wt�:`���!W����=e�=��<盽�
�=6�<��%�U��ī=#q����,>�Fj;�)�����Q%=L>-��;�ߋ=�M2>���Dۻ���=&���=���;��Ӆ=��c�갈>%���y/>pȸ=&b.�q�J>Dy���L>v���� ��>�<1^=;G�;*hg=IN���z=QT�<������"�=>�ｎ?�=}A���=�����|�i�}=Y��=Y$>4S����)=�$���ǈ��P�< ����&����.=^�7�=,�?=r��<ʢ:=q�>Z�.;�4>KNc=�SX=�g�;K����	���v����)>w#�=5l�;��=7(-��$=�R��Xż�?R=��=!�U��8p��@#=��<�tL�5>&n=�5�<��O��7=�*̼ZM�=���`���cq��j��a�c��ۭ�c�M�6f<�&[=�>^��A���m=W��=��=�N@���*�ع>�ؾ<�<6�>�(=��K=�4�=YEZ=�K�=)��<Q"��3�E=��{�P����p��v�_�T��K>a�=�b}=G�ջ�|�<��k���:���n7=XO
�%ˌ��mq������=;e9�`i>*%>c�p< 
��D]<��^<[⹽��3=�p��J��=���#��W��=G�?�1��=_|�;H3>�9=ޗ����������H:<�vi�4�P=��;�1��=�=��:.����Ѡ=�w���8�bU4��᡻|��|J�=���=2@�Z<���n�=)�5=�_����A=A���>��D&�=$�ͼ�>���L��:��`=+��=5`�=�'>��/���ƽ�I��Dȷ�q��+H=dlo=�Dߺ�C�=9��=d)�ؖ�<B����E<�׳�w{�=O]�M>^�t=l6����&Ί<J=%��6x/�SD=��_=W\q��T�<M �k^9�<��������_������S��;o��4oz=��N��+\=�f��qk���M��;RǛ=����摻O�ϼnvü�1c>a�[����(��=��=�\=P��\���9��<$lJ�$z�=�>=҉�1��=+&�$��̡_��v���<��=l6=ӑ���$�����<0O=�h#�t]ƽ�-�<�X̽+e#��8��Ћ�\Z����=o�;1)��˝=�=������<{~��q>w�"=΅G�'�����=D��=u.M=�s˽��ƽ�A,>v%��Er;��E�S��=\;�=fy>���AL���=�ٽJͽ�ѳ=��	;O7<�L/=̷�=�P��.�)<�����V9��f�=���� �ܽd�%>���>+���mɽ�2��lཅ1���ᐸ/1�*�=�\�<*�z��f>�U�<0~=�V2=n�_��;���Y&���Rս�+���E=,��=�ҫ<�>i�=�]ȻZ�>?l���Ǽ|�o,�=��k�	t>��;ܑӽ1�->;���OI��4΂�h?�=G�=�M(=�ޠ��md=-=>-0��0;�P������|����=#�B�q2<+��=���=�P�*K@���`=�%���A<�v�������-)=m0�<�%��=� $>��u=���;��]=��3��v�=��s<���=�*w<7�P=|=�:�%�=�c��e�*>�*��r�����<Ѐ�=��=�B;�{��@ƽO�E=�}�L���^<�;Fm�<��=  ���>�@u=br���K��G��=�j=u�W=��,�Rg�=A~=-��=�=�<�A��)a�SB=�<@SD������m=]�V��22��<<��)���e|���սMb ��	�=@��O�r�}�콱'~��?���P�ëK=��g��r=�;�A%=���;қ��>+�=�>"<=N�=�g��~����W������<�R�=�=S���;Z������<!����(�.�r= !_<2�ؼ(>�r�?�Gƒ=��3��H=����̳�;�>���I-�<a�=�M�=Β=�	<��=-��=���m%�4s2<�y��d5��R<W�ѼBC}���o;�Dʽ�t<�@�;_���=uxd=Bx\> 2�{^7�/���%�
Z�;�����(?=a�ɽ� �=�F�<���꛼�� ��ׄ=��u= ��<A7,=IFl���Q���|=�Q���=A�d�=��<�[=� �њ>6��>Uv�=﬏;�==k$��y�D�Y=���<a��>fd� �> �<�m���>��ҽ*��>��~�yB�F9!��]
>�=�v>��>�ܨ=�M�'�Z���6�;isE>Ţ9��s�;�C'�*�P��V�=5"�=��Z��6=����^>�'=��=FV���l�c���"�+�lş�ݽ>I�>#�c�z��ﲼ�Cѽ���<��U�L�vi�;�2م;����P��j��=(����\�V:���=�=��.�=�ҷ;��=�eT<HTT�Ur=<�H�Ƃ��+R��m���+�<|�=^��<�ٽ#e㼯�2�P��<�"��!E�=+�)=I��6c5��@<�X�<���;�W=�Ķ<���=������6؀=Jz=��=������=�0��~g=��b<�@,�kK�<��>Rɞ�d?�RJ�S��=�_)���C=Vs=�V4>T'��* ���c'+�ުŽBr�= ��<��t�v9<4��P�W<���=-���Gۛ=��>�Ϭ=��0>o��=x�,<dq=�7�=��<��=�0����;eW�<���~D�;��Լ�ݙ<�ˬ<8�=%J=��>�⇺��=�7��R�=@o�qX8=�ޛ���=�>����ϽR��tu	�Φq�����-�9��=�<b9��l�A�GR�<w��,����Y���9�<������v=c���f	��˽����*��<�ѽ�:�=tb��r�= $ɼ]���n<*�&=�F]���>��V���^=sY���h�<�2�ǁ,=���X��<�`�=<��;c���
=N�Z=����CνŮ�=��Խ���=-�>��߼������ӂ��;�=��<*oW��:���1�O�=�q��;�����T<���T
�<0G��ɰ�=`���(�����ƽ4�̻�H�<~�p��ʽ>J�=�>!��=�L����=�ݼ�.�=n?�=<��i�=�\G>Xs$� e˼d9ǽ�T��
��,�=�tL�*�;�p�3t�;�=QP=�g� ��=&��=1���'%��͔=�nݽ5ޑ<`��=�@=��X��(����=��>��=:kO��H�=�QC���=����Zx���q����ҩF�o=�����7P=�Y>��R��Ў>CCj=b{9<Ә=�{�Yi�=������
�ɍ�=`(彷�<vٝ���4� ɚ��ڽ���w:>�6=�b>�+��%~=B�=��N�&L >��T=� �����=$@<�ߣ2���Լƴּ=�k�#=�L��eX��	��<Y8�B��=��=M�������W����r�=UՂ�MX��Yª�.���B��=y��� ֍���<]���J�=D����^1=�IT�m�_��n�<4g�%�=~�=S�=�R=�i����;�h�=�s�=����\���٤��=o���Cɼ�(3}<������'=�q�s�ȼ��<"r���<�}���r=������=�q=M�=��ѻ3�=y������k1<�{>�א=�~�=b#��Ƴ�jR�<*���*�!�FL�T����B-�A$��,��=˲*;",����=���=Wԕ��[	=Z>[ >D���e=ѝ⼻Q=ވ8�D�=�~��SI����=���֎�p~���[�=��|=Ϳ���U�=3���M`=M[�=���ő������m�;S,�<�;��5�T�K�2�	�8�=���<�O�=c�<HN�=��E=�=:�߻�C㽆����Ѐ=��6>dw�=����r� ��|��T���<ge�<�4<i�W0����<�x	�@��=�8v=�̮���=�B�[�����0��;�<��<��=N��<�@�=\v�Id�11�;ײ�=W��;�[����=��<1o<��=��(c>�꼽��=|]Ͻ;�a��_���ğ=��(��9�=����V`=8MU����ɮ0>?�=��<�h�<A�Y=�Z�=�V���q�=813=|�=O�����=`_}���h;tf=��p;sL�<`�p=Ty<E玼�U�x�E�_]ټ�%¼L�7=��/>��-<f糽lp�=��ͽ	証��j>���=e�W�6�=w-<�F}>�總B���u�=@��=�t���ˮ=,�=Nr��+��ɷ�jH���^=k؅����"������$-����=|�=�|�<���8=��S��!��cC�=�Y�mvټ�\��1X<��>�oս?�u��Ic�`+�&�=��ѽ��=O�����1�u���E=P)��1���,��0���b�=��ؼm�(7=�M��>��B��=�z=i�<���=�C�<)۽�F6���h���=���i;s�SŐ=|�w=��ź�=�c��#���ͨ�ǻ���=M;���<۽,7�=�5�=%�=Q��=�w=W���N�T�ܼ_�8��W=ܗ/��Rj<&��<"a��h~�g��w�}\����#���A=�І==�=�E=t�p=�ҫ=&�G=#�=�]�=�I��4{�=�g.=��˽-�r�Uꐽ#�=��X�����=m��<J�:/��<�Jn���H�y� =�i�፸;����Y=�ȝ��v{=Vh<���=U35<�v=ς�<@8v��Z�=r�(�nw=�xԼ��=x��=�JĜ�#Y�=t��=E��=���w��=����&������ڴ="��Pg<<�ŋ9J}ݼ����<�Qe�i�Ͻ�^�=�3�=#��=x-g����=]�`�?Y�=}����G��%�<~.T=Zm�=iNM���=�n>;�>�;˧=�X��'=e�<kϽH���{�=h�.<�s�ѳ���=n�
=�p6��-����n���G�:f�=��y=כ���!�����r��=#@�����$������<�{=��߽�G�:��3��x�=Dݐ<��=�(�V1>A<=W�1�z
z��<:�L=h�6�g��=X��=��</��<�	������M	�=���|I7�g��=?�,<���[�ѽ(���H�n�7��9�g��%>#���xϫ��a< �A=2��T/��)�}]�=��3�Ooe�f/��=�=���~wa�?�e����=G�=���X;>�F�<��L=�#>��=|��=̈́�<h�s>B�=��=T���`�$��@�P��.'����}�<���K�<%%=D�'�F�<���<��Ľ��e=���!�ӽW��@�ͽ�x���(>M��=����rX4=�ʇ=�h=h�=��G����^����< C�<��y=0Q�<��1<�㲼Ҝ<��>�y=�%�=�g�����<uO%��p�=��<��Z�>=�ϻ��P<t�ٽ�� >����-�;L;C=�?=x	�=" ~<���=_�ڽ�#G��r�M���T�񆼼��� ��D���g��||�<���G�L<Be��^b=�Y>���S=�e>�Y=���򡑽�x=�,	=�\E�]�	=������=���=LW�=�����1>���6 ������`=��9>ݽ|�8=��$�$#�=��=n:�<���]=��=Kͼ<�<�I��z<l���Z�=P/�<Q�<!��=}�d��\C���=�� >�.���z�D�d=hJ=�S�t;/=*M[�F��=(�f=��#>�����{��g�,�$�ȼֿ�=,�8K���qh�D��g��+̗=�oP=rwV<���<������=n�=�?��*U�ͤ�|㽼�[���=��=.�>=��ҽ��=��(�(�����s����:���<7��P7"�R�*����<n��=L�
ý����ɉ=���9q�=��F=#ɖ��1>H�)�Mլ���=��=�n>����I��=.7�SF=Η��y�W=xE���H�=V��=<w=�s#�aYx������n0w>x���"��=��i��9�;IiC=�N>��̽� �������h�7|�=���5{>k/Ž��B=8��Y���<�l�=j\���:��k|}��K��o�=6���a���[�yB�=�g�<$M�=WVt>h��=x����pS=_+�=��=;A)�&!����<�h	�U���
�DxC<�7=>��{����>؅*�@ē�n�l�Ʊ�=~�=�]c�ҙf;��<��=8x��`W=�~�����Y�%��
>��ݼ=��)>N:�=���=w;m�o�5=��0���= =�cѽ���=�l�=E��%�L�tJ�;]��=�w=na�u.�Ni���.��M=���O;�e�<n�4>���<i8�=�?�"�=R+h��H�<Ii�=8K=g=��=hk>�M�=����=Ӫ���<Ӱ�=4-�S����l�=�<
�;p1�<��н��=�&e=L>(=Gᅽ�(߽����@�=魜��s�K~7=��q�� N���0��5�<*;a��(���ɽ@q���o�=�1>�o����������=�K>�C�<l�=��#��C�<.M��qz� � >CU���F>�G���ë=ظ �Y�;��z��PN>�;>�xW;x�޽��!:r�=@e=MgI����u9Y=�9���Y�=�i�=&�=��H�� ۼ�M�<xM�#�]����7>�=��Y�
�+��	ܻ�;=��Ld#>�JQ���w�A�+���=%�='VV>!D��!����<�>�~>r�
�S��	ټ >��)<�d�a�G��0O�{�|�J|j=�t�<!�<�h=�h.�;ɽҝ>\��<��=Kۍ=�"<�8�=`d=����y�H�����w��vDȼ�C��M���;w�ѯ���bѽImp��F��:��)�-:a��fἎ�����=*9(�G�<pwW>���<x96�Q����a�<f��`����<�5���Ъ;V�1��H���V;^�=��ͽ.g��4=K���r=��=owe�ᮃ=s|�=6��1Sj=D�>1T@=e37�+^�=u��9�X�3C(�@��E}����=MP=�0��=c�ʽ_jr=N�>��$<��=�,=�������?�<�n>!�ɽw?�]~��S���/=đo=�𡺁����*>{-� !%�!~�=�&<��z=؁Ǽ����xY�׬5���<��E���(���@>vN�=u\O��G�����Q^2>��0=򭝼�;>:$> N�=�߽,>m�>�2��_<��B�����C!;�|�
F�g>z�=����V<R�2<�(�r���1X�T����c=}����ߟ=���I�f=�&<cO���m������9<O�ݽ��m=fV=�ٽ"K����_�-��=�r���MV�q=�&��N��G����A.>T���<���=�8��W��=��%=N�!�ZW�U�Ǽ6�S���ļI8�=߲���<>D�.=V��=y5=˸�=���A-l;�]>�߷�;��x�=w{����L׼Ȍv�+e[���ȼ�X����=ڂ=����&k�=ʟ�=��߽<��<�>���<e�=b[�<�S�=W�|����Y/��G�m��/�S��=�_½�>���iպ;�d>�U;�nx���.�4�=�/̽���;���ԹU=j�[�*!=04>b���D�R=��ͼd�f=Pj>c�F<� =�J!>��ҺLp�=�è��"�=:�t<����F1=>C���f�kL5��~���<`�<���<ÑD�D���p>3f������=>j�����8=E�=��ѺT%�<�$��>�T�=���=J1���^��ʼ��,������ؽy�\�^4)>^Ҭ<��Y��ڶ=��m��D >�#����=�M��Ј=���g+�=�Ƀ=�A?��;�����_#�=��ν1��<ҝ>�f�=f��<�a=K�= ���3&��Fg��`>�	��\�=?��*�8\�g����'>�?�a���7>7��<8v,��O�=�M-=z�&>��.��W�=B3���1�=��>`6=� �=�@>�	>����I��л=58I<�沼"�;aE��~����9�s�<m쁽���,���]�*�朼�fE�X[߽�B�=���=�32��;x>Uܔ=�n���<�j7=N��=T>X���$>'7=p�>|/R=3��� )�=e�ս�|=G�����;5 ><��=�P���j���5�]Q�=\��^�\����=�o"�ͤ���P>=��=Oٽ��C�@�ȋ��^=\��=�j>��U<z:�`ƽ���z�i���������0�$=��7�%<Գ�;���rN�<ԙս3z=�S~<#��=���;��;�c�<�Q��i�E�������Y=w��=�v���^�wF=!�=��=�B�=Aa={�Ľ�>��6�]:�31��<����Ә���w�C  <����,	�� b=�F���p"�y$�=��ֽ�I��e���K�qͤ��W�����a���=�>��-"��T���}=�.½�3Z<
�h�
*t� ��M��;N'<��>t�9<YS�<����a.���;*�z�kĆ����=��=�t==�Ƚ���=(3(=��;�[}�����=���<����B$�=I�	�*=���Zb
<u�����=���=��ܽ��'��ག�]=��r=̏��pʼ=��{<䣘����=&F���y�{=��<>��}��=�>�=�����ɟ�J�
=�^�<^�Ƚ�⦽��ǽ?0 ���s<x-���۽C��=���=��;O!���o���H���
=;�N=���=���=ç�Y�<�L��{����=5Y=�bx�.U��\o���ܜ<:�����=Q j�z�Ǽ��<l>��'�=B��L~���H>� >U�<��=fm7�;��=K�=.ͽs�\��	4=a�>��y=G?��׼sw+=�~m<��=*̙�hp�=�<>�=�)���l�m=Q�޽����l����:�:9�-e����ʽYF�_=����i�<A��=9n���,�;�M>S���l��=�A~�Kf;��y)<�.J�X\���:.����Y���a�^�8�$�=�
�z8>�))=ly��5�=�#9������>%�=�\w�Z8=�xȻ䋌;԰ڽ��=�6���D��=[�4>WL>\r�=����w�s��>UI���N=u͐>��=Ja>�J>*xܼ��Q�<@�=��=04,��R�=� >ŕ1���0=��B=VI���O�=���,ʽ�l���-��#�=u��<���=k�@=�K����ս�*�9ŽQ=��B�=�ҫ;���<G��<���=o��=�|X����?ν^���ټ���;O���Dg.�����5����=� {;�Z�<Iq�=8�=y>=�,��퍽k�Q�xm�q&��@�<W?�ǘ=`��/�����J=�4�=�"*=I�&=�׬<kb�:�=Ur}=7=��X<%)�J;<�7���쉽���=�H�PVz�2����:�/��� ����f���<��=����@�=�B�=��� ��=�
������	�=@����2>�<����k��	\�Mc=�h��D=��k=�(��/��|c:j�~<��<d��3=�ͽ�]S�ʿ�|���ˀ�E�y�G�bٶ��B��& <dķ�6��;�p*���<�=��}��=Տ>l�ֽh���u�������<�ֽd(�=��b3`= N5<E�z=:>ri��wM��=��<6 �<ZeH�r)��G����<�v�^��=����J!>Ws�=���T���弞��=I[��
�_Z�<��%=(���e=m���Y�=��H����=��@=:k.�ƛg�qŽ3K;�`��9���<�*>-�9���+8=#���F����;�2�=q�S=@�� ���q�=����c���"�>o�8=�[;O��<ś,=g�Q=�
��|�=�����������=�߼�����u���E<�f>�b��ez��h�,�s����q�}���Iʻ=e�>;��ａ`���qi=6��=D�<���Z��=���6#�<K$�<<4��(e�=�I�<�H<�l;]����#�<�C=�I����q9=�<�=���r��=;ȅ>?�����6)�����$���%�Q�߽�)�=L�=~@�=i?����6=�,��t=�/�<`"^�~�<�n6>��v=��n>8|��ً=e��<DlL���<����/�L�= =���n%=�N+�,�����<��3>�ǆ<V�>NX�={�Ͻ�u�;��><Z����w��J'�<��5=^�=���=y�=�]4��=u<�K�Ej:�6�n��U=���=�<ƴ�"�➥�o`����	�4VE;3܂��.��20x9�s����x=$�ɼY��a�V=s�����;��>�� =ũf��A=��	��>=-	<=Ǟ�/	=]z�=5��<l�=y��=A��;���KB�<���������	O�����k<�$>=����O��`��]>*���b���=y�l=pU=�g ;.�V���<�)������½^Rܽ-��=fY��1l���N �ԍϽ��=��"��/�=[�>��<|z�=]�<1$�M�<SŠ=��>�	S��g����F�*�b�E���ϼCa}�ϝ�<n���Յ�^��< ���)W��6�ߙu���~�c�<�%��e��F�<�=�=�n�j��&�v9�=�o�<`�9s|)=��<�=$o�
w�=���<A?���"�TMK=q��-8==�H=4�½�ѭ�����= ����S��L�<:�˻��<CD@>�D<o=k�����ڂ<Pe6�ܥ-��|3��Ƅ��I�=��=�?h<7�>��=���j�
����=��潌�5��>=���N=K=AƯ<:_H��N�"n�o�d=K/�=1�^�k>	��<'�u���;��=8�=_��<K(b����<��4=*OY�A;ٽn��=s�����;9�n=��V��8>W�������p��*�A>���s��=Q�<><��C,�;�(�9��=����s1=\|x=E2��|`��>�1E<�c�u�Ӽ�������]� >jʹ=�'G�TQ�=z�[��*o>�!=��"�&�_���]<�/�=կ�G���q����N~�B́<���e;����=��4=�����G=$<���*����<�N�d���=�¼�k佴��=������=��=)b��~�';����i���|������|=<.d��.�ɘ�=|�=�<�����r:�Nȼ�n��k=�fu�z��;6� �
� =|^�<D�Lh��4��<�>��!`�=����W��=��T=˛U����f��=��=k�.��}=��e�v��=�4>>9!�ȫ`�B��=��v<
p ��E�*��7���E�H��<Ag���+>��=�>}ܽ9�=�t��v����<X)��3/�<R�=���=�t	��B=IG���%�:���Go���ֽ}h�<�5��y����=�h>�R�==��<T�����a=!�^=�b�=�(=�
���Z����=:y=����<�=0��H�4�g�R=�ؼ�y>]����=1��=ť�]��<o��@3�G�*�yO�=��=;�x�/��<�JV��Z�=F�;=S�<�>��>���<WAu=3�轻��<AuP<S��=8<=��<�G,=�*=�I=Ep��h��3� �vt��4���V�c&=��u��=��<\����N=�-�<J*�=�.�/�>��=Q�=�k�8U7;U+>�;8�����:�F=��=8��=�(��Pi<5TQ�����{�O=�f��š�ZM��_~�=rȍ�S�7����=�d���>)l=���=�&���>�	;�7���á���%���1c=1��ً�<|���=����L1J�8�<n8$=��=��=o%�=��>h��;w=3;1�(P�ȁ}�j�=�V@�!�"��l�=�.>r<��0���x=u���z�\=� ��G�=ci����@a=�8��0Խ&>���0��e�=��3���<�_��V��2�<�-b���1=i�=���PA�=���=t�<?2���#�K�����G=\����)}=���<���ߧ\<Ʒr=_E�=��!>X>�4)�!���xȻL	�X�<M�&=2`������<��h���9�=4+Z�/Ў��I��%d<�	�.�=)���5,�Ѩ�P�<���=q�ǽ� �o;9<� ����Y�ç�={_�;���=b��<�W����ҳ=��ڽ�H=�ܥ����=�L�s]=�==P�6>��߽Π��Qϼ?��W����#>�=MK�j�<`��g�Ž�#=��N>�O_<	'�=l�><���=�vr=&��<+�>n�p=�򤽗�n���=�n�<�ft=h��n	��C��a�a���_d���A�Vm+=��>�0��<�ʖ�;:���̽l�*�yWC��>tn>^*)<�U��ǽ�H�=�=�\x=[N=d��=�]=S�P=���A<��۰<5>�W<���<�;y��)�=�f�=4�Ͻ��$=�!0>�lp�{��<~:<[���$�C��<���= >W��<uE=`2U=�?�=s>l�q;z��c�޽�M������7���=�{C�̸q���k��cc=�W���.��3м(ܰ=��|���C�o�Y�}|�=z�=6�ȼF�"�D�=g��V��@ϽH���F>=��=�}=r�w=�
#���r=<���>�����=�t>r�Խ���'�����=� U�d ��а��&\��/�=Z[�=H�=���+H�qBj��F�=2�c�����=�����G�)�*=��!>��>RFI>j��L�H=���<�<�<�!�����H1�;3��c�/�N��=R�w=�=�=��9��a=+�̽����a1=�Ih���T�*S��+(=�������+^<$Xν�>��#�=��=���=�>�=�A���R����<M��߁;U�<�9r6�rX��d���p��V���ּ#��Ԡ#>�����]����=�,����=Z�$�҆,�j����7����=+�r=��=.�ȼ{�U���=��T=�	��蹽�=��<��o�yz����^=-~�&� <���-ud<2��=��<�Y�=��]�^�V������>�=�����"<wHg��떽}H�=��żS�!�a�f=�b�=�$����=�&�<��޽A̅��&�*��=Zi<~Z���w�<<i�����9���=��=�d=B�=0�v=f�=��+<�(��&6W���p�u�l=���YL�� Cm�Ɯ�=�!>h�w=�+�=dO���|<��}=|
<a\�<Œc;S9>=U�;�-)��6<w����=.��.�<_��<��<�=�ϗ���O��K�=��~��U���6 ��s�D��=):?<�/d=��==�MO����:DP�=Y,>V����*�BR�?����ƽ!�=|��<h��<< );_jH>�'C��� <�D��AQ=�#ݼk>�;�r<�ǵ���%�<L0�4cĽnCC>�
L��+���G�=vb�S�&��d����L����=c�=��9��"ݽdZ<u:��C��+��=H������=��<��ps�;���T&Ƽ��z=�!����r=����.���Hý�B�N�N=ܨP���Ͻ�,�=]��;��=1��-#
=S�=�|���3�; ҄��\=@ۑ�[<?>%!=e�1>M11�o$��Me�ƒf�'�j=����|��-V=�����Q�w��=�t�����=9�<�m[;�@=|�>��-�(�����=�z��4��k4=M�<�x���]=:��
Df=�Ѕ<��Ƚ\�ּ3����=�Q�<֥s��> /=7V�=������=�}/>�f���Ҙ�=�=սʽ%�G��F{=/�=yVR��\#��=��ͽ3I=q��=�\=W_=\)�=:=��u������3C�=\����/>�O��i*��5�=�~=�0<Ʃt��,<$^�=y�.�e�<fz����|�k]<�w$�b �=j�%<�q��w�=���>r��p�P�ۦ^��RJ=�B+�I3��u���8=ʗ���̼ ���t=�\r��}q<r
�<�|��p�=��<�栽�E��g�= 6>��E<��=�/��������=S%���:�=8�=�.>��t�i�=��l��,�=2Y;�#>h�l���E��t�<-�����=��y��o#��N>,#�:��<�@�=a��<v�A>��ټn)�<���~�V���Cc�;#
��o4��ܽ0BZ=��F�?�o�u�>pę<A��=����:;�u�;�Q�=(�=����<v��F����H=�H==�<n�����(��=_F<Jܽ�g
>��=�X+=��<߱�;���=+��<�l>��Uq=Ai���T9��[+=���=��3>/�6&Ǽ�������<���=�Ӷ=���;r{�= P7�J�n�
&=!��<�Q�/�=�Yc��Q`>�� ����Q��-�:=|�'�I����,����������u==vR�S�>,��B�A6?��Uq��̲�2��F��ǒ��zμ̑>E�>̽>P��=��̽�Q=4�H���=]҇�7�O���[;~��|л�$�<�ki=BS=��0���>ȚŽb�+=�+=�ֽeLռ���=C�=��6+���p=�ac�C��=�l=��E��-��)۽���c ��6��E;W=h�=��.��	M>~��JJ=���������=��r����<?����V��+*����o�=���<I3�=��	;#��<4$Ͻ��=o�<��'��1�=g਼+3��@�9|������<3�<�&�<C�(�[g�=�!>�R>;�s���=.��
��ٶ�S1�,(�=�X0�M����U��p�=�	"�$X�=�`
>KS�!��E�a��=ɦ��Hl8��=ɔƽ����ȿ��3�	Qk=�l�<ÜN����<���=ج��3�=e;E�}S�N2t>ͼJ=(��=�����f>�r*�Q������x<=#s=�~����ػX�=�*��ń�<59)>Z���f��=��� ���Y�<�xl=��>%�=���=bL�=�����7=5p��X�=G�N<��ͽh�^>.!w<�D���n���1���Y=��=�/<$��<�0=��L�0/�=�ԃ<��>b��=�h�9��2�}β=��e=�$���G�Fd=z���"%=kM=5*b�`�=2�R�lz�=����<=���9t�=h��=v���LF�W=r=`��=�м-��=[D3=�*�<�v1�Y|z���=9tܽC�Ƚd;�=܍M=�	��7h��ҙ����=�=�*s��ɱ�L��&�N�y2i=0�.�;��T=�x��4�ۏ=���;��; >�?=���=Z}��P��==�o�e:�<[�<����z�=)9��eG+=m&���j�2�>�����;��=�d�=ކW=�`6<*�;D��<XU���2���=�Z�=����V�="e�&E�=�%�9Շ=q��`���J�<��G�8K�=t>}o׼2�R��q]��U���=1t����ܽ;��{$<�y��i�t�G�H=ֆ��۽,;���I���[<h��;ڇ�=��T<�5�;�s@��C�N�=�(=�?�-<�D�:,��͘<t�j=��F<c9��;�}�A���>�<H_׽�j�=}~�=��=-�̤�=!�=�<��Ͻ�=��)>4���#=���ؽ3�'�2@�<�	C<��������:�=��<�z��	�=�*�=�eV=��=�z�;�q��k�=��}�{��o����>��=��*>�@��6<���=��J=��=�놽�]W�\^=Jɻ�T���m)>Y�;=p	e�h.=d�ܼ�f�Y�=�5+�k�=���<ہS=�w��'��=���x%�@=�_޻�����>�����8{�Dx��TR};V�¸ɊB��%#����=Jn=��-����1/(9a1>���wa�=�l=Џ��f��<��,=I����ټ��G=�\�V����ҷ����h8���3�����=#
�<PA-��o��;嫽�j�=��=~����_<V=Ʋl=AVd�g:�<���;�q�r9��P��=9�=`(X=)����cĽf&��� Q��/=딺���b�t�����<X�=}���w�H��9��˽��J�;`�8���C�=@&�Q��=��=v^�=�A_�wY����=gM��`i=d�E�A��=�n �����6=�<O�=��)����=���ʮ=�/Ž��������N���9=��<Ig�=I��<�f׽z-�=n�l�!\�=,�,>���ɦ�=�߼�;=��:e齣����C�=��E�)c�=��=�=���=\n�=���=�ֽx�T�P��@�#=tX�=n|�='M��|�nĵ�Z/���`(��ͽ$����Ͻ�2R=G���^�K=�^�=^�۽.��=X6M���<LU�=- =�h�=z�t�lRL={�ͽc���#�
>�L���(�=�{-������bM�Sp=��N=?�=	�N���<�;�|%>�E�/Y�=���<7g���/��w�GT=7��/ѽS"�=��5�i e=���=LN�=�q=�蠼�?�=1zx�h=t`E=��^��N-�޽R�T���=pk��3���a;�n�;=�<�2���k3�B��o��<�:��R�=R��=�Q3>�J����i=�i��+=، ������m-=N��qֽ�,�= 桼;��<��̽Tz>��F�ټ�n�=���we����=7���d�$�i!�8U� >e����<�oI���a��R>���<�0���=L�ཥϐ;�[�=��<�<�4 ��>��k�L��	=�;�j����<���<Ë��4��\
o���������k�.'�_ԃ<����ů��4�rd�=�f=���>�-��\�<��>�O����0>�g�=�P��>�J5����=�����H��v(��ѽ���`��=�H= }��!*E<Op����ͽP<b��U=��Q���}3��k=���<�S=KB���O�2�<l<�x�d�=�N�=�U�=�6>��>�2��<M7��(^F=(��<L;�����Ǫ�=w��=��X���;��m=n�ʼ��u�A�=���=7\ >�IS<#�&<��I��ٟ�9�=��������J=�k�=&��n���Y<��>�a<aO=M��=�M)=J�|�C�=�=!���&;��\� ���s!���& �Y �9����BO�n�H�J@K>�4m=��x=%"���`�=���_�=Ft�=�a =��h�0>�r0�]�=uc$��*$���6���>ϳ<N��=��!���G=kY+��u^��&��]���!�=w}�<H��<uhF=�X�<�O�=s���/�-=�x�����=W׽]�=:�+=�@=_w<���=F��>����":=n��;�n׺��<���<�d��3�<�<I�N=�R=�p=��=��Z��.=���=+�ܽR�<��!���N�Bx<�fu=�
�;�q�<ô�<��:g����ཁ*>J�4=��>���<!G� �D�x�x�R=U�=��\:��r��!;=�֩=�S�=;�H�"}��_�(=0�.�N+S�<��<�x��"�=`��=}�)��I=�8�=�D��v���q���}����<ba`=;���C%>�c5����=c�o<٫���4=X<c&弅�o�=����솽�>�K�<�W��D �����Ǽ����Ĭ:c�l=m1\����Q�M=���=+]<�+�=-^�=��Z�:���EP��6`>j&x�R��<���=vj7>;�ۼπ��8���R���N)��_i��v.��^��|(��!Z >���<ފ��)�r�C<,��=� <$ ����p�y,=�����"�t�=���<�P�=۠��w=:�>��>�#D>1@>�>�d���'=>;����؈�0�>x�=/}�=�h>�5�=v�=.r�=4@�Ѷ��qK��D>�SQ�~b�<�L��Bk�<��;A��=4�+>V���oY`�P�^��=\U.=�؊<<z=��=�c/=����Z
���~<�k�G�'��P="��=�_�8��*�=SKj<���<F���>�L�wFһ ��f�< ;K��4��΁<��=ū�;ؖ(<� =i�� �=����<�?>'v������;��V=�x��+��=��j�!-�����5=j$==��<3߼)<���Yu�=,|*=X�}��E��2Ž#�L����=y��<x�<Ф[;�->>��4%=�F������\a��ݡ�A:�<t�t����<��>>t�]>�X�=����l\�=;��<�}�=#>>k9=g1,:0:�<ɲ�s���JW=�ل=�� �r�=`sn=T��=�6.�`��<�'��贼�J<�%=�|��$�=�{�=�,��z/�=n��=��y���3=�-��<�&�<��<bY��wq�O���9~F���=�ޥ�mʸ=8v>ܠ�<v�=��j�^R��ॻ��IH�=�#R<qǃ<~��<�҄<�i��-);�ʽ����^<�YA=��{>2X�=�=�,ս\��=��<�`l�(�<��mӊ��&�=��Ǽ�|���8C����=�5���g���B�=ټ��q�=9/@��р��K��|�:��=3��$�����HJ��j�7=�����=�+˼����&>R��=N�<�T�=PzN����=�WO���<�=���;8���S'�SI�i>����1e�7�<�����������=�/�'.�=I��^i#=p�����=��\=���x�7����=�n�V���J��/�='�:���=M����D>��=w<�<��õj>/�X>���� 㽈� >�=V�=T=>�ҧ=	Ç���=�'�=��z<��h��=4�<	�ҽ�ș���_��A+���m>����ʓ=��<F��0I�;s��H�;7��{F<��<�<J�qn(���һ�2;�Q�,��tZ����B=�/��k僽�ނ=�K<�
�/�ƽ�r=ӭ;i2�=��=m�޽fka���=mp=�c=�t�=�6�ؗ�=�ρ<�*��V,*����}0��$R<���=��+=F\���=�g�&���=Wj�<�R��,��r�<2I=���F���ؼ���<�߸=��=�nͽ�zN����<8G�<�g�	W7=����䛍�� ߻��ؽ�K���HX��=ڽ^� ��i�=]B'� y���Nl�3�I=K1==T��pkh;~ڐ=D�=��Ƽ�54=uq�[*ҽM�H��������<���<o�*��|�=M9j�y=��;�}Ƚ=�ݻ��q��أ��,�=���=�=�ט;R�ֽ�����T<�w&���;J�;����_�;�����	=6��=�|P>�|�=���=�ц�C輱>�L:U=[A=kk�$�=<�m���=�L����=�4�%���G�>c �=�>�ѳ=�^�<`�=�Qý��\\���;�x��r���C=CZ��q�<�c��3����=��X=�J�|��:����A<
pĽϭ���>'9����=N:��^�=�0��_Ժg	D<s)=U�f���R�X�y;+	�=U2��Y���dO�f�a=�mb=��'���=�:�=��<�T��z>�����4�<�L<P���&�����<K��<���=�P���Š�d�>�E>qȗ<\�Y�w�ּ���9�<ֿ<�_����=�e���\Ž6��=j����qk�ճ]>%�Y=(ǲ<�e۽�	/�vhs�ܯ1����<�װ=e���	�L�>>��V���/�F*����V=��d�?>�>=����d>�J���OB=�b�ߖ�=X|����<���z��>�.&>���;&��;�����-�����o�;ǽ�\��=���܉ؽ�u>^6>�I0���>:��+�=�n��U�=iƓ=��O�O>�a-=�����</=�G�=m�>��<,�%��b�<��A�X=^rc=��T��Ž�Q���>Xi���$>��0�5༒��k��=�&��Qc�̫�=ί�==�ƽl�c�vs���?��P���<���r���c�m<�jϽ�S\=̖U��v3��a;�Ղ\��Q�<�	�=��!<�_̻J1��˽J������}>��#�����=��P=L�&>��=����������5���=�΃=g��;(9��r��<�w�<�N��]^!�f�C>�5|9H4c;=xI��<�-����=�:C=�Q�=t�=�2���F ��Y�=�M����J=z�<��=G#�=P��n�ƼY>E=��=��"�� ;�++�;��=×����=���=��ݺ�����r.>#P��:N=dhG=��⬿�~�=;=�p���=�u=���=i{�mxH�*�=�;��k���9>tS{���ֹO�{<��,=BD����=D߽����=�\>�<�KUr�D�:�oAU�3��=�ř�ǏF�	1��FM���$�&�=S����<D�>\t�=��;/���wT�ڦ��^��V��=�s����Fm���y=��K�C=�P>5�<�[y<]y�<4��;\��T�&���~�=-��=r��=Z1����=e��ߦ=2�8����6���]=W�^=��=I�(>OF�<�� =%��;SW@=n߷����=�����0W9�|�=�;{=��=�Z=Kuϼ�h�#)L;��T����=��8��<�L�=��;�پ��
�<�jY��j^��:��d��=W�н����a��~p�<����M<�����=Z.p�Y�!>�@��@>�B�f���S�=�
����=6�=��+�&��<��==��򽴈>��/>l$�=Cm�t�8v=6>a쀽O��dS>�=^�=�J��<.����s�=h��>Ǌ<��E>�$<��D�NeC����ҵ��Y=02 ��3=��ٽ�����>�S�=������w==FI<d�u=�4��l����:��Ev�3��L~(=$�L!�ӛ=��M�4!�<%a��s�=�T>f8�=�t;���;}��=�7�^�6���,=�]O����p���4�<��V���g�2��yB<\�=7(;)�=J��99=�={��\���X$�<��"=�&��r�;��LҼ�O.�郣�^��=���p*���=Z<=yb>O�����<�L��sՂ��������=����W��+编W��Y�&=<n>�ٲ�X�[=>h=25�=>P���?�\:)�X0&=��5�lI�<�:/�qq={.�:�p����=��>h��<�>/=�0=1%�=Ҙ�4"�;���=w3=n�}=�V5��z�<�Ɇ<��;�ȼ��+��G.�#=`>=l��<M�=+U�����=x����?�����^{�f��<�غ�:?�=uΟ�WǽK�=��L��O����&��Gs]���=q�<����gr=�K~=�Cs�f��<�)$>�=X��<��缱0Ž��㽌!�<�k@<% �s��=��>#w�=��<�1�=��:��w>?�=�Z��Z�=wD=�w���Q���9=���<r��=��5��X���{�A�t<!�n��=��w=�g���U�=p��;,�;=[�y=����˼f�=0G-;���=1A/�a������A)�=!"�;�ã�V�=�>�<�S=�c�=O�>�!>��ϼ��Sp�==/�=��r:5>��%=GG�=B�	�,=𧉽�q~=dG>~qҽ3T�,"��y�^<&��=�""=���<�=d��"�Q�ս�¼>�c�?^=�
�1����G>�D=�2��.h���=���<����>��>%ڵ=���'����>�O9=.拼;! =¢V=��N�����E]�=N�=�=W<4p����;�>�b>a��=���֗2>Ƣ�=*>��Vi��@����|��ʼ��b=d�ѽ�r�=X�:]X��C-M�Z�<կ۽�댽�#�=�
�=#�ս���<ّ2=�I����`�U�:�R�9=5>[�>肹�ᘺ��=�WF�:"ǽ8������������=@�=��S��s3�M�����=5�\���*�i�<�VQ����?�����c�*(�@d=��ȼ�q�=���<�ю:����@.>ep\=��F��D�=�V��3����2=���DO˼��>�1��=�Ⓗ��=�k���=��V==$ƻ&<���<���=@x�=D����P�VE1=D������=Q=�X<A//�2��=f��8)�=�4���7A<��̽�c����;�;=g5�R�3=�&̽�u2> �(=�'U��%ʻf��<Eؼz����`N=���w���U=��<��l��5�=d�=8"[�KR=�����߽O�;Nӽ��9��=��(<Œ�=$����,�=���em�t�%<�ҽ��o��=.��� m;'�->��<Z��7�+H��@�S�|=�߆� }�RIк�ӝ���a� ,z=���l'j��q�M<�78�<t�(=�7��4��u��ϯ�="G��a=��ֽ��=�� >����d��z]8�]�;=���<���Ļo!�hϢ��>���������=Gt���L�=/�K�)�=�}�=�l��������� =Q��=�>�]���V�=*`н G#=��=�ֶ=�I�r�=�7=Koo��%ü#(�=,T�vT�=+����M�<��ʽgPü��g�'=�:�=Ǣ�;��=�=/���F�=��=�f>i)�=�:�<��1�p�}=E+>���=��=�$d����=�5">����*=�S����4>1(=��0>s9;�������<�|����=���ݘz>��i>���=~�t;�O����<��"H��0�C>S��4`<��>SƼ�=8=$n��ݲ�i��ỽB\>Z�(��9��@A=5��<z��=���9����4�=2���l%q=��7�{>B�=eώ=4�>(d�<��������xu(�bk�=���<&/Z��F�����ͨY;�:6=���<X֙�P�n�F;ݡ!=�6=<���=p �<���P���8��w��������%86=~�J�$�*=ff���ཆ��B=�b=*p~��F�e�J���=r7�<�1�=�gf;��&=���=a=m��=��9��/�<��>�6<�5<�,= 儽?��; ��<���=�_D����=�<�=�Ƚ��;?���=�<͸�n��=���=p�N=_L <R�=�
��`p<o��(=�<u��<#⤽w.=�#���r=<=+���&u=D�g���Լ<+>&r/=)�u��~>_�=��R=���y$2<r�����=9I?����<og �#p=]�>��O��L��:�����@�<4����1>J�����#�d�=����	�p[g��d�a~d=��໼D1=۞>�Aҽ�:����8�ػ�V�=De��g@Y�|��7�S�jp�����=L��,���=�Q���?=�=���i�^��=�Uк���=c�۽K�a�9!�O_����=�[���<6H��(">���[K=�<ȼ�]Ľ��A�Q䇽���=cm�=^���+�=�)��ʽZy�8�G�����=ax��0y�=��=GK�������W���C�=�,�<���;nRɽ�Rd=��<���#6>߈����=��ƪ#���>��l�fx�Z*�W�����!>*)�0UI<~$;���!�5��iQ����=�>�+ڽ�߃����P�<WZ=����C=[$=n�A�h��ZJ��_�X�0^8=��;>^w�X	�vu=�P��5UC>nx<�	 <���=�>�=�����u��&d�(G>��=�,=5i�>��,�2�=Zo>"�G=����H�����>�?�����<YI��N�A>�-=�=����ĸ�+3��t�!>K0�������<�_�<E�7=�h�?χ<�Ľ'|ż込����H�;N�=N%��!M�=�M%�v3/�u>���d+�kn콭�۽
���#f==c�=�<x��PU������^�9ˋ^����<]/ʼ���o[=��X=n�����=;��;�+�?��=��]�e��<v=�=��=�c����켻�½�f���+i=������4���=t��Zo8�̾<������<�/���9�l���'�=l�ܼ�^���<�=�c�<�����<��=���:𺄽'ϕ<Q��<4�<�=�g�8�j��+I�����yZ�)��3o=L{���=��=k*�=&�=j�)>v��+x�������P<�C�<!�E�C;k=��	�����C��|��/�=�h��`d�A\�<�s�;i~=bz�=/	>��h��^�[�,� �����c��a9�=Kw&=ѹ�:�=_4s=�-�<D�L=lL�=#_Ľ°�H��=2�H<�����J��<A����W���������� >���s����L�=�n	<��H�T$�<�M%;��D=?]t����=� ���%�=��Q=��8���=ِ�=s�9�>B����Bܼ�Ҟ�Lπ=���<��=�ξ=5�潷��=Ӳ��+�@����=#=�=�
==6�~=�V�=��P=f����8=^3F;�&=��=.��<a6��9D�<ýX�G�>xL38]�3�@�c<�h�8
�=��L�X��=�Ȅ<��ؽ��w>���:-���{�=�3����VM=,r>�״;�J�PO�PՒ=�y�=>r ��&�ce`=��=*id=��g�2љ�e�=���D>�P�t���k;R�W=D/=z�b��伭��= �<� >Wo�=��t;Xl�9� ��qK#>éX��M�OTK�$��89�=j��=�!a��y�����=O�=���;�c�,a>KSP�W_�=��o=�i=C1I��q��M3>��;=
�=Y˽$�3>Ι�=��@�:M�=h>�}���8���2=�z�I�0<A��=���;R,༑��<\��==�F=�c�����=}*��V���=�[��>�V>^�^�=
�<O��R�1>d|�=�����H�=.��<�=lY�<�>[R-<)C���T�=�2���^�:��==�稽�Ln����S^�=������<�5i�yH>Y!�Jp�=�X�<������>�I�<qv)=�4t��\}=����G>.��<C���]��=k�8<���<R+>�B�;A�����⼛[��K�=hL>_��=�\��3 =���=JPJ���ܽ0�,���9;W=��L=OK��̙�Q\�;hO�=޷7�غx=�A�<I��=�8_=b�:L��=9�y=/�b=�=��<?��=��`�r�z=k��UK�&=>��=f���6 =�u	���Q=
=��%*ƼQ��<�b=�w�=D�b=�����M�,H��T�9>�SD�,&=4u�=�>���<��.�oX8��`�;+<Nʔ���=,j<Θ;<w�=-Ɗ<D4��H<=����=��<ji�=M��<S` ��^�	���A�j�>�{�b'm����<�;<�"�<��p=��f�1	1>=���V���LP<��ʽ�oZ<{W�_��=�`@<����%�THX<�D>��%=�����N�	>�u�=����b��½�p>hs�;ǁp��z�x#v=)J<�J��c��Fcg=|ED=w��<�^)��X�<��=y���G��v?�5�Z];���=v��m�(>��<����1?)>�F��&�=��ƽ��0=�{>��{=��n�X	��>��q�>P%,�jr�=ߎ=���<8�?�ز$�LhF����=�J)>�� >�Y�<�������=M�����v>z�@=\>)>�2̽��>��=Rg���W�i�	�u!���=F�}�����T�в�=o{�=XC��9��Q�W=���Q���Ӷ<c+�e9�<R�$=��7�h���o��@���Ǽ���ia$�ю�=Q9�,JԺ�4��v��Tn~�����A�̽TH�6�/=�����<4Dk=�j�=��!=��S=��ŽXҐ��4;}ۍ=��==5�<��5�ԩ�=_2��XЄ<���=h��E�=B������r-�=�	��Q��í�<Z��#"m�/s�m	�b+�<���}�'>$��=!�ܽm��<��c<�Z<��3�=�1��r=h>=&VT����=>T;��=�G!��'��^=�H��d	�8�=�ּI�=�̈=��ҽ8����K��:=Jwz=u�P���=�<�`[=�=��=��=�Zh=R�<o3#>�-��=y�<�v�<e�=
2�==��<A,=Q�"=�[�=��=��[Y�(�
�9Ƥ��,	�ɑ�=/F����=.4y=���=����ʀ=8l���|�X]>���=LE-���wb�<4���ٷ���@=�=\��9�����>�3���U��=�v�=��$���W��u�={��=T6
>�`�9��=�h= �l=ҡ����=��;'8ȼ��ɼl6	�a��c�\=��= �+�~�=���\oW;��<��>	Ӭ���=�Dr=aeJ=l9�<(?>�>� g�9�=�$�=t��<���绁��f���X�Cnd=�3����[=�v%�o�'�����3=q�1<���:�7�fO�&�$�>ɪ<�^��5�=�h���,B0>,>���=������N����=H��=e�ֺ��C���G�<=$�=��4�pt=��=����=M^�<8 ��[>�ۼ�fǽщ�=	�9>��[�#<������R1��Į�)��=}��={�L����QM�6�ü��;��X�=[$�kH�ےL�N�<�ݑ��Oj=�a<�<��F���=��D>���t>=���l\��8O=�ض=���-�����/>\(i�~����F=e���[�(��8=\ ༘�=8˦�rG�y� =@F>�C�=���R:�������H;q1 �Z"K�Z+׼栏=��=c�<�%���<}��������������N���z&>���=1�?=V˶=��E=�>׽�ࣽ��h��V=�&"F=��=G�Ժ��<;�)=C�`�_�g<N����D�9U�;�� ��7<	����$C>wy��jy�=�q�<H����i=+�8�}�<�չ;�q����'��T��3�=U�e=���=CV����=�����K�m{��/�j=�^*� ��m�}�AK�=�G�<L"(>c
�z?=�Mw����G�!=s�R�Q5>�(�<#=Ǹ�=�\���Eܼ˲��Fϼ�6�������=̹����y<B�e�����ԅ<���<���ܕ�=��=0$p=A�>��C�	>�Խ�g�<hd;�\=�~^��a=��B �3۽���=ɭP�ڞ�<�	ܻ`=���2>Z̽}w/=0����C���<|Z�|#�*�����I�L�=kg�t홽��I=Ѿ�=�=�ʜ<|�y�`.�;��)����%��<�0ʽ�!9>�و=���*��=v�@=�彷V==��`���=�_h�I��p,潉�O<J{=�+�=����� ��N>t�<T]�=&{�;��n��)w<7l$=hu�/� =���<+��=G	>N|�K��=�ّ�S�K>!��4}`�C�
>g�9<�'��A4k>$>y=ӽ�e�=�(���z3;c�=�]
��ߕ=j��<�t����m<ׁ�;ng���H�=d��jr=��;��Y��Ƚ�'�=�>�46��<�;�3]=9��=�)���z=1����N;y���L8>�q���=�|����=�n<�����ν	V�=�ഽ��m>O����b=q1��d2y���<{�<y�=�@�=I	�W,o<3dv=��L�U�;��ͽ�,~=13="᜽���*�=��=C��OD_�!_�<����4��&=ŝ�;tf:�F�>�QŻvXɽ���Xhs���{;��L�^݉���[�-�O=��f=px=����l��=��+<ܣ�<��[����=қN���>��=�v���1���nܽ`x�=~=�a��_dc=��=ro�5�̽gk=-}<��w�v(���{a�K��=�ʾ�\�ս�-T>�����|����$=P�=!)�<	jx=0�=��<���=�^�;�I�=���=�(0<�柽3ݼ�4@<�n�=w�����Tp�^!���
>��U<6���/�=��<�hļC��>D����ǽ���=�7=&O�+���1��=gF��u={�X;!��=��ҽ
7���Ҟ=Kj�=�z�=f��� G<�O=�=�<0����M=�=X=�i�=���=���=B]�=�،��Y��ͱ<�z���?�=y6�=f��[o=�c:��>�=�}0>�w��R��T��������K��Y�<8�<%3���c����~�K�ս[Ek<�0�=T��<&!ɽ��	;%��=or�<[��;$}���j������$>1�<jF	=�|<��=�ǼUi=ǰl����+��n�ԽKd�=a�v���=-�=��缷��=��;8�3>�K=�G�<p����N�=R�&����������=֮�X��<l/;� g=���=&LY����=t��Z��q��<�.>�):�}׽�>�bH���=���=	2�&볻�ѽ��+>����Lɽ4K;�:tH7����=r�"��M8�l��=�為�f�<H"�EQ޼��S=�L�@P�=_jƽ�4�qכ<T,>ʧ=��iuQ�^.���=��=���=W��?#�;�E=���=�=�;��م�=F<F���7��H����=oO3=,5�<棏��E�9KV�����%>�"�=BȽ�脽 �]�g�>��">g�a���>��=?-S���;�P#��m
>j@�=^>�=�о=��=�C�8'z#>Δ>4����DV�vr�����������b>�����^y�ɧ�;�"�|�<4�<J+r�\�1>,Vn�Z好Ι�?�q�'T
>LZC>#S�KC�=T෽.��=�����=�0ϼ�֨�P�>��Q;~�>X{�<�+�<�s���\���B�=��M�b&>2gq=z�P=�XT=�풼�V�;l�
=���/`!=��=���=� <pT�������>Ü�=z�<���<UC�=��=�;�=�>�=��ӻÏ�=j��=�u�e'�<�z��0�;s���8�H12=����ͅ=�v=���=��={o�,t=Ŏ-=2�	=�Xf��s�����O�='��{��=�	��:o�=(������=�����O|���f\���<��=�V=��T��`>���Gqѽ,�F>�>�N�cYڼ !�����Sܽd��<�X��NF=}�ݽne���v=͔���a�p��t��=d� =%l=��9;>/��F���A��Ss�<�O��D	>\>�H�=�u�=oQ=��6���$���=Z�o���ν�T�;]�==��8�u=/>�mk��<�A<�6<ӵ��ݹ�����/�/��NA;�~<��=w�2�%B��k���wh�fc</�=�5_d��<�}>轍���F"�|^F���8�ǻ�j��mي=�bH��9�=VM˽�S^�~�+�l�&��삽���=�3���>d��u=Q���T��S{=����o���[A���(��%�=K�d��|/�r�;>$>���<_*<~�;i��=$��=�3�=�󘽜�=�Y
=~���s���U�w=����.;h���n��=ỻ< �=j4K�q�������xe=�:�=m����ʚ=ԩ�������O�:����J� >��;�J��=��L=�)�<�V=����;���<�J1��ǻM�Z��80=`B�=l��*pc��̕<O��=r����<We�=-e<�2���Fμ���=r�Ƚ~ls�[����ǽgLp�%Of=½����Y�^%��4.�a�=�o�S��@�<���<�J���Cw;������=fѽ�y�_�=<c�=��z�0�_=V=�a���{սd@�=��/����=�Ţ=p�(>���<8U�>\ؼ�лo����9�j&w=�;!޲�>>q=�=�AM=�:��`�m��>Pm��=�/=��=�=��=[�<�<�=Y����=5�<[�����<�p𽉙l���(�f��=���]���܊�=�᧽|c�=�F�;nQ=�i(=��V�� �=Ű�K'���/=p��<�6�
ĽV�/�ox<�X�=zw6=m��=_��=��$=��m���q�R��<�~��[&���軮�����a<=����=rzʽ?4�=N���<��~�P=j��=��O���(~=l�s<I�<HN꽍�m=8>yļaG�=jl�����#���Ǖ=1��̓=�D���*�o�7��"�ׯ[��ҽ̘�<�<��=L����Bٻ��?=� Z�-�9�1���<�����	���n���j�<L�T=���b� ���	��=����m�����=��>\��=^{=��>�g�=>�:� F�r�X�r��=���<H�*�=�s��I>�õ<�&�=Hd��,$�:�E�wG��&�Ú�;���<�p��G>�׽����I��槨���*�� �=��y](=�K��u���߼����� ���.>u�м� >�ŭ<��>w����P��F	l=f�=wI"��1��0=��\	>�՗���=��˽.�D��JK��⼽�;(;)@�=I�
>�~�=㈺=�����u�<�]���߃�ݻ�Q�������u�aAڽ0�r:�@��rѽ#o�=��d���<i�>s;
�Vk�<�>{��=2倽땽��μX�<�n���������<a{�����<�S���~=�
���Ũ��\��)<����3�ʩ�=I�w>%��uK�=.�>��=�U����=�f==Nx=ם=%��=�a >ސc=�����E�<hڼn7�F_�����=���<E���ta=���y������=Ԕ��b�f�p'������n8=��<AL�{a�=�>w�>��؀��1�<UE>�4=9�B�tм:�	�M 
=�����=s��<L��<"�=�.^=N/F<��ƻ�5�=�=�V�=fS��}�>!�q<�6�<W߼��_���=i�8=h�=���d�X=�a��+���Ž�,=��>+��<�y���=���S���ͻ�=�=�L0��d=�F��V�.��=��<��_=)�&�"�<��{���=�+Y\=m�U>�za����T�=�V����<��+=\M�8I{<eU~=^4+���=�4H� �B��3��̃=�<�;�=�W0<��c�[�鼌Ͻ�<Bڢ��"=���\��(���=�g�;�:B�jU�=yXT=�{�=�-���3��1�1mw=��uV�cV=$'�<�{���-ڼU!&��r�=�sD�/D��$d=��w*Ѽʨ��'��˽�<f>��=�'=θ =
��<��:�ᘽO1��|�;)�=c&g=C�Q���~����<�wf�C��k�5��@׼��~���">.n�=��ֽ�ſ�N>�\��S���=sG�=F>�}<Ջ8� k�bxq�V,t=TZJ=V�����]�:+ "�Qð=(d5�)w>@�!��I��������5�N�=��䩨����=wF����e��Õ�Ax�=��k��L>��<֏>#�Q�)��=�0��4�=	>�=����=(�t==Jݽ���	�4=">�[�=7�ؽ�V<<m �<lL�>�D%>�{������J��?�=��%���<��V=��޻&;��-�>}9�=���<pPc>�k���.$>i�<��4;��`=�*�{'2=�����r<����0\=�e>�@伦�W>���==+=�57>ýet���9�N��Fu�<��
�N�`���(���z�J�B>��ܻ���<��=P�:�93�k�w�����~�/��~���?�C��<]	�<8�~���=�*_���>Ѓ��� �T]�=S�D<�5�=m ڽ3�l�=2?"<�D��fԽ���=fFD�=]�����;�1�����=�U����N4c<�{^���=+筼%=Q<��:��-X����<�'=9���U��<�.��z}+����<���='�1�D�(=yJ=��5=��*f�=y�	>�Tн��ѽ� ���˽��m=��<���=+�=u�>Z�z{:�y��P~<1)>�d4<	�=N�ͽ�<Z�,=P2:���<�c��34ܽ�D�=XG�)@�����W��<J�a<`J�=��(;i�S��<`��c��<�����=�]�=��K=�U=�:�=�9���uh�o$����=?h9<�����<nƵ���=�)ۻ�9�(7t�_?�;�ە='���q�=^�u=$��D��b=T��<�>8�=��킽v/��i�L���>��l=z�Ľ�#��ND��!�%í=3��N�;�jn�>"=�
�=}�;�w	�)_%�u�<şd=�q�z����dw<����e=�&=���P>/AK=�m��s:�]9�<L:R�t�R=�8=�A"�2Vռ,ļ~3{=�0>Q82�ڃ뽀6��M,�����ʝ=�	(>�_�qa=�t�=LXƼ�R=�r�������=��E���f=��5=�e����2=M�=V4�=?i�����=r�A=�_�=(�����=�-(>!���Z��XBŽ07�ro�<ɘ��̆��(ǽ�����M<yn0=��=[l/=JƧ������C��Zu��	�=?�=�a3�rE�<N��iv�=��m<f�e�7���{<��<&����aE<\��=����]��_�{��<{P���F&=�~�3Ĕ<3Aǽ�%��cl"=t/3�M�o=$; �����o�>�p�:���:v�/)ϻ0�I<&=D��aʽ�U>�(ּ��
��녽�<x�E;ֿ*�#����8�<�\>:�ʼ��f��P�=���=�]:<�>��>� p=��=a)�<�U==�=�0��0M�<v�O��ˢ�mE�=�ع<��>�雺<�k��[��0����M<���%�=Q����ɼ�J��m	.>���<��̼p��,�$��ܮ<�	>h�>6�i=�����=T��H���!�2=83<�R+��E�<YK=Gk=���<������ >�8E>�؈����=��;�=R��<�I=4J,�;\#=Ȓ����;X�����E��;5�P��=�%���;=N8�<O��@g�=�D�Oݢ�ד�<9��=��=�)g�]yϼ�F��/Q<�7==�l<�>�}��/�(>L��<�$�=�@��02��&��=��I��* �<f�=��=%�l��G=�����a	�,>�^�=Ҵ�=	����a=�$��xw=�I=H�Z=z�>���=��Mի=�nv���.��W �����b>ҷX=��@=���=6�ѽ���=@?�<5��{ڼ%>�i�<EB+=g6=��-�8O"���=�K�=!V߽;�H��;1�+<��`=�=L�h=G�v����M��膢=�
I�"���=��<���"<&���O=H�B��	��]pb=�Ͳ����k�u=$�y��A$��a�=SMֽ`��<~(L�2��=T؞�`�T����=�B2��΅;R1=@7]=���=R�7�沓���s��=a�=�%=�|ܽ����&N���˽���=(Ef�>��T��=Z��}�O>0�B=�Y=�*��<?aA��jQ=Mq�=��1>LX=`��=�_�=𫏽i�=螺=B&��!}=`�H<4� >��;M�ֽ����=&=�)>�?b=,Ľ�����0�=l�ҽ/K��Uߨ=�b��Q�=�<t ���_a�j웽��=J'�"����X>�fD=W�=Z��<���=8E��r��V����G���������1\���@��}�c=_���o#=�OѼ���i4>!E��T�����f�S;P�E���r�<��=�Ǧ�}6�<���=�IQ�v�<;�5=��>�]�=�-�r���A*<%��[���1A=!(�<���=��\=����=�e=��<n� �|���m��	> =����i<@�!��>�\��gެ�-B���-=k�=�-���>��ݽpJսţ�_
��7�<:�T�P�=*��<LX=J�O=����e�=�u��`�=�湽�q=�$�<����V[�_B�=�P>ؿI;��=�r�=b��=9��=諔=��<�	��� 2�1a$>�b=�����*�@ɽ���<]/��M��<9��=���=?��=�z;
ݼf2E�NT�;2ʽ�]=���=��=���=����3>t�]���=��g��[�=���>�bg�z���� �7f�Y�0഼>�=�O<��QJg=P�s�`S��� >@����BS=}-��(<�~��2���B;<u������˵��:�<���>�$<�T�=(Ǽ�����0>x��6��[>�5:�^��=���v��v=����<��c<�=bI=nD><����&��c�<���W��=�v��e�+=��W�i��=�j�=�~:���7=K3��X�I��"��\��N =B[�=��<b�9S{�=b�J�!AȽ��[=�����2>��ؼ�>�= ��<5_�=)��<�j�;�I]=���=i�<AO>P���,	6=p��=~�=��ļ�Ȁ>�qb�?U=ҿd=��Ż;���_ٽ����~=ي�Z���ʽ���À�J��=J8������'���5�P
�v��/<N�>�/�='�<��M��1�=m5f=�2�<����YT�ͷؽM�T=��&<sL=�S=�Uٽ�~�+5�=��<S�:�#�L=�/=nZսR��<Q�м�p*����=���h���16=�=|����BK��vK��ˑ��ᤩ=����?���p"=o�ݽ`��7�i�=�!n�<x%���ܱ�T6|<�)��:=��<�9�=�݇�Er����<�0>m�<��F����%v���=��q��v �C��v�+=��=@�����<[�P��������;��K����`=���3�=&�=�p�=ξ��S0��[{�7�̼Nj�={b&=J}y�$�����<�&���v="J;ݣ�<���Rt�?|<�9�=f��<�{μo���=��=`R�C�佭�<{�-=��;Y{=Z��:��=(ME�TG(>X��=�B-=S�=����|�[����叽Q	�=ݳ�<�ȋ=G��;T����/=fr��a<	 �/.�=�ŏ��-U>�A<y�;���=�A0���2��bk漲o)� r��3ь=S&���Z=�v��.��=2Ua;L��;��<⚽=�,=f�i����gt�2JP=�=����E���8>=�*{�w�=�w�<���<���=�h�m>�﮼嶚=�?2�pI���7x��W���Ӽ�^ ����>�=�/Z;�7=%�=�&���܇;"xD�JLɽ���=��Y=0�/�z���ʸ�=�ɽ7��=�� <'��
��a�=� �<���=	�km->ڏ�ӹ����"�Q̈́=��D=�%�zs=�8��>X��<X"0�K~��$V��٪F��<$]�:��G��,M=���<%۹<��:��=����kP,��<�=R�>��H=g
/�7-��=-(��T���$��7QR<����@��J�<д���_S�4A��VD;MS���{��ʽCd=���=w�*�V�Z�\��=1�H���<�P�
��"���C�%�]�>L��<��w�Zk�<�3��Ⱥ=�H��^��F�=�X�����h9��-������Kn���p<M�Ӽ�>�?�=>7ȼ�S߽��=*,�<��ǻ���Iz�=A��֤�U��<��=���l��f��=��p��q0=�;g�c��7!�>=0�=�^�>^��=
�N����=��=��<���	�O�A#z=�亩��;��m< J,�˓<�uP�yP=�:����RU�<bʞ�<*���C*�{6>�S>~4���z�<Pr�����K�<�V�� �<��=MM2=� h<Z�߽���<l�=Fη���#:��7�Z ,>3�(��������������=�B�= ��<�z=��3=?��=��=�Ͻ桋��}��=v'�=$����m<�_<_F�0���� �L�~>I���7��}ɓ=�Q>�`>��H<���=�����=�	�=@�9�=M�$%ݽ���=�.#�Å�!M�=48=�=�~=p����>�����v����d=�],<�+)�辋���=Q轙��;=S�=Һ
=cE<a�g��t=����fb��).��Z����>>y!��Ձ�h�=�����>Y��<	�>�ὁ�=��=����=L9����=�������
p=�+_� ��b1�==CG���9|{�~^��k�m=i�ּS�������=�ʨ;�X���8����u��=������JR���b�ʷ�=C�;M-��R)�s��; /�!L�x��=��B=���="@t=����6:ݼ�Ž�Ռ����=ɧ漿��= �+<�^�=-־���%���}=D%��j>��)���`��d#�Y8�/^U�3�=��s���c=�rT�!��=�M%>-ѥ���O=@�`=��=�� ���A=W�D��3��5z����=Ŋ6<��������?���6����>�Z^�H�=���=���H� �*�=ڔ�<�U>4Ι���ɽ���<Y'>�Ƽ�}�=(_��U�ݽ'/�<�tc=�Do�[|����.������p>/R>����`=&��=�i���wn�=��m���<�|�=�L�=��W�k�]I<��6�Cs�=���;�x����ŽҐ=0���������=�PM�Puy;��9=�a��1-�v��;k9=��=��<:�&;º����<^�<�=��>eE%���m=��==���6Ԯ<��f��=t�V=�
̽�˽�����Z��Q0=��>�=Y�B�C��=0�,����<���!�!�G�<<z�A����{�һu�K;Z�3�6��k����&�<���=�B�p�1�>r{��;�2�D�"=!5�=�j���\�=�0f=!#�=H��=Ot�<Éz<hQx=M۽IF7��Ks=��K<A�<��f=�㑽��i�t'[�Jm�^�5<�>/)�=���=M��<��=& �=�:�=�HL��D�=�j�=��-�Ru�� �=���==S=�-�=��=�0`<�0�=ݝ#���=dZ��Q@Ὁ��_�M=��>�b�=G�����<��4�t��==�=�a���3�n�ü��=O�<IR�<_j��n��=�7'>CwȽ����k�#<;
 >-�Hk=��y�Yr`��.�<��i=�=�=7�<qFo�>�=��ʽ��x=!A1=م���">lk�<
W �!I���R<)�>ޚ�=x?�<g��=��=�>��<j���Qޭ��9��,=x[8�h���tE<�1��8�r���0;���G��=���꘹���2=)�R=���=�1�=�00�ʄ�vѳ�9��<�2%���ӽ4��<���/��=�[�<Ds=m#����;͡�=C2�=3�N��/�j7��tE�3��<&��ť=7p��I�T���I�,��x ���!�Q��<�.�}����{�����Mּ�-��=���I�g�}��𔽧�>9�2�s��S!9��zN>�⏼��=a� �@��=��~�;��=���=��?��ɑ��-�=1h�18>���Ӭ�&M��P>�'�=�ǎ=��D��_�=���=6�=W��S�=]hI�Dɽ��̽.�L=#�>yݽ�~�K��=��=�(
��	&=k`F<��=5Ւ<7 >�'��z�>�jc��ґ= ���|L�ڝ�<u�Ի&�e=�������=G��=�ե�GC7������[=ILG�${��-:>S��=�'�����=�����k����E��]�<�G彬>½:<Q�q�:ث=0c=.+q<,�M=��L<g�>�M=�ǽ9"E=]��ɝ�j#O��Y�=%��R�=�
�����8>;Pּ�Z�d������{<{����<zi�r�=wg��
l�=�_C=}�>5���7\=i޹��ľ�v)��x�5��Dռ���=�����=�$F=��;��+4=$�j=�4��[��<�h�=wr���޼oC���z��<V<�a ��#7��jR=w��<~<��;<�'����R=h��i�A<N��sA��>�;�=r�1�SV(=���;�=I�=h�ݽ]k8�� >��:���*�I���>��!<Y�<L��<q�R>b�2=Ly=�F��U:tCּ�\9�=5;=;H����'=�M�<�-���1󼥧�=��N;�v8�b�=��¼�N�h�=S���Dt���9����=�p��R��=Gߋ���0���*��0ˊ<�	�=�~�� ���"u��}�<�AO��|���ֽ�Q=vZ�<�ߞ���ɽ{!y<-彶aɽѷ>Խ��b=�aZ=/:�A04>=�;�EZ>�C�=@9s=�s<��?�����㞼]L�<!�@=�&��͞<�r=HO������E�8=�</=���%k�s�#���=eR�|=������Gf�j��<r������e���3A��l)=KS�;+m�=�=0��<�7�z&=�/���t����ӽ~������P���yԽ���	耽3EK�k�!=$�=�j�=���;��!>r㛽&���-����Y=���;�Z4>i�:<�n�<e^�=�-�?���+���(�B�S=Am�ܕ)=��<`{u�� E>�Gb�^N�=�~8�2�c���>�[6��}��ꧽ�g=>��x����4=�/�ۂ�=D_�;��ýDH�;��)<�-|=��;��=�ͼ޷ɽƼC��I�=��<S�i=>�#��>�M�%��iϼ��'�Q��D�=uYݼ<t��M�<=�<�v¼�j&�
#=^��=���z<z��=�%��/����<��<ZUY:V�&=F!��\�=j��t=2��<�ԕ�A��=O��%�<nx�<�?�i1p��[�|�=��=�b���뽽Ě4=G�<�^�N����;�4�=̏�=�D�=x��w�νH�(=U�=3�����<;�=q#s��u3��^>���=�1�<.�4�2�b�U�;��;�Vƽ �W<A��;_�=� !�'���o�Ƚlc�=R�˼�>�G�ᬽJ<:>=�I=���<I(E>r9?�BԪ����=I>�9==�=))��&<%m0>.�+<������;�8E�]�����	��tʸ<'j�bE�=ـ=�G�=(�߽������m�:=ٖ@=}Vؼ�y���d�<�j >�Y���N�<6��Ʉc=���<�9�<h��=����~�T<i�=���=a���X�=a%>�{ƽُ�;��=�Q>K���L����R{<�t�=vP�=��=�������0�F�/>W�^=q�M=����c�=|^�=�ʽՇ�=bWu=��=�j�%��;w�\=�E��2��;T����<n�A��>�?~�cĽ�z���s>&;�ߌ��<�Q�=ב�=9�9�M=�#���!/>�=]X<.�=Q�л��4>"J�=�K�=Վ7����=u�<|��<4ax��>뷌=�\P=R<[�<=��&<PB=ײ�=�!�9a�;lQ�<2ʁ��,>����{t�=Xo0>�����I>aA<.�=�.�֭�=�|���( �=��>߲�=�� =$�2�2�>W��=�9�;�޽�
=�=�?>�;揋<�Ո�ʦ��K0ý��=8��<�'�����G���?��Ӌ�3使���@� >4��<^�����/o~�-�=+�ʽ�C���	=ҡ�<ꗽwA��<�j>�7�=/�H��������=�EG=Xg=t�<�4�=���i��<�g�=%�W=���2�����=�@��9=�0A�ζ =4��A��=Gf�=aZ��u|���%,�gtG�T[(<3�<�	׽�;=v���	Q�>��XX>ђ7���U�#�>���:�\*!=��P=ӰH����MG�<p�c�p; ��T�F�xd�M��<���~�<�7ü�T]��H�=���h��=����;�Q=pJ�s�=��b�K.�=9+�=�|�=���=�k�=-N_=a���f�Ľ�Q0=�̘=y�4=З�x��=`��<ʋ4<���=�֘<�ߊ=1+7�J�
��>#P�����<wp;K����<��<�q8��=彆�x�Ɔ6;�l�=��<���9,�>D�#�� 輔��<Hg=sk=5kмw�0�V���\��� ��=��=��<�{��vWc=C"���=�M>�g�;6P�=v㤽��I=z��a&�=�]�<����Et=h4彪A�ETǽ�#��[u=f�<=t+�Dd�cs>��-=���=�!=��&�1<����%>x*�=
\�,"�;{;<؛F>M���|B�\g=<��=j8�<� =�z�� Z9���h�"�RW�9��?�8�=�N=�<��a�Jjd=���<mɸ��;=�L�{*��"�!�8Ὄ��z=_��=�*!>7�8=�}e=�+>E�=H	�=
��=Z������oY=�d�k<�=�N����>�Ə=O&[>L�=��$=����>�4>:�=��꽋��=J�"�hz�<d�O�X\<A�<f؏=���S	�4���N<8Ib��}�#�����=�j)��xx=�#ƽ��6=)�=�L�<k�;+$�ptA� 4�>rf��MA���C>#�%���k=
z���Ku<����>�ܥ=\I�Z���)w;^ԽPg}�����_�>
!j�������=6�,��+���=2��/s{<���0½��X�mk���.�<�X�<ձ��A\���<<���;;Pֽ�r�=�d!>4�ͼ�ϼ�_�b�_<պ���晽R�=r�<�Z�����˳s�w�=ч���	��Q���v��4�|���<,f`=��<�ϰ<�4ǽ�o��7�<�v�	?Q�v�}<�:������O=�C�=SX=��y�E�&=(׽��u�˹�=o����&��}=�f>d�==�����<j�h<t�#='LF<�5�<T����2>��~=�K��ả=J�g="���K��<a����=����""�<r ý���;����=�LB�n�#X��ӎ����=�T&>?[ɼ���|�>�4=ߴ��;n�=h���ל��-ﻬ�$��1S��M��!߼u�ļSŲ�_�r�$�׼
<�g=�(�=Ρ����<,�۽����b��%%>�1�=�@x���%��I=�H&�u�:p~=���	�=�2�3:p�Gk�H�"7Լ�	�����^�=�^
����r�<"�	���<>��'=�%H<_u;���Ϸ/�� �=��=�m�;m9=���1�.�4�=;�E>���=7Y����<o@�=C<F���X�ʓG��W=��>��ϼ\�l<O��=p��<���c!���B�h=���=v�����=�_�<\����1����T=sY��K7	>��>���ܼz�=��Ժ�-���=��*�lq#>`����ļ[ֱ=+\�~M���>�̜��2�<�_:fz���!B<���=� H�`�>�>�q-��n=BG�:�>��U�ƽy9=�׉<Ĳ�=c���{U���=�65>��8��ļX}<�>�}�;<j�`��a 5��7�N&�=��==����	�=�}=��<�����J�Z>}����K��̢���ֻW��h�=q]�=]_=�-_��|���й[üM'+<�M~;_��=0��=P�b<rV�u2�=.P����&=+�#>pc.�ã�<�D��1����{��_ �yc��]�<<S�=�P��E�=� ��[��3���{@����������>��Q��
>m]�=vD�<����ps���KȽ�T�=J(�=и	����<g۰=|��ֵ�<2<!�-=�����<�Х��v��ߊ�<7��<�Ȋ���W;)J��G�
�5*6<R�Ͻ"�J��E�:,S`=/��h�=rx5=vv=���N�;=&�4<N}>ё�<cļ��=�6b�e��#!�;���=J��m=�y=Xܪ�1�-<JUy�~|>yG����P>3��=hz���Ȼ��4���Z>�ؽ�&2�㎲=nt����=0�G��R�=��W�j=�����#4k=�ҽ��7�ֱ�<B�)�3u$���=�q=z�����=6�=���=9lf��4�=ϙ�<�s���`2=xN�=��<���+��y��<Q*9=��a=-�=��;(�_=��S=h.i��_�=�H����D=ܬ�;A����d���J=!�u��V�<J�˽���+����.����Cչ=@�ڼ�h�<]>�z<X}�������\<إʽy%�=M���%�p=�\�=�F�DrB=:���/�=���=�bf��	��@�z=����h��=��>l�;�唢������ =��=��\=�կ=��=뙼�+$�����u�=K$���ּ��=����T���l۽�(�Qʞ�9y��Ƽޚ����>D�">��<�e�<���;:d�� >�J<�m(��Ի�Ƚѝ�>�!�o�~<܋�T"��?�[<�9&>��=n�ػ̩�=�Ý<�Tx<��\�\H�=-�Z��@�=0���� ��̪=L�N����<�[��_�=+�<��=������=^�=iQw=�[�ZN���1��Մ�+?����d�[����<� :=JBQ�0۽B��=O��5P�<(��=M!��}��c1�^���)�=�v�=+��<n�`�*=��!�=��[��K8�.
l<?#z>��M<�M���/K�/��=&�7={��<��|=q�|;Ĺ!�:�2��=P�=��=������$R�<�qȽ�B5=�.=�S4�;3����J��<ω=�b̽�<![�<��)�v��;��=��B��=Bi�<�,G<t��;�Y]�'�@�X/�<,<P�F<��L�2�<i�=��-��r���<���xs>���=�iv���]��'1=���=ԟ��⭗����=�Q�=���4�<��!����=��=Y��;�73����;�������=v�=�㔼�h�;ٞ=��4N� 1�~�<�h=JY=�R#=��S�h=v)�ƿ�=0/���C�, �=Hn��W�7=<�;Q�<$��=��C;ڦ������=Bn�<�@%>C�O=5C��OҼ��=p���P{ļ���=7Y/=�;p��( ����=5�<�{��=�K��	�=nx�=Wi��ɵ�uJ�����8(��E_=2�Z��SH�����U=�Т��^��!�G�YݽŞ�=��y<$��I)��+�+�'�>�߅;�ev=븁�!�
>ݫ�=-=o5<|�N����=�^��y�ν�.�=ꗢ��#�;4ھ�	�@�ϕ>b��=��<���<x�f=25Խ�ν�>�I>7��9$H=R�t�HSP<=L��i�������o��:�:��<�o7=/</">xS�=
z�=�^^�g�G�gP;�����p ��3Q�W�=��a��	̽!_��p�<���=� �ʟ�=�$����(>���=E%=M��<���1x���p<s���x&�;����Xv���9=�Jo<򌶽G5=�}>�Nӻ(�g�ybG=�3��Ӝ�=�
�=���<pz �$C><�����=Ҭ����<g
���=o�u���<Ǝc=C�w�>��ƽ��"�K�k���>n}O=��=G+>�`d�y_���6<��Ȼ�s��=���=�@����0=�T#='EQ=*�򽂹罵����ֽ�>���=,�=��	>U<��*>Q:ȼ��'< ��Q�O=�T<H\+�s�u�cX�=@�={�����=����k��X�л�ӽ�H>-ھ�a���<,.>ҷ�=��߬�@�=�f�=����,Լnq�����~����)�j��=��;�e8�|4=����	/�=�Ժ�{<��=O��=�]o=�<p~����<;��=]�#�N�S<�y�=A_�ȱ�=?��i*F>�,=o�����=�:>9���y�=+�ӽʯ�=�3g=Z|�=*ɡ<�BT���r��7��& a=|��;��=�.:7()�~ ���	�|��c� �-�=L���n=n�(����ޢB���������_�<L@ȼ���=@ģ�^1ͽ�� �W�iM3>�w=>��=�l�;�\=�j�+0�=��=�mQ=�j=:�x��HKe<D�O���=�#��ʧ>��;'8=������\>�����f����8���$�=��=M��S�<�@��R5��X� =�?���=�Bf=G�#<��������սմ��/-R�K��V_���o�DM>&��#k>=[ّ>�ýё�=�%=Ph�kQ�;����݆��9K>�=��T�01N=��3;�p<d���t��C
"��3��DEټ"ҁ=dX=�Ȉ�G���NA����o=�"=�������u��<>[s�QX��~<�<�]>�%e=R,R��q�R��3>��0��H�=�����ｆ�5��=&�:�ci��Vv�]�ýGf7���<���;�>�<�<ǉ����5�S$8���8��|���=��>	r�=dz$>2��!�F=�}�:�՟�I�/�ȳ<�2q>S���B�=��<V%�$�>1.�=�B{��º<#��=���&v>�h=Oֽ�wb�?�=H+��m���$,��x>b���QU*=�G->�����Ի�S3=L���_o<T��<��=|���h�=����>5=10�<��ʽ �I8�;����=�|>Àü�<2�\��R��T�=?\��&�v<�����>��<N��=�����ý�~�O��="-]�v�4��<����0���|=�1����<t��<0:�;�k*=0��<gu���ݼ�Җ=��Ͻ�)���N�=^G=)��=� >2j�<=�-�+Ɖ���=�>������������#�K��=Х<��=�闽�K��c�WMh���=ҿL�ŉ�0*��.	�<��f�U@�� ,=r����Ң=`��;�ļʅ�=��[=9�=s��ˋ=p��=,/*<R�� ܑ����<�u�����\#4= 
��e�w<*�;=�R�:�ƭ�y;7=[�>Ob�=ʷ�=��<��������������^�$��8>���_����H;�>��
��1�@[�ybU�/V�=���t3�+_<�酽0�>�@��l�S�����*�T��)��1�� [��
N=52=�L[���=�c���u�=�����P��2�����/^�<��W�o���iL>B�=MR!��}&�){���z>P�/�D�%���`=��M���`�����S�a�+��);=,��D,������5=�����׼��>��v�������a��Ζ�;F0���y�<�g�=�[+��d�<vD�<�D��ؖ���=q����Ľ��=2>��H>q�)>���p$�=ɳ�=v�=n��΅3>8h�F��*?��Ń=6C���=�7��&����#�� ������o�,���;���=�W=�f<��*�5�>� �=[L����y=�uC=%�;>c�;F�=ݫ�33�V�$�� �;H�Y���߽�Z�=�-��4;�N!�:���ʽ�����������<�=@�>9�λ��-�H^>�Eӻ���=Y�F=m�=o2l<�[�< �F>�K+���>����z�=�@�<&���!?��v=š���Ä����QB��
e�=h޽jo����<[<z��<��=��K���<:;�=%oM=��1����:cFA=�� �����=�;�=WS��%P=��=k��<��E=,�=t��=�����=`� >��7=�s<<3��v���^����=���=d��=���<Ŝ�����K��.�5=�(�=�f+=�40=ٓ��3��<Ec�;�
4�ME����=䰏=p%>�A��)a�懼Ұ���޽�!1m�8�d=��=|�'=*���e�=w#E=6�=q����<��M>��H<�m��ܒ=���=�=��$�=�A����B+<�=:=D}ڽ<���H>��] �5�;��/�vS��y+=����Cn�������1��f�=��H��=�"T�������;�\�����Է��9���<-P&9��=K�=��R-��|=�D<��=�� =Cɻǜ���B�ƭ2����c(�ěX����W+#>IӉ�Qld�l�i=�Tͽ,-[�^��)���
)=���<Nv��'G�SjC=��><�U=��=�u�=*
F����{m�=\ۼx�=+����*>�XD���[<�o=M}u= �x=�U#��/5�@�<6�R>,S�=��n=���V�r�Mg=�)�����
<�<�T>(�ͽVsP<�*;n3��/��=.'��?����=�n�=A�=�p��W<�����;�I�=��`=�*�-Y]�E��=�d�����r�G����=�J�=���;V�� ���{'��FM�[��=(g��=A�i�f�{)�����p�<�s=û	=�'�3��;�=��<�O��cl�>Z��0��e�P����������:�t~=�l=�� >�`X:n��Gׯ;%�[�9]�=�v�=�ܗ=꜆�ܙq���g��9�=[e����>��$>g�;;$Ͻ���r=��;U&)��-�=���Z�ﭫ>O&��н��>z=�\��1����=)�>	۽�g�=�n�3E[���= �S=Dl��^���*U��H]=��=%�=��F�q���=��=��H����L >摼m�*���#=|�<M綠tE�;��ԺxY�r�>ʤ���.���ʔ=i�����>s�>�
�v��p��;M"4=�B����Ҽ_~h��>�=�-�<O@�0�$>
��^�=�?�=�l0=ZpD=r5����=�3�=Ñ���'�����=�0׽��}<����H���+>��ƽ�Q;U�|=S���0=j�=c�.�j� �<���h=wQ�=gK޼
=�=Y�B�O��^����N=��ټ-��S�=�P2�!7+�1��>󷖽e��k6�=!��<��6<�X;=�7>�ޏ�ڣ���>�_�6=>!-��N>'��=��>ӿ=���;�L�����?�����=�,����!>5�Ɗ��ꎂ�d�=H]1�yԱ=�O�����D�=�k<Q�:"�k=2cJ���=���*x�=-Ͻ�2�w=�6I=���e����#�����T���꼿�=�����۰=;쿽�4�<4p�=�L�<�iὡu�<<S>C=��j=�6�=^ý����1�=�=i�e=�׽9�bT纂NH=��n�z=�E���>�D��=���P�<py+>�j3;�Gm�D��n;�=�Fw���G��D&=�`y=\F�=��>=�y%�!߆�y�L>��.>�T�<n9�%�.>XsB�+Ba=�eM=��L��
���o>�<���T��i=�>t���a���.��l=�����|=��6�;>���=_eb������>��<��=x�,<`�;� =�s�=-?f=�v>"*�H >t��=k���,�<5��f�̽iRc�E�=����35���������ٵ��S��7F=��H>&�=����ŋ�q�>�X ���#���ý�ý}䰽�f�s٪�ګ�=�YӽN�<�b�٪�<)�;�L̻=ß>�w�=�#�=#��Q}�=|�@=��=zb�����:�[>I9�{?���:껆��=8�F�aw-��a��-���V�=9��vk�d׭�����Be=��;�>лb����<k �=�Ƚ�X佞�Ļn���|���%)�=*�q=����ͼ���Fs�=t�?<xf�8*��\Ę;����j�<���7�<&W��;�4��e��Z?�=�����uu<󶣽c�=ݚ|=��Z�=���L���KE>oL��y��<�;Ȃ����M�vAE<��=�h�p r;��<f�;\9�<\Z�=�ཆ`��������=�=�����;vV�=�1�&�x=�/�<�/��&���.�=����<�D½kX>��r=v�W���>��=r���/��'��w���.ѽ��=�-»A�
>���j=$=�C�=4�<���=�
3=�u��߇=8;<>w/>7 6=�ک��SA=��=��<�ψ��H���"����=�e��.���<v��z����ڼ�M%�^;��шF;�,<<L���M����<�kE�;:�g�������ؚ=���<8������s���V�����w=����ĸμ��[=�0��9��:mS`=���;�8I�^Tڼ��^Y��)x�IV�=���!���o��2>�/=z��=ޜq�=<q�k��=y�����<:�=��u=	GG�x�i=�=�<���=n5��oܽ4Uн�{P=?��=������-@=q �l�w�;����=�{�<dq�=>��m=����M�:�m8
����=Q�)=�M=I_>=��Qhۼǝ�=����M�;��-��%9�Z&>_+�=���>B7���x�=�=���e8e�;f�=�"��0r��H�=�Vn�ܲ=C9<��ܥm=;��,�F��9��=��ȽU�!�����_<�	!=]���;�=Һ���=���<��O����+w�bK��k�=LL�=�[�<�-�=��=?�D��@o=�]L=�e2��̕�E�=��>�b�v�:��S�Bz	��yU��Қ=$ �<+���5��)�<��.����=���� ~=�K��^F�<rG=w�B�2��=�c��M��=&��< =|�<���=|�����:<�v���G=��7<c�=^���`����Y�
��������+�=pLڼ�ն�uGE=j2=��=H�<?��)7�<�(�=��ݽ�;�=�kK��.c=��!=�<`O�<#�ڽxB�:4g�=��>Jj�7i��[����<@��=��r==���F���`(���<=�!z=�"�
K�=9#�@+Ѽ�>�L9��螼(T.����K��=޻<<��=�x��=���<��=� N=z/�=1=����p��/��VA������u���b>"C<:��<p���H����������� ��'�E�:ķ�<a�=����-�=�E>�6"���e==�R�ǹ�e��<�i�����Fu�b7�<򉅼?0m=��`��Zû��0�\ ���<Wyۼ.L��a;���C���=bm��ױ��h1�N����D�����=����ޘ���]�" ��o.>,ۜ=���=�k��ѼT�=yđ=C(߽�����F����-<�˽�N�=�'�=܆=��=&��X��=��=�.��8�����u��=�N�=���<9��=��ڼW�U<��_���B�B�;�s�L��;���5>+���F=��)<�=�U�=o~�"{�T��Ex�<g��=s��`���J�j�L��=zT���B_�=o�#�4�<3��<u��hq��"ٽ�,v��9�<��=�88�Kb���c�=z<�j�=��q�X�w;��>��ڽp��(���+���-"��醼G�ӽ�'#����9?��<�H�=�H�e��<�r��6�=N�9�X�u=�j=p;d�=GI��L=뫵�t����tX0�Q�｜|>+�˽�MڽS�<���]��=�����;�� =�1����G=$߻ɺ��Fi�=�ʏ=H��=�JG=<Hʽ��ļ�Ż����,T��>~����>���=��_�D�=�x�ϋ)��B=�t����=��Z=��->4��<Qc5�����<���<&��=n��=�.¼u뎽��B��̼=��/�R���4<�6S=H�3=?�m=�z�?�缁�=L!>7n�;��==C	>3vO��<1]	=Eݽ!�G��k�Q=>�X�<f0�<��o�)��=�.R�
�8��k�=�W��k�k<i+�<yW�^v���E=��&�?�"=:�����-�������1���ϼ$D��{��X��TY����<a���q"���=D5b=ע�d<�����>R#���4�5��=�J�=|<���<�A0:}��c=#��;�&��_|>��ɼE]̼����4@>D6�����<����쿽Y2>�
����Ἐ�=z�|����Ch�=I�_�7���If<��;͐Ƚ*�-=@eH<u����޽�bQ�S���΂<���� );7KĻ/&�=��,>�5K��v����=fV3<H���A��->e=}�<���=�ӕ���+�<p�a�Cq/<�f�=\P�Z�<�e]�=RT<�<
=�v�=is���_�=R��=qp�:P���?=��">|�=e;�;i�4�!�ƽ+E=��=����J�=����yS�z�;��{�A"�;���{{=��=�]k����R'�=��[>�c�=���u�Լ�E~�a�=��=.����>Xݐ<"�3Ay<��o��=1�����2<�:�;9�<����1輾�
>�Q=���;ot�����<r[^>lD�=�䜽�㚼����<��9�+y>�q=�k�����ଅ���=~�ʽ����{����̽����G�O�5=�"��lI<��9���g=1a�� 2û�3�=�	>�E�=�B��콠h5����=�`�=�(|��B9< ��<�#z�QM=��<,ҽ4F�=��<�I4������k=;ߣ�7�{�^2��H=��f>���=��=�兽۴@����</�c����:��=��ҽT\��>��uj���<]d��v��<��C=���F��K="%K��J4�'v��?�½���:�6-���;a�f>}�B��<�Q�=�v]�bdh�B�R=B˼~�@���ٽ��=8��H�<!㽻X�=F~<I9����3�1>��fu5<��&�=�߈�=A=&z9=^{Ž���=n�	=���	�<������ｏ��<y�Q=���<L�QF�<�[�- 7�;;>t*����=��߼3պ��E�<3�">�1�=L�v<y ��e�x�Ƚ�Y�=͙�����yȼ�=�2H��r�o\��x��=��S�W�%���A=�[��i��| W;���w�>	�Y����<�!<m!n<#���W,�=�Iƽϗa��<M��2�<�o����=�U=p]��*K����=BP>�c>����؆�=��ͼ���Xн�=`t�G�d�HƘ�0>���<C��6�>��T9�Ҽ�Aͽ�4ռ�>��K�=<����x+�x�
=>q���*<���=_c�=���=W,�<��<�Nн�P���ȑ��dd=�ڽ�S:<&�z=�_A�7�3��q�<fݚ���!��*���A���89q�*>I�P���2��a����d��`S���>�=�f=���?�=7�e��xƼt/�<�����K��z��4�6�!1�������}�K���x���hYV<W�2�0�˼)������?��`���T�Z>}���Ķ<It?����,�=
�~z����	���;��]�xa4��ɽ���=]�h�5�W�xn�-�<s³;�	<U`=���=[��@�Ž�%<�=��d�ɛ�=��= �Ǽ�C��E��=~��=�ά�/��F��=����uv�{��=�3#�tt�=��q�,=���O�=�/G�%�ƽ�[�<�i=�f�=z�.�ioG=R=��,�5��=FV>�f��ƅ�=�9�K���w���;�����U�>��>�)F=D���y]=d��|$E�ٵ�=�mf�ļ=��l<���9М<)�ý�j׺UF>u�:?ʰ=)���o���k=yJ��:��">F�J��>=ӭ�="P���.-�9s�<b8=z�W=�Y�=�4�����<|&�<J�=6|���<�����N�?=7e^=u�=:�"=[E
�f����]>=�p	�ݛ�=3��<�#�P>X�">���<&X=����K$�=q=�?�*��������_o=��G=,�>m����<>F>�=_!����>�*�=k�O=W�`�=������ʽ�5 >-9?�Sbл�&�4%]=�9�*д���(�OX�[���\�=�/����S��U���o�<���������P۽���=�8���)���>��X��ju��颻�ȣ=�SJ>�]q����<��=+�:=;ѽ�= ^�=�I�=�����<��>�aw�����Q=��=H>x<����O��:*k�:�=��<Do8=A.>>b� =��<�?x���=ehh=�P��n�=�	h�����~G߼y����g=��8>,҂=x�>�\<��>�~i=^=bZ��#��<�)�=f4`�ʬ�=a�D>�ڻ/�\����+Un=���o�<�}&:�T#���,|=�#�=�����?
��#D�:��<�%�<&��f!<�A���50=?�8>�� >�pt=��>���[�=��<��⼻���N2>��%���g=	Z߽��¼�!��Z;E��lG�m��=��!�5�>�n�=L���\�G�"�
�-�i=s5_�t�=�F�<��ٽV��=�E>D����j<�����f���w��+�=�M�*Q�<5��=�J'>��<�o�=p��=9��=�"὾+½�;<v����=0.+=�﷽��X�����A>½�&O=�b�q�=+~>+�=��sռg;��H����=�5<Z���>�����'��.�@c&�5�#��u�=�u�<�Y�=D�A�@���V8׽�̽�S���Y=��Ӽ`\>+���/�=��w=��2=X��=�璽-�/���">��X�קȽ�������d���f�k�WV��޸~�UB�I��<r�4���Z��7�����된�<���>�	�g�9=�q��� <��=&3ݽ;9�<�=�Y��"Ĥ��,~=�;�=�xH=d�4=�� ��A��륞=�=�N�=0��P��rh�<�7�;���<���=���=5��=��K=RA����:�w�=�n4�"\�<�A;��\���>|�I�i�=�Q�|=+�],>�7h<�����;Q�0��=D˻�d�=jU=F�+y�;kI�<�8�]���;?<�:ν��<�����\=22=�T�=|nN=
�{=u�����=�w�=��=�½X�����%`=�,s��z>�p%>|��0�=������<l7 >Ƈ��gP=�.>sٽ�xܽ#�+�k6��(�@���<�A�=.z$��F�O�==��=�+��]<z'=���޼њ�=t��<ߝ�=��E��q������~7��c�<���=�T�=_q��m�</�s=|=K=�?���ٽ »�w��VJ>[{��J����q0<��X�=����~��={f�=�O���= F��9�=�s��X=a����B�=�>X�E���F�=j6`;EΞ�ʿ���¼cK�<OL0�S�L>�:�?I!�%������������.U=~�=�gE��C=�׼T�<Av���6=�C��Vk(��a�=�X!>�Ǽ�i=K�3�F3�<��=\�<�!&<�;=����)�=*����Λ�����m����!�9Ĝ�=
R̽�FS�FnS��^E=Y����>=ͫE=���<Λ=53�<��(���E>�(�=�Žmۂ<-���s���@>���<��<~
D�tY=�p��4�=��Ǽ���<u5����<��ѽ�]�?�����	=�ʞ;�᭽��w>��+<d�G=^�f�h4��C�=~`g=�틽#�>�U�����'R���@�D�ɼQ�|����=��U=h���j�=�D�=����=�n½�>��=�r=�b�8�t=����]\���W��{e=�~��tم=��=�V�E��<�6W�b��{�<����G�P�_U�=��t=o¾�=iB�P3�=�=o0=���;OX:�?$<'�=�� �����o�=�'G=�N�<&`	����y�<?�<ܣ��� »�)=����`�=4�1��õ�S�h=�����	�r�;6�=6/t�.���u�<_J4��J�E�h=1�<�=>�~<���$>��<�,��G��|� =K��#T�=&{}B��f;���w�<oʹ<��j���)�!��=+�=��.= y���1�V�<4]�=��9�vO��U�<q)���
��da��i�����=� �J��k^�7�*>0g���=�# =!�=��
�N���h{�=p�=lyؽ���<l�<�����<��2=֙A��U��>�=�/ؽ�Ԛ<���<�:�=�..�h�C=�H��^�����aҚ=�Y
���,�T5�����`�<� �<;g�=�x�=o�<5fF=��=a�_�3=.̰<yR=W�=a�ȼMp�<��L�r�=��m=	]�=��=�.�=#=��*=++���=��}�ڔ�<g>H�B���g<��=Ⱥ�=��
�հ�<�^R���P=�d�<��S����<�+��>�=z�b=�P��b$���p>J�<D�ƽ�Ի8)�E�N�z�ٽ\�׽�_-��|���&i=�r�=^�ӽw���9�R�>�a<�c��� �����i�5����E=je>:����M=2�/��w��#>�ҽ�I<=3�Q>�=�B)>� �9a���r�;�Ѽ�VS�l�X=�/��ۏ5���%=���=� ƽ�z�=����ۢ=m��<��@=9E�h罶nּk%��)�=�~�<s�l=�;̽ ː<Z�T�
Hc�ɏ=�%J���t��/ ���?>�=�vm;@v�=�>Q�P��|����=^�s<��(=��=�;�P��=k�>4�^=�I��~	>�ī���=����������*U�;eS=2`�-� =�'���m��Hs�<�ޢ�+ ��.7�<�wɻ��k��xμ�O�4��dcX��F4���)�iS >�L�=�e>g"���:�=�8L=��;�y���'�=��nGo=���`����	���m��*�=U��#%���9��������u��i�ٽw>g���͘���<s�>�V���:J�'��=Kː��V�=!5�<ӣa=Z<�8=4���6>�O3���껈ȗ=.ӽmꗽ�>�=���9^\���H�����| �`�]:�-e<e�̽���=��<Ħ-��Ͻ�
=���=���<�dm>d�~����U<���m������Qvg�r��<�H�=�;�>[�W$�=K���h�&�$4��ds<��ؽ�M�=�4�6Z<��/��R6�:R<1*��(;��=]��<���y��~���b&>*� = �m= =���<i9��+�=}���&=t�<M��m�=�%�=�x�<v J<<oh���5��ߢ���"��rU=��ҽf�c>��=��=����=B/�=��>�ko=��=�}i=Jv=�^�i��@F<x��=98e��E�=�/ɽO	����=H >��=^7'��J�=����D�;�_5���=�?n=����8=��=E��=%���Yˀ�AqE=]��<�)&>p��<�����Ǽ�~ɽA�]�Z&�=�=�Vk=��ؽ^��=�ƽ�@>�!`O�T��=\~���`��7>�� =�cŽQv�=�i={��=ʝ>1{;;{K��<�<�2>U 9�=��U<''�>���=���*v���8��!͓;H�=�ͽ�2&>�'s��;>���<�!=��*=%/������DS>Ĝ�<Tw�׋�@�=¯D��P!��> =S���p���!��$��􎽺L�=�FL>2�bD�=��s��d>
>b��;�Z����=2�>��4�� ��`N���;>
����wW�u�H=z��<�e�<���=RC �Kd=3�	�=��=v@�<@~@>�Mc=�S�FB޽ZM�<d��=#���h��X��<��0�Ӌ�<7��<>�W;4�=[n�=\��<l+4>���=[&=���<��=�;���">��ʽe��:&j�=G�<����y��<k�߼���=�
Z<��/�P�,�f�<���Q��<p=	|��P6<�`��7�۽����`p<����މ=#P���ν[͔<%�R=�BH���=%�$��4��)ϼ�yؕ�~⼞��;���=^�r<�U�=q1� u�p:��䍽��^���>5Q>��<V�s=���={�b������=s_<�����꼿��=#�
��Eƽsu�<�ѹ�5�὘q6�>_[=�ȟ�ಅ=�oQ���L��6̽�9���X�=����?>X�<�a���h�<AOB�e	�=�����(��2�<�눽��Ӽ��g=��]<,(��w=��	=@`�=��=�M�������ɔ=����c$>��{=�ב<5�謪=J��=��@=�����=��= b��kM�y9=���W`>׃�=��=�M�=�<Ǽ�%=�Ӻ���ý
�<���2ߐ=彙��=բ��yԼ0�1=�����6=cv=�]/=S��T`�=_��=��7<�r���4{�2��=��>a������=o�<6�ٽ�0��<P@�=u���h�=mQf��B�/R'��)�x�Q=W�=߯	��{��qY�eBY=�^��C�*�Z��<7�^<4޻=�:1>%C̼f½���<��ν+:�_�	=���E�=dX�*�C=�}�4�.��GӽxW9*��<xH>ur=�d=+b�=n��ډ���~�D^�=�JV;�/�:�>�?����=���>%m(�>���}U>�ۣ�,3�=Fn�8]��;�>�6��_�f=ڎ�=ށ缴�����<��=h�4<;�=��<�X�+���lqM=%�r=!�<-ȱ=<��=��=CA�<""��D%F=ϭ����R>���<M�L�]�Z���<��z=��/<��>�,5�zI��^���X*F=�m�=u���:�!>v�=`�׽���=*"����,L����=���7?�=�z��\>��Y�;I�=ȣ�=Vٽ�)�<.V�K� >p{s�ȡ��ziW�E�A=���7��̺>U�Q�/�������i�=�� =ʀ������N�|W;�ȃ<�ٽ_Z��G���U<OD=���<s:ټ Y|=X�c=!��;"��=�.���g�}F=�~F��E>��.>���C->����=�	Ƽ H�=n�=��5=�f�D������]+�<�����,s=�0
�1x����N��W>�]$������6�ɩ=>���ʧ����黺=�S%>�ȹ<��3>��f�.�]=>����<x�<�u1=f�ʼX>�>=�s\�^�~=%��<� ������������T�B��=I������=�Kt�&��&��z�����`"����=)I��%>O��Y|�|'G�rZڽf�4>�ť���#=�jH�5(\=&)=Y�r<��<��W�<��=R��=!�=8M<��D��;0O<�=+�ݻѼ�<��I>6���G�����A۽�箼7���hؼ�.,�im	�a�y<��<Wƚ���=w^�U.�=������=q;t<5��=ę�Ii]=)N,>��=���0~�=##��:���Y��h�=!�=r�=^�<���=<�E=f�~�џ=Fg�NU�WΛ=Q�>=OZ�<Jզ<w�g�KD��lM�<eZ�=�C���\�W�+>vٰ=�<�E��;=δ<����=�5�=����=23����>��ٽ�_�͇L=ß��XX�=�#�#�$���4��^��&=" ټ����m߻��n���<ݢ �5[:���<4�Iz=���Dq�=��>~��u�4�S�����)��=���� ������z��g(=멖��h�<�ȼ��Y=��ҽ���{��=�p	>X�μ �>��˼]T���U�=�'=|�b��wi=�>>Gr�=-J�<����������|!!>���=}:_>K�
���h�+�A�j>���A輫��:���<���t�=J�!����=�g�<C�
=�p�=�?��A3�=��=�1��==-�>U&b=~x���V�����<�<�<�/�<���*��=2���]8���G������>��q�?O5<��:=Ԍ�=��0��>�<�)=�.�G���b̼."�=��>�=��)>fb��`мFh�=�T��!	=�����p�����='>����O=,x�<����pfû��=���=y�9�=/V���B=�.����<X�>[��<ڕ�=���;$�Y�g������
��3�l��6�/����ݐ=�ڂ��ED=/\��^����&��j�1n(��d�=V�>��=[�=�=�a�_�6�S�=ŭ=�<%���=�ٖ�[��<
�=u
� �4�ϼ}aP��R�=�{����;�T[��R��>>�/�O���^n�<QN*�V�޽�V�=`ٽ=<��o����~	<W��<�MG=Cu>��E��(>)����@�<�J��(����=	���1�==��>�`ߜ<��=#?�=���=Y˽I	>�SZ�7�н����k���=�']=ɺm�j�꽕_=����*K=�p�=e�=R�=�=:o���g����=�N�=��$>۷.=]R�!�;$�%�< U�I{���;��ݽ�=~2�����='ȼ����c�<��=����|㷽�ܺ�͡=z�R�*})<H|>O�Hk�9���jL�� Ƚ��>�ÄE��>�{�;�$>m���S�5=jw�=��3��@A���5;F.�=@>�UJ�<M�=���'7>�=�jF<^��^Y'>O����=�rK�<q�=ދ���<7���\>'��2=W���y
>'�=��M=62���rڽ\��M'@����_�S=�+ ��Cݽי�����=g����= �=�P	>���=�<)ѽ_��<�����ɻ�>��9�,nm<+��<8x&=YT=���;�e���RT<�|=�$½����?�n<K��=wP<?K�ϩ<'�<G�/>�b��V-k<��>w�8=�,��I�=b���g�=4��=.�z�����]���&].>���EQ<�M;=1D�=Ά4=s =���b=U�=�d>�墽�Z�:ƀ<҃�s󆽈|��h��B�����c��#=���=�М�X%=k��=�#�y*���.I���V���<���:<%<Dv���2P=�f=,\���>$�ջO[U=z����>���=�е=�=�H=t��K�=�L*��=�m��W\B��n<_'�=���8�=O��Ğm<���شo<���=�d=�w~<.�ڽF���\�<�J�=:�<�.����2�?�u���۽��>��:��Ｌ���D}->��'�SP���Ԍ��o6�t�k����=3�˽���<"��<ܪ½lW�����<o7�=Aȼ>_=�^�=|Z������G>��=0` �Ӊ��=��j<���=���<��<�}���{����Ũ<��I=���=�_>�K <��=�i�=qX
�4`h=*���E1�������9">�O�<˒����O=I;�<�گ=Z��<q�R��%ѽl��<^)`�1y'>�P�<���=�G�-�׼|<B�TA�;�����E�=J������=~�=C6>6�ͽ�s<pD��������;(v`=a(O>j�P���=�윽�������9oCܽ8�νR<�=�}�K�>d��.]�c���Q?;�=�
�<����� ��]N*>����}��uy�=r�>�X;)W�=���욼�^;L�<@�;B����=�-��lp2>'(-� ��M&�� l��z>d&1>i�o�|:��\?��p;줽��1��=K�O���=���=���]\�=��)<�&�`ﹽ�錽�g=4�=����M)���I<rm�=�F<:�[��|�=1r=^�j�$��=]� �o�m�#Uz�Ճ =���-kc<�=j>>��<-o��<�=�Y<��=���j��<_�_��=�B�=v#T=��=�6���'!=H��<��*f=Q����W���䳽�Q=�16;%̃<�%�<,�=#Cнx޼�����d�=���=nʽ8��=C�@�X��|+�g������<e7���E{=�!�=��<�;�=�白�;#�0�<k��*8̽v���1�=e�v=���=����.=޽��=���=X:��B<�g��<��~����=#D�����ܷ&����Ɣ�4�>�,G<�\[=š0�ԥG��M�
�=u��<P�?=l����=�н�>=c%5��; =z���E��:i�(��;vO⽻�:��2�=�MO=Zo�Z�=
��:��<~�j<_�=�o=w��:�u�=����@�b�Q�l��<0N =�-=V%�=�j�=�
O>�B=X~[=��o�U��=P��<7��5q��c���>�R��6|p<ט����=�����d�=��O����=^c=�a�:u�;��'>�h�=�콬$���S]�Gm��� Q=���<���l=�b�=�a���D��Ľvpk;k�\������=_��<�>佺z	=$�����w���7>�u¹���=C(}�0S��j����:�����$�]�%����fD=�X=�ٽ��� �6��<�=�<�=>������|�ϻ������[�;���=l�=w�k�g�O=��R=�>	>���<���n��[�H>T'T=ee�
ɽI8q>m0%>Co���	>g��<� �=�(���h�^;>���=P��(����;Z>����z����==>,=���<ԍp<y=�(�=AU/�K"=�н�W۽>�<$m>z��=%�>���F�O="�=žL��PE>�A1>�j��@�=�4;���j<�+�=�д��#<��Y�eV��*�=C�w�
�CM����s=�'������k�=ڔ�V~�i��=�����>�����F2;&�=��ͽ��>�#��Z�T�� =�b���P5=T=�<L�=8|ǽ�%�=�T�x[=�F��bB=>>�5>߰�=�(K=�}=z��=�2�<�d�=��'��=0`w��@�j�����W=0���̐��*�87�=�Y=��=�>�xBL� �=���<
����<�+��LJ�K'�=�d���ٽõ���+=I��g�뻭�=�ş9�]��<���gB<��=�A�=-�[��M>��K>7$����
��!�=⹰����=C=��<O�Q=����*C�=!�3���1=wM2�f���Ց=X<%~��WTc<-O�=�>G{��X��".��8{=�U�=���!bZ�K���X[��ώ=8����
�=�����ک<t�e���Խr�<`�=W��=[��;��p=�_�:@ �=)�
���=�-��&�j=�;5=���
��"<W�8<��z<��0�rl��Nڽ�
=6�0=}Q���>d}���e�<��K=Y;�=����"x>���������u	>�񽤱Ҽ��!O=j��='= 7F=~ =rO�;�(�<��&>.�><��<8_�@�4=��J=�I�`{�<�39=R/=�9�=��;�\�=�n��ܜ�=�F�'�����=�������}=T�1��}�X���=�4m����=WC������wQ���{����<3q�i�=�ؒ=�Ϯ=���4�N;�Ys;��h=�����sǽ�}�=`�<˝�26<�ҷ=�F<���6`�+4�����<�%���=d`>�#���=,�����=�WS= �#��=�h#>z�]�G���[����<%�ܽ�u�]!�=�l=�鼈�=�� =~�=��y��Z�=��N<��*<T=@!m;��<�=��{=Z�����=�7�:�����	>�>�M&�4_F����W����-ɽ-jU=����,��_�<7�ٽ�w��ⅽ���0x�30�UO����7=��T�{>S����=����Tp�_��=�;�=�<g=L�v<`��H<�= ��=�㚼�X<Zaͼ?��|�߽\�*�9��+�Z��V"=7>�#E��3�=��ֽԓ�=�j)=�=H5���ѼU��C�>��t=N�2�md�=��F=���=K)���TQ=t�Q�/<�>��uD���a�U��=�>�����oJ<�o<��<R�y=�`��;<J>��X�$R'=�㨽���<#�=Ha�=q�Z<����3�=�/꼭��<M��.�T� �!<=ƾ<�7�6}��<��:��K=%YT=�ic=��q��<��*����=Mr�= ן���b�u�=7[�$����U�']�<�*�<�>���<�@�=�=j�v<A���=�S���˽��B����<��>>��]�<���=��=j�==5����w�Bc㽴�J=;r�<3�q=�D�=t�O=�E�<울���=˥��N��pM����=��9=w��<�D�=�b�=�j��eJU=/N�=���<w�1�4j�<�n|����ѧ{�H>��S=/��;��=+�
=ks�;8��*DU=��*��M�='-���e�<�C<�'U=���=7g�g�;>�=� �=�>����P�<���{�-��j��B$d����=#��=����������L��9@�J�.<���:*<�}>֡���Fq���J��:x�
>���=I�=è=)���Z��=�����#��� >���=�������U=�2�=�&=��9���>���: �<
��󐢽�+=���R�$��5=rڦ��~ཁē�0�!=qW�<s��K�=�5��K�5>N>ؑ=�J=����T�;d����0��������2�������q�����<�O�=��ƽ�e�=cIB=�P�=�D����=s�1��.<>6�<�wfཅ������������==�@>�����n׼:�5<|Q�Q铽�=�F�,��b��-�=��^=b�����Mn�=|�,<n���=/4o�����,�\�� =9D<?��=c伎�D=�@ ���l�=��>=�k>��^��hw=�h���c�<<��m>�>.;�Q�ɓ=�	�<I�>�㼽ּ�d*=���<��ɽ��T�1x�=��=�s~=|#=5�<z�>C�ܼ�뵽%���j�-�[S~�k	\="�=v�q�B�w<U=c�h�0�?��W��F��S�+=󼃽^��[�[��嫽��=��w�k�+>�c���{� ~U=GVϼ1��=ۡ�<<�K�Wp�=�-O�A���ev�J'��x;�E��F=>��@�=����.��=z&�=�s�=��=1%�#G8���$�°�l�=����G�=>�=9j�<�=Qm�;�U�9��`ټ��p��v�n����<�S>To�=��� �Nz�H� =��=�1��[؀=Ԥ���0�>�
=�qw�	~���=jY1<��<��ӽ�5H���9=��<�݂���=�]��e�&=-Qw=��6�2Z�=9�˽�c��k>�D>�]=t��m�O�f��=H�=� {�L}�b)8>	8��ڏ�yw����b9��7>����`<V���-<�%��:�<2��=�=���=�U���s��͏<-��=<i�=O;�;�	��U����=#V<6��z߱=�/�g��=L��	E��Ü���%<
��<���=�2j=T��=ܒ���'>2��=$��c�%>>Q;7�<����E���۽�+-��w���<!	�=	(��F���5����<��<>������A�r�>=+L��ʱ�.��=���<��ҽ߽~���~=��i����=���>���:��f>�c*��t_������H�炙���q<��=��=+�}=�O>�Y�����=۫���&^=1�>ݗ�=���Y_=��!=���%������=Ԯ�;|�=waR����=��=��6<�Ŕ=��Z��X��
��� ���	� �{<�[�=�l��9jʼw��;s󡽼��~���J�ܽ�H=��v�6C;��6�<v$8�U��=�r�}���ּ�~�=��޽���T�%�<���۪�=$�=�}F�@�|<�g2��0D<Y�=���<�Y�����G���x[�-��-�G��{;�0V�+)����y����XV<~:����i�̼%�=➘�
��<�`�<�J=�Ҽ� >�$@���ǽ��=m<���ZF>���<��X��<��<�~ �+�2�����<R"z�W�c�D����<��<�y�P*;�8�=�ת=��:��=�l.>^�&=�랽��s��Ҽ]^�t�����=t}�=�؜=��'���W�)6@<��4>=�H=�,�=A��;}@0�l�����;y6�������<�=���=��j�,y�<l#�=���bO��ÿ�C�y=$pT�) ����<q6�1���	����L�]7=43->7��:2>�c�<�>��,�vt�=�Dּj�=��<�S���#�&v��穝���>��=�t���'A=~���(��{�A=�h>W1�#�0�=R���l��ߴ�=B/q<������=��=|��=�&b�u.��D�	����=t�(��=$
���{��o�=�������a�<H�<V�Լ^1>����=ǔn����;����1'½ǣ�bk�;�*��k�=�ԅ��w���>��⽕R��b��U��`�8=��-=�<)F<���=�A��A�=��>j�]�Aߓ=v�5���$=�73>X�ռ��=ĺ�i�(>�4'=�%�<�i
=���^�>E]��`��=�h��	��;H͵<k��R~S=���N	r<�#>��꽚��=\��<½ּq�����o�k�j�g<%P >���=��	=K� =u����4=%P�����=t>��A=w�ѼyE=���y�Q�M�n=�v���=�ȭ�m(�<3D�=%���P�>�U���=��Q-9=�׽m%ҽ�d�=3o����ȼ�٨<�vS=�b�9ɿF�Q�W�.:���U��|�=��=��5�,��6���"��2��=��1<��w�1�G�|_�cW4<Y���"��H�7��H��.�ŻD���2�<���r��=k��Ż��ȕ��.e�<~c-<�v�+�ԽI�C�0�<g#ּf.o������Ͻ1k��O�%<S��
B�-?=V�=��KF<2˛�N�=�Γ=�Ɨ�I(�;�᪽�>ӻ2�K��_�R������>�)>���� 
>�W�q���Q�����=[� >'���a]r�'b��d8:�r(���8�IؽYO="���^�=��н
 �:�V��A��)���=Ե����м%����=�R��ugڽ��
��Me��d�=pf�<�y�= Λ���s�|��;f'��-�'���H�<���;*=
��O���ܼ�{���B�����< C��p��<i��;�i����=n��=Y�=��$=������������;�!�<����)���d�6�y�:=ہ��`���N=#�Y=��|�b~%��1 >�E�=���~����=|[˽���	>ç�=V��=�T��	U��	J%;��==�y�w���.�=��v<e�że������.�h�G;��d=k �=����W�1$̽�J=�{C;u��y.�=�߼ W>����S���%�=������Z��;���[�S��k��H2�;Wf�<��=S�e>�x�Q�=�5{<d�i�&�;<��㽄,��
3�DK_=�Y3;��>�wb>V8��u����<z��=ĩ=E����7O=lh���=�F�<�k�=J�+c����麽��-����=���uU���J�=-�=�6�
�������3�9����;X��; ��������=s�ż}��\Kr=�ѣ�dc�=���=���<��¼}We�$�x�L �='�k�'� ��n��=⪮��&!�'�4;E{½�d@��}��UQ�;h���1>^^6=��3���<�������������I=�~�=4e��[�C<�#X� �v���=�]�=��=�]0�@����|�<�{߽%i$=U��b�`=a�(=������� X=k��	����Y>\�<�.<e�,<8セ���=�2S�^f�=ۙ7<ߊ��:<��d��F���XQ
����=30>���S�]��]=�*�:�y�<f6�<���=�c7>�5���>�s���ԝ����=J�G��T��&�=.Uɽ��;�-=a&�=�����p�<���Ґ@���#�4�t=H�ȼ(�ʽ��=�@����.�i�C8�=��<ʵ�=P-�=E��a�<js��cý{��=�4�~����=I�:�u�7<|{q��$���}����=]�;,R�=����@D��{;�=a��!5>=���=�p�=�:=[�O= 逼[�=%FG= q��]π��+ �鍽!]�<Δ�=�� �@��=x|l=�	��׻~Y�GJ�=ݍ�;�D�A� ��`"����B45<�%Ÿ{B=>�3�=� >?��=�Ҳ=ji�=k�.��"&����=8�=\�=�Kr<nZ=���;<�w=:o)=�0<[1������I�<.ǻ:�,]�����E�=�UH��#�=��G���=��x�a�W=4��=��	�ғ�=������<q��=E�;���k�=Fh�<2�G=��i=�Ĉ=z��=��=�	�=7���=�;/��28�j�z=�N�Q&�=��D>�&>џ�<�E<��=�q�r〻�΅��冼�낼D��c|ܻ����<y��Tޓ=X=_�
�D=X��=��U�D'�<ń=U�\=�����<J'>����=&>�����2<��H=<�>�<�:hA�<���=)��=VG�<$�=+��=�O^=�!�<�ٻe5���O(����=
��==&��{>��u�=4�7�����8�;/>ƣJ=]��P�<�=0��=��Z�{�!���ݙ!��f>"�޽M��="����[�u��5^�����,>����}'�=;�>"1o�j�м[����4��P�!=��=j��=S�n��<��=ݴx=�1L>`Ӵ��=0O�O*c=���<w��=N�=�Y�ކX=�%���"�<�Ȇ�8���������K=�(�������3�=�^�F������->�Խ��<��=��<��="��:�n�<)L9��}�=��N�-���$=�싽��~=:/�� �����b>; ��w�&#���2�O��A��CG<Sf�<c�B;ª=��$�μ��id��I�����<Ca^��N�Z�� �sH$=D�����׽�'���#޺z���հ�r'O���q���=��=�R�=%� =���=����/ӵ���H=�0����������,��K= �|��^=:Nһ��ӽD�Q��CI�^���I�->׎w�I>Lޯ=� '=�߻���a�l��팼�Y�<����n�^�.�=����7��~���Q�s��=~�`=�@�=�=?=*7��7�;lj�0��=�����jv��h�o���U���=6i���w<l4�꛷��d��3��49ٽ`�6�6�V=��=��൯���p=<1�m�x=���<ҧ�<)g�;4�%>j�Z=��-����=
`�<G{������'�<�}��Z�*�y��=��+��y=`����=ܗ�lɽ��
;�����=�#����<g�=)�U�O��<p�ʽ�[E�*��<\zK=��ὤ�U��u�<NS�;��=��N�ʴ�m�>�=ҽ�D=KC�B�{<"��~p���">Z�=Zk\<�@=}˽����.q�J����(=zm=@s��S���z�ܓ>"�>�e=*�U>@A�8m�Ľ�\��=�\.=j��/g���3_=(�,=��S=�
=4߂����<�$�< /=ML��A�<ҥ,=���;9�>p�Q=�<������p=��*��oV=\ۀ��=��A=���;�[��[��z�<���\<8V¼�ȼY�{=��;𣼻Ni�b_�=L�ƽӘ1=L�1=�k�=4���+�S=R��R��%݊�XE�r�B�f0>w�=2�=oO�;��<�H�=���<�e=���:�<�BL���;��/b�㝓=
$>�U�=�0>dZ=������<���l%<�=�岻jR߽@�	�ù>m�=�=��=2��x�O�+���l�8��=�Z=m�=�S�7"=�՞�ŏ���,�=��N�ף�����|�3<)�t=�� <�ֽ�t@=&��=��B=�O��l}�;�Ai�	,)=�Vٽn��<.��=��=�QB=��#>�$�<@l��t�9�.'�<��h= ���%枽���=��սx�^=�o<ۉ����V�n�A�U�˼�:�=�A��1ۻ�.�Ǽ�0�@��=י�=K�0�;���H����=h�;�O���8뽙�J��ӵ<��%�)�����[<�|	=� ���ye��E;�p$������+7<7Eg=�j	> �k=��<�f=u��;�a����=D����c;!~�<���=��=
\�1}%=m�=kr=9��=���=,b =GR7�%#M;�o�= �H>�1ཧ-�<�,)�����@i= ,=���<���<Q����7(�1�,>{O��ml�=��<?W=g�*>�J#�G�<�4!>괂=s�e� �<�:�<�`�=�P�=��<��λ�Ɇ=k�̽�G=+��=l��=��'>��=6�!��_�Ȕ�<<�%��#��^̽Z��;����Z��<�����=6ӽ�dҼ�b=Lz�<JN�=��齾hO�&/���Qļ��=Pv	� ?6���P��䗾��ܽt=̼��#�9�-;�����K< �_���.�n]S�;=�ؼ*{#=d�����0�q�^=u�w�uv�<�(ý��5�&�����=�ږ<aW�=\�M�p����-f=�->�Z=Ⰰ���=_B,��]�<>	=/�<���^;`�<i����$V����=Ǯ����>���^ü����k���&��k��IL���V��=v	�=~��<u��=���<�-�=x�>=��<��$�4���Uك<��V��k��=/~����=����->�;�:g�R�G�M]J���x<-����e=����K^>;I����=��E�������="��=�輽�����5=�(���-=�K9�G��=~>p���)=�j���&ӽ^���p���9>�),=�lL=�~9=��C=�ڛ=�->�;�޹���ڽq��#1��<	�B>�E�<�y<%-�T
���͎<:�<��_�^���ʼ�﻽,z�
4>��C�=0>a^׽�
��F+ ����;�F=D�2��v[<of��]yǽ�� �"��$�7{��<�1�=F��Ux��"-W�B��=S<|���	I=�*>' b�i}t=#�>kH=}�����T>��<��=��=�I�GF��S���u�$����=��=K7���Ԗ�����s�=�F�=����f��<�|+���<�� �($k��"�<Ռ��t켨uA��䄽h�<�P�=��$>�]Q�߂�=؂߼���"�9����==�j;�þ=��"����iں)X���MQ<R��=T��-,s=Br=eТ��4���%{���ͼ�Ӌ���=�?�<�ý�vl�`�=71=W�����������[��򐼹�'>3Ȍ�&T>0�=�Yp=�����">F��<�Z=�{<�œ�v�#��+=bB���/1>nr�<z��=�������[ ӽ��L��k&�%�+>�g�=͠׽�b��z�F�E�]=O+n� �Y< y=>GǼ��>�ݩ�iA���=~!������/=�e-=�y7<D+��#�<A�.�o+�<&2�_�=v%�=sS<�u��A;Z��<2m<0�<�[��.'=/Zz��`I=$q`<��ƽZy;=}Pu�Tf,=���=!����a�&��=�(��J�<-�k=�)>t=-=��x=Ŀ���ѽ�N<��;`ӻ��ѽ��=
���X��G�=L��=V��<��i�k�ݼB�9>=��<�`C=�~"�曀<���=��ؽ�����>N=��=�=:��<���=�����D_߽��=ad�<я����=���=8��<��~=-b����-}4;�k���,�g3�<�_��AR=�g!=�Z�=��缁l">А�Dk��>,<�P�<�Db�ځ/=%��=Ѽ��1��݋�= �N��y�Ӷ>���jǘ�lK�T�D����.����Q�=��4>Ju=U =�SĽ�	=�x[>��3�q�,=ȓϼ���i�=�
��ӿ���t=��=�\�<4o�<�r�=
Ω;L��=հ�=.j�=�e�:�U�<J��?�='.�<M�s��B׼-��=��<=ӻ����<>\Z�=�>�����֜<�F��C%>�u	�D̽�����ۗ�S�s�U	�<`� ��V
=GἼV�<���=�̫=�܋��3>80=�(�<�q4>������w��=��z�GQ%=FG�=.v-��|o� �X�L��:L`V=V�=rȌ�GCX=���<nf�w���u���=� ��f�<r{w=��<�=������<#ع�sV>&�>�����>|o[����*O�=Xo$=��
<�Ʈ=�Ώ��fX=g��=�)�=,����>�z˽�t���/=�]���U=M��=t.ؽ<L���>U��}��H<G�=�@=����)����>r�N=�S���L�=L?=���<K�=��{=!�=M��5�c�eTŽ �	���<�]�<z�>e��=��b��x�=o">��= D=��(>��=�;�W�ػis˽s�Z���$>8�<h�����<g�>=^AX�j��<ut��<U=b~���<�Έ�ʴ;��/U>�����i;�3��2ۼ��=2���î=�."<0
�<�lJ�����u�<9������<[m=���<��
=��=���=��)9�'����=Oa[�G<GÝ�H0��U���"����=��=�E�=7� ��[O>�,�=8T\=@f>ySӽ�E	>�B�<#��=�+�=		=�����Jн�=�����<z�ֽcx<Y�f<�ā=�'ʽZ$�=�A���Wl<Xf��o�=0=��=Y�����d<���yԷ=�ے=��<\��;1�u<);��� ����7���4�n�5�i�|N.=[�򻄄�<� +�(�M��_>XJw���潬�<=�3 ��i��7�>�c&=3�������ʏֻ[���(!=������<n��<C�=N��X\�;��D��|<_,�<��½g_+=����P�������&��O�b�r=��=֛�=
��<�"�T3���B�pe���;��� ��=db�}P=#�.��>��輊��=,m�<�þ�1�,��g;���ۀ�<��>=1Z����ݽ���=���=[a=^��=����E�=}�<t���;��X�A�B���-��<�ރ=�u=�P=���=�ł<6��ÿ�)J�<�V2���4�RG˽�,>T�+=�' �{��)�~�W>��/=���=눪���$<�Si=B��=Q�=�=óB�\��8_>��hMK>���<��o� [[:y�=ǆ����=[DG=K��٩�=ʇ6��w��x���5��g?��F>��s��M<�=u<�<N��5�#�d�>��=ֶ�=;�=1'����O����M��=��ߩ�= �C�󳛽�<T>�d�#��=[0��ӷ=0��=�ro�E(���N�=S��^R<�i��D�'��><>KkX�?8۽Y`+�ŵ���/>)󍽏������<>�=Gj�=�^>��=����(�=0��:�1�=n�[����<}>�=	R�<`_k�&�H�HN��*(��NO =+5���.=��=�{=�b�;�/a����=x��<l�<���c�>>�=�ޠ��)O>��u=�b���Q�;@�K<QAS�C��z�k���q��<v��,i=�< <*!��k⨽o�C�Y�lit�ܿ��dR��.�@=�"�9�<㚩<7Ϊ=�4V���=�4�=��Ľ��u������3>9%�wj�;1=����һ��<�R	>�=�[>��J�	��<U#��%��C2�������u=Ƃx=˫k����g0=?��=[>�x>�?�=ã�=rꔽ���}�����n��d<���6=�!��=z�s;,u���Yy�Otn����=ˣN=,{T=a>Լ8�k<��Z�I=:=�@�<���;|4\��vW=q�>]�ʼo��<�f�<��$�b��UA=�|ּ�82��X�=
��=�|�=�6�:&7��h-�=G­�퉧��V��E��=��>���;������/=)�����=�� =���<S�>S��n�E9�Џ;�ѭ��u@=%	y<�a*��2?=��Ǽ	pX�Ax�=�=�=�I=Ѕ�=aa=�lW��;I�*��˽�6�R�W����=����⚽B�>���<�&�=�f�j��X��=m��=@r�x=}=]��Js0=�4��=K)>F��=6�=���8�;��>|>�M9�/�=��5=���W��Ψ�=p��<G�%��&�9�=F��<�&����=t�q=uӿ=T/=�ך�e��=�;���m=f�=��0�k'�<g���,������dC�=)2>���=�*X=%(��D�EW�x
=��u<;X�<;j�
 z=�_l=_gս�e<��ed=X��El�<�#�=���y �=c> �]���>[a��l�R>�~���ɡ�R�<�.��&b�=� м;��=��A=ٿP�]!�=k�A�b �;U=4��&B;E��=���y^�_��=�˺>;]��=��S=�p��o�X�j�\�^�s������!�=�M:$�>����4��ڂb��_c<�"�Z�ڼ�Zм�X-��V��&�;k%�)	>�X�v�=f����%<����E��l�Y��%y��><w׼�����=��=թ�=�B��U��4=,�F��2H=�u�=�,�;9��m�$�~���e<�PG=������=9A�=��.��ɼ<~��=��o<E�u<N����|��Cp��(:X=SoN�5�����?<�`�&c�<�8��f��=5�>�k�;b����F���9=�Q
�I?<�=�=�����@��Q0���3��ak=֋2;zI�=��=Y�(���=:��f�?=���=d�����0�4=��*�E���(�;J�	�q�O>e�㽎,�����<f;�Pd=�`��H�=uN�;���=���<@�=v;H���<�߼=�SG=��&='��{�w�>��<cC�=���X>$����iM=�L>r�=��ڽ��=��=MXe<��������He<e8=��U=��Gh�����[h8 .�<3_�<�`=��=�3O=��ӽ�)>�C��=�ҽ�;j���ؼ,�g�ԏ�<��O�	��������P-G���b<�p|=���Ӱi=����|�<Ƈ�#P<μ�m���^`<�f�=h4<�"��=�=��Ľ��
>
w��r>^���z�=K٪�����lX>ᑩ�˘=�c��=��ƺ��=�s�����
�ۑ�=��q�R����>�	���[�����<��۽���b0�<$<�����aL>|�&�=Q��&�|=��F��ǒ�v=/	��ےX<���=[F���X�����=�ܼsPF=�=��d�W=�Jf=9��<Dk�o��<  �;K8���=Ƶ=�%i��&��� dL>�ټ�Le�=آ�=z�r=�'y>	Wн�>�=��=_����W�= ^��>r=����z��}=",��(>��=-Q(�C��<�=<ǩ�QH�����kw<oB��)Fh;g8�=Cp=�:���@=�����Fۼ(V���[=>�!=��9z=��&���Լ1<�=U�<�f����X>�4�<�O�;� �<,C	>��s1g�V�T>�*#��(�N���6=�d �#k=�����U����Q���=�:=mū�C��߆�:D�=��V�=T9���$<�S0�lc�=������c<�5-��2�=�E�>%�=Y��*x���:=`r�k\���m;�q�/4ǻ�K���c>�n<� �;B{=�nV<!j�<�V��s+=H��\�a�=f�'��JV=h��:�xd=��>�b!�\�=Q1�<�`�Ć�<?�d�=(�Y���%>�>���5Z=�윅�> >e�8�v�f��g��K��s�	�+������=��	����=�i��CX����	��>[=z��=P��;�a��l�>(@ּ�WͻH[�=\=�:;�����@<�����v�\�
=�kͽ�%�<j�y���=1���U��=Pi�0X"<�^��ϟ'��1������!�V����v�=�������=xv��R<&Q=������=Ѐ=h����{=hӗ��� >�'�0�<-�<=r#�=-@=���=��"��;�w�=��'���J=�r�����=�>J<M�K=��;�Ǽ�U�=�AƼN|�<MҼ�ץ�_��=�p�<���=�t=�&�=?t<�=�����	0=9����Տ���W=:�C=IG=�X�<5\=�
i���r=t��,���Rh���׽�>��{0>���< 1���\�o��?6>o��z��Ϣ=���>�3�|�=Mg�<P����:4=�"1=r ��~\=�-�}�=��b�-��%�91��;��=���e�vy]= ��@�S=�	�'��=:�=���;Rҵ��D=%~�<IX)�Ƽ
�A�r��>&=E(�ˑ��,��@�F<^B=�|~���>�G �4sI=\�xC>��K<��=�ٌ��?C�=�/�3a�v+�;."
�����P=���
�3���X�	R�=5p=�ѽ����� q=���=1��<l��k�<�4��b��=��l<c�
>wg���I);�f@�@b��kj�[j>8��<��>�,���C��o�>=����_�������=��.�&4<Ũ��^35�� ��:�����)���7<���=�B��
�I���pR7������\�=*P���;=_E8=C!�v>6�\=E49��E4���@�z������<��������<�����6.9��د���u=�瑽�w�<<�<
^=��M=�=E,�=Ц<��<>�����8P�<�1%<��˓>c�_>K�.����&+���J��Dc*>ws�=�'\��.��n�;�B�;�8V�݊���36�<L��=x�A��T�b�=��=�	�<3=�?�=���d�=��a�>
>��=|�*<�]2��u�=�e	�k�o�X�ƽkE9=)8=/��=j��������<�?�:j������*=^�*�I�ͽ�X�=�n��	=�>Q��<�=⽹�R=�#�<h��<��y�=��=�{�<��<v���h�=t.>B��=MQY����u"=�eO=��F�%���ҽռL���q��;\�0�<���=�ּ�=���ޑ=g�=�B�XK��~�=m�=4��]s=�������u=�3[�� X=b�Ƚ~�p��[Y�
`��G�:��:>�M������&�c�����*>%�<�۲=	Y�:�B=7D��7���n����U�<*ѽ-%��P`=�B�=V9�ބ,>��= l�;�2ݽFf��d�ѽ�٭��J=<O�rX�=q�x=%�����(�V^G=�&�;nL>-�=y$�=�S���=��3>����>V�=w������(dν��V<����Q��A�=�Ϸ�^��q3�;����z�����=���9�iX<K�=1G���"�=�E����+�<�뭽|�x=��<��Ѽ�AϽT�A=s�aZ�;�XU=������>�=,��=
������=b����)��ϧ���q=�68��z�;-�"�G��A}H�(�)���;��g;]��=>O%;����de<`TJ��~m��wq���H��k�=�l>��4���=�1(��c=Й_=����8Wֽw�>�p�����=�K[=��¼�V����!;g;&>d����;�	��#�>��*;w*����3<��5=Ow0��I��ְ�;tܽ�*<�W=��~�ߡh=2Ot<t>�����=]�&��+3=4Tt=\��Ww=�T�<6��q5\=��="�s�C/���o��xQ��:��=V�B�u!1��4м��H�J�[=��U��2�Fz�=���3��i%3��e=g½=�`�;
�����R幽Xc1�l8�=����t�;2��}V��x�J�F�d=H>>��4���<��Ž>�>����e�<Ӆ��=ܼ����vF<���=��>�Ҭ�ġ���
����<������=�̭=vs=�-5�Z^���}�=a�Ž�	�������Ӗ������
�L�彝�o//=Z^H>�2��:����&��|꽜&=��G��A>O뉽T�4=f�b<��3>:����W��͖<HD6����?������O7�=�Cq�YW=a\�=��8�Xj���̺==K >���=�|R<`�a=��=�`.� v��f�=�]��zi�����+n�_lO>I�=:����=���>�~#��.��s�޽@.�UU��wU��W>� ��*%���{�X�V�L�[<r->g�=��>�δ�<_�>�U*����I��=�pp���p=2���1=� :�aS2=�">o�#>�~$=���C>�%�=���=$y���v=f��<�-�=������=�T���=�H>�/}=$$q<�$���=\��6e�<�V=�&�=i��^�=o3��%>=��H���s�,�>=K�=*@J�gE�A>��;�U�<)�����"��;��=�F�4���*=�&�=��=�Q�=�9���N�}�_���=��<}i�;����޼ap��\�9��:l2 =.�=Mٽ�;/>�s�=�<y�H�ǟ�� �ʽ���=0B��B�=XWM�E6���[=Tx��+����<W���/��&>�#��b}��9żJq��(�Լ򠭻{:�<�����=�8�=��"�<���<v<G�=�A>v���H=G#��m�3�h��=jɎ=�(���4=�Ix�v��!e=$O���MV>딳=h"��[r'<ru=��<Q g>��8=0aM����=�م<���fC�;Vν���<8�>9C�;�ƺ=�u=~�<�ֽ}k�=B��7�=�z��e���8U=p���P@��Ƚ�b=P��=Y�/�b�t>	�C=��=��K�^q���=O;=�N�bAB=4����/�=,'�=�<��㕽d��Ll�V�)=�W�<�
��]���BW���<��c<�Q<�ǻ�0M��Xλނ	��e2��f�q�<j����w��\�9:4�=��m���>gQ�=����ʇ*���߼�f�xE����)=����]�н�>o��+��܇�<��=��8�a�u=8�O<H4</'��5��8a=&�>������8='�:��R>t7 �ڢ.��֎�y�wH�=��-�����)=�W=�	;�\�V<X�c<� �_)�=� �?�>�С=L0�=�$߼Z!�;Y�ν��P=��[��g&��x��4��
�ѽȥ�=���=�P.>�ٹ=���O�J��d�<��E�=�����s������=!~���ۚ=� <;Xc���X={O=�'��vhW=Rr�=Z�f�T=��>,K�_|�;a�A>bI>0R�_����7=�Y�<���=p��=!-y�cvO>�m��z+n����l�
��f�=�����	�6X�;Ej��+�<�0=�T>w`2=��=�C��~�E��˨�<�2%=��w��*q<�m���U�<7S�<�9�.{%<A�%�_ׅ� }�R4���6�=*kѼK����m�e�=�/��t˙<$�<����@�������҈<.��=' \=	 �=�K������(��������=�:-=�<=�N�%�=�R��1[;�@��6R �	]=��~=��=�`�=;>�=V���EX���=�3 ��|�<�I��
>[Bü1�y<`#�<���<�Y!��4۽OC����uV1=�+>w��=���Sӱ=+>�aW���3��9��t�=�]���p=vl���>=�?t=Qc��p���d� ]��c����c�fǽ
�=�d�<������/��< Զ�����&k�+7�={ɾ�^�Zj��Z!M� �n�/>C:���z=�0�=:z�=ڒ��V�L�=X{�=x߻��=��l�gS��M�o<�u�����<���=��?���R=)����-��=�Z���t�=�Z��l�=^���o=�o�b~����ý�Q�<��=x�ʼ(��Pk���"<�0$�<0����V'�3M�}<�������=����\�ӂ�<��X<�q�n�=֕���û��:=�(����=b�Q�载�u= 9�=��c�y}����;m�� :8�~B��[�<�)~�K�Ͻ���N� �o����~���]�=,Gj�Q*��n�=\�����ӽى�;�=G�>�͖��̽�I<��3���<���¼]p=��DU�~��=T����6=!T뽧&�=肼�φ=�5�=ի���=>��y�ZA޽�8�=�� >��A=�;�����z�0>Ӂ�=]�q�h*��}���E�:��<=���<��u��>ɔ0�gVü�5�=�|�==o=܈u=m�>G$��{�+= LJ=,Fq=����kI6�����j�;7������`I�3��<S	b=e��=M�=���=����X��N=ljd�~*
>�u��|��������E!��۽d����\��R�=$;�[U���=ΐ�=�6f��g�7^�=mQ>p���ArL=]==>�����=U:�g5��G5q=M#?<�h<#ϼ���ҽ�Gk��D�<�Mt�*F>˾+>R(>�U@��.-=o3A���+=뽀�?����E<=3h%�c!.��$'��4*=�O$</<�䂹<��6��i ��QڻD2�=?�G�n=
�V�S�=@1D=?�=؍=f����<^�<?�<��=��E=�0
<�.��?ػ֝�:�A�=�
=����ܪ�������μ�ؽd�(=:�=Aʚ= oW�����bv=��<�=
e�="�0>l�=�\�]��pV=-S3�X�<�gٻ���<�f�<��*=�N>`>#���ѽ�닼���=h��5_�=X'n��0��*���m ��|=F쌽	[<�u=J`�=(<޽&>]<���g��C��=�u��)�<��ʼ�>���>}w�}�T�����q��>�=+�R������Z��.׽����m�)>+��;f�==Ec��氽M!A>�*>N`K=B}o���=5�P�?��V�,<���Q����9:V=pDx�@�C=L�u��=�h��v�)��|�<qn�Ť�<��<�K�=v��<	·����;�G����>-="+*<Ʀx�����c�-�<�?��\<��4=�K�`��k��.����xl��S�d=|����e�:*�:��\>[��=pe.>��=;

=��꽅�ƽ?�j<�T>�G>e0ۼ��2�#�V�bH���!t<j�=�E>��<�(�5������B4=���=
Q����I=�{D�DS>�U�(C=�ɽ�dϽY5��f��=���?��E�=P@�F�0=���;��=k��6��l�< #>�����弲\<?�j=���=_�=t�E>������#>�#���_>GzW�ݦ!=z�=#�;�s�=򋤽��<F�9���=7�M=.��=�j�=\��rM�>b���
��\6_���>Ε;����m�>� ��LA��,���=���=�z�k3!<��<��<��V}���6=:�d=\�!=�uɼue�L��;��t��և��{�="ÿ�f��݌��zM<@~y�b�:�Y�8��u���"=�+�`�����̷=�P>���=�0��H�;��"��8�=o���=�<�oL=US��+��sK=.�>FAP�I��<A��=ˡ�=�^'�b^��� �$>֡n;Y|�>��Y�J6�8ս5a;s�<?�:<}�7�˿�Y�Xn�<��0=0���Q��&5��<'$����=��<%1�v�=T��=�N<`Q�=�:��m9�X���!�<�J����=�ڃ�$�=�%=��G>?W�KǷ<�� ��d���=�{"<[_Y=��$�L
ѽo�=r�F9g��=Id�=-�F�-�I�(��=u5��2��̑=��J=�0<�KB���/=�~�<�	=���=��=�=��eE�_D�m�=���?���0=��.��h���b�9p��Rk<�ʸ=Ӵ�=�=�"w<�>P�$�W����9=�>�:��=���\����pӗ:B��rg=��ƻ���=��6o~���<�u���F�=��=R�+����=��;=S������ی� �=�ɜ=BO;>�Q�=Wp:��������t��'U㽾G��B =�z�>{m<�Ũ���ػ^���y�=1.��(w�A=��=�E���/>E��M��= bʻ|R#=c\���M�=�n@��,!=��)>C�%��=��ӽ|� >�F�<U��Q�>C���vdk<[�6��D@<�̨��}
��OT�,��ν�P�j=�*�0�=6��_�b6>ܾ/��l�mJ��o�/�i
��y��<pG#=f�=3�|=���={=$��N&��^�̡���> ��=;V>��ԑ=���o�<TN_�������[�f�D������}�=_�u<p=�=ЅQ=Z�;=A�Q)���W<�B�=�����>r7��f��=��켎R-��?ýk�=c�*��� >ْ=V馽t煽�3����[=ͥ���5�=c�=�-��=��G<�U��/��К=�.������Ɍ��J�<��`%<�>��9�<d��>�T/=�
�`���{��3=�閼��?��t,>�o>?�����䟽'��~��<�0����S=l�
=�,�=`	B�S�=Cې��G�P6&>��N��@<�<0L>�&�<l'��U>I>�����<=�N���,=����\s��7�;aB�=Z�<έ���=R 뼐��=��=�"�=�Gr=/Ԝ<�������=��ֽ�K!<��F:=ֽe�(=�?^=��׽��'���=R6i<�b���w=6,�=��;>��\��A ��A&�ՊT9�w��z�=��::��=�Kt=p����=h��'W,���<��;�A%��U�=+?i=�
��B=V���qW<(���L��c�w�w�>�z=`����O=��K�y�>0��=.뎾��O=`9V����<a��<ِ��j����<U>���<�G���<�U��(�a=�>؆%=��).彲~m�Pn�<���;ҝ6��0>K>=�= �|=55{��y�F�=)�=�ݵ��X=@��C�B>��Ⱥ��߼�K-=m��Ϛ;�+ּ�k�= y�>ר�=�$���-�I��<���:���6.�!>���=�Ŭ=�cd=`��	�=J�<�(=��<�F�,��=Z% ��Օ��Q�;�@�<3  �M���PV佝g=W��=�%�5����i�f�=C8��۵=e2o=��B��޽�R�q��.��:���<��f��b�=�c<��~V��,=p�=e����㼻V���R�罤���*��,�=b���E�껦�>�N������b=����c��=_Ԑ=�0�?�q<�k��;��<�_C����D=@�� ��<���7����|��{u=X!̽�_�=�h(����u�j=���<��:>�*½>�(>(K�=�����V��aIj=,
>�EZ=��\<Z��X��I�8��=e�'=�^��Ru<yfG�?m4=/��>�/$=����v��=��G�z�{k�=>>JDB�'׼_O>�z�=H>;>���#�
=C�����=�&L�W�^=MO5<A���o�=�5�FHx��o�<٥b��¼q܌��S(�'���I�{<��>a)�=:P�<'m@������� >��Q=SR�ϣٽq�[�b&�U<=WI�=G|;��+��f�:= �<�����=��=�`�<�f�R=!p7�� >֤=�!G�9�1�<w�Ҽ��l=�^���8�z���ׯb=������=�����V\��@����=��=�7[��=��<��һ��;�W���~�����z���Ff=���=�ي�oN����3w=Kv">�*�=�<ɼ&��="z��̵��w�<�;ýW���e=�K�="L�����\ϽFze��*{����5)�C�=2�;����=e7��_�<��;]���~}ʼ��3��K ���k�a���޽P�:ui��*	�=5���<%��=V�{�������=��ҽ!o漏Q�Z�=�	��Bފ=���vb�<b����-۽l���!�= J�<[��=��G�7�=х>��6���*���@;o���4�2y����J��r�=�mP�|b�<�L^�c]f���;���<Sfż�����M>O=��V�=.��="���(�����Po=���e޽�]Z=�>�P�=ND����)>`/=��g�u�;���J�<׽����>���������"�U=�ژ���w�Y����UƼO��J�!=$C��4�,�}y��ֽ�8����=�����0R?=����P�=���fn_�Y��:yA�����=�'��F��Y�=߻����<���=�ݽVpc��|.��Z�(~X�8k�;=�<��<L��F��<.=^=I/ԼxὠO���; K�X�=�7=Uk�=�?G�ڪ��z�v��a3=�0q={��<b���\׌=�5=����,Z=�w�=B_��~1=j�\=��R=�����<~X4��V޽�ˇ=,�>}�+>%=�k�=VE�=�Z�=Md�=�M;��)=��V:�����Ž��
���=�6=U��=�6��D�3��j�=0Z�<!d���
��x��h8<#���k�ܽ��h�{{>C>�	�=?�=7Ϗ<����ZW�������<�z�?�3=t+̼`ý��d����@h��C"�<��߽cz'����ju�=�'�<U�p�������7*���ѡ�,/½��<�EF��u��Rؽ�瀽�M �h�<� ��X���~l=2̀=Q�=���=v�^9C��<� =�<p=/ �A�=m��<��5��=�<f0ռN#>����@\�=�-Ǽ���;�=7-b��9�9����N�f%>A��؆�<�KN</j>�́=6�<۲�<�,�=)90=R�z�'>�$�����T#>5'�<T֧�Y��=2<M<�b����<P�`��Y��u����6����ڟ���d|���P�?F�=�W��t�>��1�=�x���\�=��ٽ����dF5<�d�;3`��7�q=�<x�=���=�y�=�=I��=7!�<@2���%�<#3\=t2�'�Խ |�=��+=T?��;=re�<a4>��<4&><K/=���=��i�{Ah����=��_:���='�V<�;g<�/��#�r�� ֽ.��E s=�F��x=A��=�?��ڟ��7�=D�=��h<�'��u�J9l����<_�P�!���a�<J->::�=��;�C�<~�e>�b	��=��15>.�K=���P�=L�=[��;�흽�v�.���D�=U��=�ۇ�̳=����;B����	�eD=��
��"��VA!>O�Ͻ�o<���=/nr:q��=�b'<f��=��H��Sz���!<%�/�V�r��w�<�ly�9Ǔ=�F�=3f＝�=�v5>�� ��щ�r�B�Q6�=���Sq>�Y	>� ������d���1཰�:�#V<ve�=�6�=��x�1�������������@=�Ћ�tI�=�jҽ��'=�^��Zf����`;=o�<ּ̝��=	ά=ɽ�=%�>=�<�IX�MT�=�Y�=�@�;��(��=,⣻`�9==V$=n?�;D�C�Γ2=�v�;�7D�	�ͽ\�����=�v��V]<]k=��:=��֗u<݆G<�>��H<
`�=+�=��0<AE=t�9��Ȑ>,-⼢�2=/S=�_���T@�ǯ�=���<���S1d;�O<��A"�c�<�����`�=7ǽ=�?=���=�'_��ⰽ�1��VQ��>�|=�<y�Y��״�1����>��>��&=���<Z��S��=�V=ޓ�<"���Kz�!	o<G�M�G��;�J�=�C���}J�4���'���=��u=D=���/�!�j=#{9��{�:�����l��j.<��0��R�<�6L=n�νq83����=��㼊`p�.CH>��1<`��=BJ�=T����2Ľѥ����ν�C=R�&<f�N>��==���<��<��A=4{�=���Ʋ<��4�=<^��롽�疽m(��t�;�\��j���K=�b�B�%=r���y��`PE>�=��e=�o>c����
>+y�=�S��]=j�	����G�s����d3��ɱ�jm3=�eU>�������->��n)�	/$��=��,��:)>����L�<5%��T����� =!��<Ee'��� n�#tV=����H=Ƚ'�1>-���">��a��p�����9�T=�wf=n�H=��`<�Ϻ=|�콶U�=��<.��=�=�T���������l>��>Êq�P.{�K:<�j�<����=8�Yjü��M "�;��ZW�|����">��>h�>���m�^�/�۽����#�=�<���O8<F��Ľ�?0�m�y<ᦕ=g��<��=��=|��<6��/�5��ע���=˱ۻ�0=b5-<6��,�v��»�f������gbZ=&��aƥ<]��׶:��C=���=m�w=Eu�=����E�=�AU��Wh=���=�ă=�)i�<��0�O|=�w����^�a����je<Gc=M�D<�a�=�~p>h��=���/�Z���vb5�{���	�=z�U=���=y�V�����27�<�\�:Q�ཥ#H;���=���<|,�<P��<<c�<�f�=�l��	I����=:0�=?�>�����=C5u=�@�=��h<����=#u��C�<7�>"��=]W[�� �=�̛=쿰<:+.�����=
Kn�?|�^��=�)T=��<��<p�=acX�,��<�E��0;k=㫍<<�v��
���+�;-��"�{�=^,���V�MD=mP=���<F�<Z֦��uX=�#����=+�����9����<>X�<�iQ=��$����F,�7����y���u+<Q��:�=l��=�H�yi�o/��P���ݺ=r�ս��|��@>Մ>�V�9�ԽZ� <A��;"�S=T��w0�=ʴ
��X�=���=�ѱ=�,�<'���|�:�xt >�P���m;G��=��5�%��!=�\�<��<���=�d
>�Uu��b]:M�A>d2T>�ؼ�f���=Q�����=8T��B��V�1�Qs�퉇�-��=(
<���<���<��;m�i=�\��(r<X�a<y�=���˨��>ou��!�r==�<���<�k>�_���R<p'Z�Gλ'u��>�̽t�G��uԺ57>�6c<m��=:X-���;�X��V#����>��=^��;�
*�K+Y���ټ]������V������ &�'<�kQ=s ����
9g=���@� �ۨ�=�xܼ�8���^<V�1�IKＸxY;s*���9�0<Ee�(`>�u�u=�s��ǿ	=:D��f;�)5��L����s��"�Ƚ�=���=�9Y���7���p�q�6C&>0�<��2>�J�;�#�<��<1h[����������zɽ+�� 4.<��<<�@�<�#=�3=,��=���=�L&=b{��L�:n4�=����qA˽D'߼�=(�/��<*@��='{<�y ���@>*F�<���<��<�,ݞ=���=R(W�fh��A>�Az;&��E�=GJE=
T���y��ڠ�=Q ���(Ƚy)O����<۴ʽ!C�=��<2�V<�0�=B�<��8���j��6R�x��=bS#= XM=�'���j����=��T�x��;��=Ɗ>�	�+�d�=�<;�B�%^���0>p!���;`��=�q�S�=��G���>�:�J=/�=�go��H�x�B=�p�=Xm���%=������=@M����4�\��=@�j=ҟ�<����4T��H�=+�꽍Q��|�<��h�bf��xٽ�V=#3����=�Q=4��=Sp��:��e&D<ͫy�
2n=�=�@�<�ὶ�9�������;�N;="�q<���=y�<-����H���!�n����o�=��=�ޜ�Gķ���y�vlo<�^�����=�/=g惽e�n=⸮;̤���S��燽c{�k`(>��!=�Ğ�H����L�X���Մ=:�Y�N�o�@)�hz��cC��7>#xx���Լ���om<��2=��F�i�%�Lg� i�=�劼�Z=f�=�H齛MQ���8;��>�O7=��;ߺ＀���֜
�%?�=N���2����2ֻ��=I̼@��=�W�=����E=�3��4>��Z���->�,�=a����ۯ���I���D=���:Z�>!��<���=G���}+ͽiD�=K=��=��Y�d��:��=�A�=���=��a6+��ͼ��];���_E�r�1�}��=n����>�B>�Ko�Yp�=�zi=B�໚v >6}r�'�=��`=���=ɋ�<<䕙���1>iI��U>�Nͼ7o��g��=6��=�t�ʕ�=j������9�>ƃ��#d<@q�<�z� �,<��S��$S��;�<�L>=]�x=��<� ����;��<@0c�.Y�=r�<+��;J�Y=�=#���wu<N��ɶ�=9�6=v�*>I�=������`�<?����=0#�=8D=�gͼW�l<�o�;7�>ޚ=���=�E ;�ӽ�%�:����B=��G>��@=�0��=�:�������X�=���<��<G�2=]7<t���������k��> ��폽��=)���x/�d/������w�!RK�Wf�<��<>�6��Vu=��ǽĉR��h�=�Z\�q����k:�� �:h�1�o���>9mm=��; �<6�f��qx����<p�=6^=T�o=�R=�.<�9n�t
&�<(}��X3�8c�H���<ӑV=K����8�s�Е=*5��cC�=�q� 21�=�w=�#G=t�;�a��m=T��fPL>��Ӽ�q<��U�<�{�=����}�彗f<N��A�=%��
��.�<ن�+`9��Q��t����;xŽ�����f�<�M���|'<�ü'@N>x��N��=Uy��4���b=���=�c*�gݷ�f�>D:�R�J=7����Ѻ=qe���Z]=�����+=�鼓Ư=}�e=��e=����N>8��=��=�*���.�=2�=�uؼ�oW<���=ŗ�������=*��č��R=�×��ͽ�j�9�y�=|�=���]ݽ�ab=���= Q`<G��>j��������P=��%�n�=�"��1I|�Ko=�d!����!�>�>�`Ƚ�l����+��s�=0�߽���N�޼�t=|�u$-��eT�W=�N��� ��[��GF����?<�*<Vk�=-��o]`=�;�= '߽��/�p �y�[<�Q�=����-�ּ�bT>�Kf=�G>�R���zս1�;ic����>=8*��m<�ˎ=��[�.��=f�����p��G������=�%��V���y�<0�Ǽ���=F���9R<=|˽^A���\=+�	���vV���]�FDh=O,������I���!9�(Z��q�=s�m�:w%= iX=l�ջ�&_=@��.�[�;E�j� ���<�3��l���>n<�=җ��d�J=t{�=l^O��|<,D<h���?�=�/��白r����N3=�����
z5��M�����Ln�<3�ƽ܇�cC`��e=�4 >�{�=[���q͔=�l�=�w=@����;�ܣ=���<g���CTA>z�.=��l��FU=6�~��p�a==wW��R�=�a�=g�;�D�<ib=ˠ=wz_;�-�=�Ku��4<(>�B=�*u�==Ǖ< �強O�;�(=��F=(|�������Ɍ=���=��^�ɬ��ϛ<�¾�ׂ}=�x=�c��Uȍ<��=W#f=^A���<�4�<{m)�|"�#�T=샼Xҥ�TdD�ς�=sn=�B���m�=JC=��B���=�������<~�\�����j��p��<�
\;�G�=��J�����-;>h߽S�=��\�Խ �3>�Vy�������>=�Q=���=W�(=��=����'��^|��T=Ф���ӽ������`�;��<��=���7��=2�M�R$�=���;�e�<:�ͼp@<<n��=l�$�@gT>J���#�K�!��<l[����/��?o=���=�=yTݽ����j�<�4�:��&��|=@�=x�=�	>��W<�iM<�S�<t0<<����{=�2������B0�����qVͽ{�6�����A#=˔�����=sa�=h<==���Ó=<Z�"h=�q����<���=G <��=��=3���/�=�L=�K�dZ[��O�=�B���=�Ҙ�CPG��>�>�^�X���=�Mm=)�����8����=�F=<¼z �����۷��_6��ͼ� �r�v���<:M�=�#��=>ٸ��A`>ANQ�YA= 8P=�*=D�����=@Hs�1N�=χ�L�3<)���->p�z�:8���iἛ�=�����н��L=k&�=�/�=�7�<,��<ƨǽ�܉=9>����:A�;j���=B�Ľ���=t=y�=��<%/�:������=��=�Q�4tl=��=�d=��A<�Bڽc >���<���=R����H7�=���b%�=	B�<y�=iD>����9�d�E�O�Ժ���=E�o���;���<}����[?<��G���{�&��텻B�=���;�v������^s=y-;�o*�%n��<�ep=7�����=�<��'Yr��Un��1��l����=Q�����=L �v�K<kZ��rd�<vUz<�䒽�<�J��<��D>�\h��#.="m�=���B'��*���lz=����kcD����P0�%K�Յ��A��d+�=oCO=��>���=̆l��l=ňk=���=�Uh=���=����aCE� >�=�	>�&�=�&�=D�H<��6��N�kQ>`��^��>�9��[�=+�Ͻr<0>@=������$=��I<K���Ѽ� ����2�<﬽���<��<AL�=������=���<��M='E=:�<�@�=U��=��*=kc�s��=�o������.s�����4^=G�X>e�+��_��<=�k�;w�H�ˢe�`��u�=j����E��?>U�	�U��=�r[=�e����)9���<B�<K�����=�<=�5�<(�=��ڼTS�����y��<TB��.�fe"�^�*�X�&��I��M�>r>2:ȼ�BM=x�S=�F�=�L��؁�`$>�+�O���3=�UI;�,�<5v=	>���B�K~?��yM;��4�'>z5J��擽�:W�t���G���:�eǼ�>Е弑?˼����i<�-���R��=��=�"�=��>�3��'�="%=��k��'��E�"�`.�0����e���'�1H͹ɂ=	=��k=�1D�Q{�=ڵ)�Πڽ�
�<�*p<a�<�W��A\�:�2J=��_�'��z�!�L�==-�޽�PP>׃2�������< �M�#�u������	ռ�u¼9�"�?4ٽ�=�������d��J=dݳ�__�����<���;�Y����<��=��ܨ�=�=��2f�=�Vx=�t�=< �=���=�5���Y,����v1<M�<H>4��<�(�i73=c�>��>���������̂�<0���cq�<����=���=R���|�i��=Af�<�e]��Z=�>��p�H�,��4�=��<��=����=Ғm<��=����_U=�����ʄ=�x=V�̺��<�a���>:�ڽc^ۼ�3���8>Q�S��?�|��<��u;;Ӵ<���=��;=\$=jF��D�>N�%��Ɉ=�HV=Y�<�	Z>��	="M;�ކ�ER����c�ڼ��<$�=��=iӸ��^���=�{;J�ɼnȳ�Ӏ�`ʀ���߻tUx>��D<�eK���	>�Jj�U)b=������0>�r=�g=�}P=��(=#������M���3���k9�=�=�e���Y�h�C����ڬ=Wp3=��J=�4<�)����R=_�����ּ�
���~ս���������~�)��=O�=~D��A�=T$��P���Y>����'rѽw=�ہ�s<��M5�^d��UA=�Dp�}��=Bl==5u~;��V������>��$>N�O��>=y�N�����++Q=���Y=������=n�<�}F���n�
�4�MT�<&9|�����_���T�=��<6?y=���?� �nF��ޓu��S��ա�=������A<�v�K��ʢ6=nh���>�e0�^_ͽ��x�#�a�P&\��i�<�f_=�7�=G�<	����<�a�=�x��� ���ٌ�R�K�MJ�=��ݼ�X�;tÎ=Y'(=��;1�d=S�$;x��l����������=heY���L�c��E����q���ս6>�q��=����*'�=E���:��=�ͦ:=��<��Ƚ1=?��<�� <�����9�_�����w�U4꽦����i��O��=ťy<x�t<�wj������ý��2>vg{��.���@>j���K~ͽ�"N:�=�=���3�l='F�=��ӽX;�=��=�R��e��:}b�=��D���x��Tڙ=�Z=��c=�r�����<T]|�>�#�^�,='���=��=��o����a�>�7=��=f{�)���Ay�=0^<.��=`������mHн��L=���<�(3<S}�<:�X��;!=�.�=A�ѽ��+>�Fz�w8�R��<�2�*}��1��_O=:w��8=#4�P�;J�罱�p��.�<wD�;�]�?�R������3=��,<m��;��>�֟=�J��o�z=U�&>�*����/�:��y-���;yd>>.8�<L��=uk�7�<�ؿ=��=��;2�G>_�;-��=�g��
U�K]��Q`�<7=G�=Z��<L��=5G��˴=BV����=�X����4�����1��mB>���<L�!>���<͔��5u>���5��<>�/=:z��w������&�NC>Y���G��<��= gR��w����<MS��E̦=E�=�}i��z�+X
����<1�X=+��"t����9�v|>������s�|.�<ZJM>���=q���[�=��>.�������D�=u����:�=�Y���=*̔=j�h���x<Ւ=�4��<3<}�>t�@���W=&4���mP=�.���I���ek�7'H�S��=D(ƽv��=�%�=-�<_�=��\=��0����՛=�Y��w<�����>K������<T:�� ���A=��<�X=)<�ĺ=߷��Ȱ
�Tx�����8�<=彼L+�=������=mv�<�"���`�;?�e��=�YS��s���*<*.��3�=S]��!M�=��꽲-=�<̻'X���	���,�=�Ǽ ;"<�h	����<S�k�h�1���=�/B=(�:�u����5��M��d�=V�b�nE=�d>\��\je=���=�\���z3=	O���6�v/Z�����8;��>�K�������)>�p�?�#�%_��"k�=����H�==���8W��N���覽�����u�<���=�΃=s����)>�<� '��=4=�w�*�=ڔ�WD�O�>s$
�<Y��=D�8��y�'�T���G�N����j�F�r���=�O��V�E��%>;��?sT=�`,=�+�=f�M<�<����ٽql���<����d7�<S/(��+ɽ��P<��6<p�S=x�Ž;����s���n�U�2<��&=�*�:H�G=eXV=�N����{=Lf��m½���=��=�N˽�L�<w?����=02>�{1=.�o=^�m >��)�Y��2�����C=��=<s�=bA��@��=\���ݘ<�B=��(�܇�=Lܽ�q½Q��=p�>hʽ �j�pټ�%ƻ��a�2'����<��94��<p�m<�+��Z�v<��9{���5a;1C���9:��=�!��ڬº����6��=(���I����������>߬=�\p<&�����������-��Y�<�s>���̽���=d���|=�)�<wU�=哽2-_��K"=!H޼=;W�7s>~�I�,H���5�=�����	>5*�=�x��@�=�����,e>aʺ��+h;�T�>)J������ϒI���`�������a�k���e�h���*��ڍ��ၽ�)�����=�
���\�=;��=�`V=����@=C+a<W�c=(F?=b����ImA����3��a<��/=bɆ���꽽�I=]s�=M<pm��Ĩ�j�#�¯��5r����0���<��=j��<!\�P�<�+��k?<�ݼ׉�@>eڽh^!��S�<�c$=��j=���/���<;�ƽP(
>īĻ\A����-<{׋=���m1�<��>4]�<QD��Oȶ=�ZZ��2=� ���G�=I�l�"��@6ývh�� ��L��*�μ�M=~_��o���^=�y*�<�:> ��o��=�Y��}=�e��f�<X���M<Y��=󝅽���D�E�|�H�U�ڻ���=�2Ͻ)����d�����%ͽrB�=�J�<Z�<�!=�L�� ;�=_r����I<n&���,|=��a<��>�c�<��=�F�<p[o������p,>�b�=0�<��<ɶ�=<Ow=%F?�Z�=�� �1��:九&�9˹d<��<(s��v;>n���=B=�p��+�<�ܽ�3u=��a=�Tļ޷�=1�Ž�G'��QF��&6>�z��t�G<�w��t��ǆ=b�u=i�!ڽ��>�#t=ٳ�=�1<ش��N�
��!B=^��O5>��޼ۭ =o�=ܻ;;�Ԥ�����h�W��z=y� ��<8�=�	�Y���
7>F�۽ �=���=hv�<���Y�%=�bD<����]>&�=ik���<"�	���ܼkW���t����=���=���=�h��w�r��	<s�o=��1�֗�"UH�kV�#*o=����d��=�Z_<�,2<�텼�r��8"���|�=t4۽�CϼJ��im�=�EX<��=
��=�3j�!��a���e���=q@���֠<�.�4����=�)����=FOR<X4^������[�&f>>��~<�~�=A����<��K>m������_�=�S�=���<�I̽ϡ�=��>�]�=2>�M�=e���
]�eB�o�.�����j�>�s8�1qĽ@H=�H�=𕬽?1T=�C��W˝>��<��=�j�c�=����=�D��c#�GG���=��f��J=	F���_.>w`�;,�]@�'�a���U���l�>h��=L��=ةn=��"<����  >��==�Z�p4l=<}2��A�R�� ߣ�V\>�2?=��=8�=>����� �qh!=���2<���<�#>۔>�?�<+���XRɽ�x7=�:=�<�=�Y>�׽��M��`>uh���=��,"��}L=v$?>�����&�<v?�<���!�=(�v:	�ɽk��<�r]<�T�E�#�N�����0=�É�y�w�!��w�>��&=:e=D���$�^��E��B?�=3�C�V��<�,���<[�
Q>�K�16=;�<YH.<$��L�>�}=v�4�ֵ�<W��=���;�lT��	6=����=�4$��z��*����>hY���*=���<|N�=8�N=R��o�<�>�#En�`GS�V�9=׭c����!�=`��z���z>�$��Y�=vId�ij�=@ɮ=�@���1>q�a��N�s���S���Y�9�
#��
=&�P�>��=�5=��3��<���<B���=L�=�I�=
4
�eH7�ړ=?���벡<+����=�}=���^1��YJ��;B�X=�މ���^=��>DӇ=���=a�<c,g�K��=h��=pI��r�=��>�H@��/��Lj�=�n >�g�=TC����=&<(=.�;>}<�<��ƽ��k�D�P=����퉜<���=�-�6��=z%c���3=rR���N�<�8C�}s�48�Տ�p=��n<"�.<����71�<+����Mܼ:�;CU=hE�=^⽽]��^8�6�'�-�=���<���,�l<�h=�ҏ=ʰ��=��=v�>#�%���м;�:=B���=��o�=�-��k��=8�=�E>�|;>�l۽��c<����}��O1=!n��+c�=t�m֟�/D��,��=���==�D=Q[����<=��4A�o�=[t���8��]�f=#���Â=<�!>O.����߽�h��D��:��<�3��T��[>ۣ����Y e=�L���Ʌ�
>��%w�;��>��e�hx8>���E��.���Z��=H���&��J4��J�=���c�<+	����<<�C�-]��)g�,���ݠ� �=����ܽ:�=�q�=Xc>� �=�����ϽI|�=j�EW�=��н�-���q�P��h��[���������'b����y=pTM��qe��ҽ��F���>�ň��`�';�=�[)>1j=$/�Įm<��:���K<ܫ<Lp��D𝽦Ҽ���p��j>f�=G�}=��&=j+
�e�:=�X=b=���<�䟽AH�<��<=¨�T?�<�����=��=�v�G�󼰄2�=m)={�=�0����<�B#�q&�<$$t����T�=�\+���=�Y�<�j�Np��ƫڽ�_ؼ��@�;×;��x^���i=$�.<ls�<�/½8ט<�L���޽o��dj�=���=��=� B���v��	:��?=�>�<���	>Žl>����ֽ������:Vpܽ?��=H};>���� =��컼���s�;_3V�3꼾^ӽ�*>1�|����N�,���#$^>��v�u��<�����{a<���=\�=��ýW߼��*�;�#<�ۦ��S>᱇=�פ=����<�=�Ͻ��:�>-1�=ɋA����=���;Iz�sǆ� �)>���q�M=2�:>Ӈ���Xl���G�׸
=�<�`�~֪=��+=v���W�l��qW='�>/��=J�D��/<��ҽX=q-���c�=�j���	
=zž<yc��Q�h<༂<q�s���0�vn�����'�=�g)�S�=x h��9��c�{���=iZֽ�R�=�Eu=��?=��
�ܓ�$�?�5���?�ܽÊ�<�Db�P�t��G�3���&k�;=O�=X�=�\�=U��=dJ=5k�<vbS='�<�.��������<�x�������;�ҧ���=�A<�5v=�O�;�v�<C�H�ﴖ��=��#��5:��t�\ɼ%�:<,%���ʸ=�\�=Ћ=�.[=�xI=����bM��_;��e�&���'	���%=���a�#>G=W�=��<�*�=�j�=�= 3=j��eݷ<OI��X`"������E��./L��=<�<� ��t[�=ȧ�����;�=_"w=��<O�%��]���:�1����׼F�=�����ԉ=j���3=b���?����R<�P ��F5��G<�ъ���T�w���|�= 
;���X�ѽ�\|��U�;�"d<�� ��J�=�/>�W=�,�~)�<��D�&#N=>�+=\ρ��X�=)!>�����(k�'k�<1�=�8��yd�;�<�>�C�=�g�3~=��<�9��?=ql���c=웉�NLC<���hf=&<�/�3=����Y�+<�^��+�S=$����P��A�<o���y�Y=@ٰ�[�=���J=�ۈ����T9�=W��ωI=N�� �3>땽ւ��<��=�߭<�̹=NM/>�y9<��=!>:�=���u��=����0T���Ѽ��˼G1)<{�{=��!�E�W���%��~��>=�FO�S��;�g{�2�=~�r���{����=�5=li��Ik��bc� @���W>��<
�<hjf=Ȓ��E���&h�==�޼'ɧ�5���9d�渽����*{=Z���3>)�~<�k�4"���<�M��1=}4^=��>�@��9�=�8U=���=Ud<O78�\73=i
��W\�w�>"&>����g%��F���Ą��`*�9�?�RaP<�_q��X6= U�=���=]�I<���y��=`<��^%�~������=�I�=�6=�u��<i���=&2�;YN@;��b��0'�:�=�*	��6�U�	=ew���������=�隻*���L�}�'�����ýr<3�m*��8ɽ+�=۞��c���mm>n.�<��<Ӈ:=�n��05>6	=I���悽�໽��!��5��U�<۰ڻ8}y���J=��]���<Ȋ�=di>Y�/����ʼ;½Fp��ki��v��=T�;0�[<F =7O����½�)>��l�ĕ2�&���C��=g�9���2=W��<��^<|4P=',2>���΍<Br$=����B;>)��<�(�=�	�ڀ�=P� >%2R�����Ԋ�UT�<Dy*<Λ�<�>=�+ƽ�i�<*�X�Ц��9� Q��O0�ްм�KQ>�{�x	<��=��w;�0���Kq>��=���,�<�h=�l6�<l=�Έ<��=��=���;z��<�=3���	��=#�� �U<Ϳ!=&rQ���� ���}�=;R��ArT=�줽L0[�a�;+P����T=:;�EL{���Z=m�=z<\=J֢=�Qn<�1�r�>�j|=�=���ӂ_����� ��=3�����=�����|��F� �1�% ��9�=��8�"<&�ǅ=�s�=YH�=
�H=��4����:a�q�߼���=I�c<�(��6ޕ�3�� �=q��=�]�=؄< �N<*�w=wm���i��|	�=!�/=�$=%}��
>���[>;���ѻa.�<-u�=�X��:0�1���*w���	K�R��t3=8I��ܧ=�>2F�<�!=x�3�l=*>G=D!�l�=v��=ƻe�S��=��c�b�s</ʼ���<��=S	=X��_L >r�3�T� <.����>	��=B�����Ľ��������=�(i�= ����9f�j�f��ꊽ]�=%��=��<�=�(�<�4�.�>�1�T��=0���O+>Nu��Y���Q��=^q�;�v����3>���>s>����^� n��͉����<g���6=��">m�=�A�=i���IǽW��=�l=c����<O�(;�`���a)=���t�'=1��`N�;,Q;�'�=�zɼY�d=�7����5�o��A=�4��a�p=T=�=�Ĺ�"������={9�	�=��Ͻ̏^=r��;�	=\D콖�=����Z�H��J�~�x�y�O�ůT=� I��y(=B�N��vv�i�+���8>i6N=a���Fǽ���=�h�;^t':�팽���j�ں^�=ʾ�=�A뼿c=�E�=B����<�2�=�Ͻ}9�=�]$>�f�u,}��/�ߐ�=���=�6��U�<0�=l�ںx"=�Vx<nl�=�=/[�<�( ��6�<�G �'<¸�=-�
=N�(�|���n���g������l8�=g"��ʩp�n�=�A�!�=��>�S���Ƚ�<ػ�] �n�=�7-�ͧ�m��=�&�=l� �K#�=Ȯƺk��=^x����=�vȽ	����YDA����=�>~h=鉞<���s�P�[�=>�p	>z��=4u�=͘�=s��;�v5;��;&�_<x`=x��=q ��� ������ծ��(�@�н��W�>wP=�Z ���2�b_7>s�ս��<�@4=�3�:�W=FZb�Fyнq�U<v��B�z���=OL����=4Xܽ�E/�	�н�'�;�la=0;�#$e��[=&���V��y�ٽߴ���P����X=��<=��g��t�=<c�=:C���7��/��(ݪ<�x��(�N��L�=d+�==}�=�"j�=-y�+��<����N�=�<7�>đ�=��"���㽻��=\��=��=�2�=O�g��!>J,Z=�e*�dڇ�uB>~��=�>�͔� �V="F���{=���=�X��`k#;Xa}=�	Z>�>{V���Lj%�:悾?% <��4<7�Q=7��=�N�����?��=���F���9���
���J��wᚾwg=xP�=�=���;�mE�lu&=�h=�}��yy<�H�<�I;�7�?�¼�=��C�Z�9=B�V=F�o=?9;�G�;�c8��֧<4��=�x��.��$Lٽ�{�=�:ݽ~"��م=ԑ^���_�W�=�/�<=��<�[�Dx<�Q����=�v�=Җ��w�ٽh�x��!�-�ؽ����z��RO=O~��"*�<*+���<�Hw<[�[�s��;h.�7	�Ti��6����=�>>���`�ϼ6�ؽ/zP=�lG�T�<S�������#}<��1>�x4>v6�=��$>��0��<&9���4(>�#&=b�3<�bȽ0��I��e��
B=N�<�)=Ɣ:=�eK=XFƻޅ��t�'�8�S��=�=X{�H ��]=b� �Y��NE.�Mo�=b=�;�}=.Bؼ|1���N<@�9>���;�y�<�r�=��F;5�n�?��=U�<2=P���$�;)S�?��=�z=B������[��=[^ٺY>'�΅/��B1��R�<�?�#�2=����<P����=s���5�<�f=!Z�AӇ>R�˽�(�=0mK>����2�<����Ғ<�i�j�Q<�8>=	��=�U>Q�<}�����=���=�;x<��T��>ԑ����A��:���<���<4�=�� A�=f�~=6���/=S=���Uk�=Ó>j-N�1&ܽMM�='�^<���3��d��_�=�N�'�=�*=��<�=�W|=�`	=�v½(U��u�;���7<L�2�،�����=~����H�=Yi�+;���s,=�G>X�䇯;���=߱I>�TC���}:���ޕ�(�R�c	��,m`<�jx<.�m�����_�ĮC=�"���ɽ�(����<���;�C=��|��)�<Ph�2���g��cm���W=�&���Lw=m�"=5K�=�[�=j�&����=����?Q�����v��{h�h=�h��(.���?<TvO���:=O����=��j;����^U�����<�Q=5@>�4s�ފ��+�Z�pp�=qHR=`{>va@�a68=@�>���������=�K�=Ϣн�X=ʖ�<���?ż���Wl��^p+����=KX�=y�=`��[�<�ԽZ�<}BZ=���*(ȼ	N�r_�K�>�%�=�偽��=�$�=( ��򍭼�Ƚ��)=dE��x������[�"= �N=G�ͽ>{�<�|�<�s�=�y=X���M���Q<��ͺ��q�C�<聽:�y�)�̽32�=�G�=.���κ�g,�DI�<�l��7���=�c�=��m=�}�N���bş=�zŻi�gE����=u½�d;)j=ͪ�=�<w&_��'��!*#>j�<��½)�n;���;�-�=�a6>{B����=��>�7O��
���o̺n�=��-|�=�yv���>>T�}={ӿ<�Wּ�s���l����< "��v��=�*=ЦH>MZ�=R�c=%F���a,=ct�<�g����
=Ņ�<}P��>m|���ݼ�Ǽ��"�AL>�'d= L�r��G��=��j��D�<,[=��˽���[�=x f=���<Uݠ��}�=ή�=P/>�%�������A=X�d�Y�$=c�=�~"��̽D��<6ۏ���/���B��y����/=# ���^<:�=>��=���;��>v�;�L�<dǒ�e�=����sQ�,	=Y�=��I=><�=X)>V��;&�m����(^\=mH���x>��=z�=w�U=����F�8�=��;PI��=��:[Y=�L>�c=/,���"����=��=���=�V4�=~��=�2�=�Q>���=-O��j >�k><ā�<E� 4㼋��==�M=yW�<Y�P�)u$�d�,=
/==>��t��=�M�=`����+��(|l=��:��"��&�;U� >@$��0�ӽ +[=��S��j=��˼Z�I����=�X�<���������`=��d=-��B<ԷȽ9���}�=��=�|��%�<..�=���=��%=�����=ؔX=Jm�<���=e!�<S�o=�5�=�H>����)��=���=i���_��@���u�=��L��r
�b�<��=��.���܈��A�=~\��::U>t�	��Y<�_�=hY׽�4�=�ټ��sN=u:��$���:�c����5G=���<��\�ΰͽ��&>̞���u�=���<�ּ���}[>�)�;F8�=#����"�!�ǽ}$ýe�	<�Tb=�
�߇�;�>�=�T�żf�5���u;>ۥ
=��˽6+r<�>/u�=��2<:��n��<��ؼ\�q���1>��;������o�=��Ͻ���=���<��J<�=���=q:��5۽4~w<Huͽ�K>K$=n��<yaW�=9�=��s��'�<jH�=���9�2�Y1�<8+�=
�������ɻ�;�=��=�c�;V[����=kӪ��Yɽ�����/<�َ��y[��=�]B<+��,9���_��.��=�yԻ?��<���=e鈽�����<�7�<t��<�E
��K��������ӎ�=��ͻA��"�>�`k=��z����?�2Η=�r��������ʽ�ӽ��e=�3<=a�����=���y�>�>*�D��(v�j�:��M>�@���:{���=j
�=�d�����=���f2Խ.�4>a"�<�h:�t=\kY�J��O��tɥ;Ƶw�X�6�5��=�%������s ��Ȧ=���=�8v;�l�=m�U=���a�i�xs�<�(>=8aM��sȽ���@i���=�	 >M�=��m�3>�s�����<� =�?>B���$�������_<=��.cU=o�-�?�=[5�������漉%��C�C>ci��f�-��]
< Ԃ>���<�_^�m�fd/>o��<��̼\�ڼ�u�;���L����ͽ4S�=H�=΂�m��|����������k��벙�w'��)���8��A�½՟D>�a�=
"�=�K��=J09=�s=�M)=��¼��Ƚ�Æ;|;�7��=��ռ�kU���_;Krջ5�����Ľ�w~��h=��P<��BN{=�\�;*!�=��߽��O����;ߡ&�����Vt;`�#>�O��Q�;�/F��ǻ�ӆ��K���F�=kT�;��=���	�����1>��:>۟ڽP�n�H]�;�ѽ����%X��\.�3@!=�.=�i<C\߼��=�����S�=?	�jc�=!����/=��=Me[<���'�����=����Hl0������=!I�:Ky�=�������X�<��+�%=8�"=��!>E��=e��<�����w�I=Ƶ���=uU���)<�9���9o���={=>킼Cn��:�!���X=����X����=���=���=�J`��b�< ��+ :|���K�:�@>���>�����hd<y�ǽ�?=�ڧ<��b<.��=$o>	�鼊E��޻�=�m���K�<G�l=�Qͼ�(�=l�̽�5H=�� ��G�=l�B=O{���V�sd��f��*�=�p�<Wϔ<4R�<�Mj=�pc=w���&�>��)�����<�)��1�YO����=В<(I<���<hƽ�3,=I`=.y���a=
���.3�{%R;4��=��;U-�吽�ȶ�y�=|@E=7�>^4�1rD�~�[<��ӻ�@��{�����;��=�"�:<�8>�h>j�=Y����켒��:J��-���� �`&��뤆�΃>&�z=�ڽD��<'G*���Ǽ�5w<Ԫ��yB���j���=�
�3��<q�ּ�N����t�<��j=�,>=��V��ޓ=���=MwK��1�= ���`�=>#B�/o�3@��>W��z�vD/<bs�K��=[s&�?1�bjY=�i��o�>��J>��>?ʩ8�[��5k-=� Խ�6��'<(�=�͋<H�K�ں�=�|�=�V�<�n=
R�	G/=Ö$<]c��h�>��G=�n�=\zJ�W�w��O�<:�=LN=�����(�<&��Ƙ�M�˽���=��2�oK =ܸ4=��=���=��W>�Վ=���<$�A=|��=�W�Jeo����L����: =H�f=]�=��Ƚ.Y8=Yٽٱa<{���;k��Վ�=&�����>�1�<��%=)P_�"^\�n�ͼ�K���S�=5����B��*-�9L��=�'c=~A'�d�$��=��[�v��m-�����[�=�ӊ��C��K�w�E�d�U˽}��=
X�a=~�ֽ)3��ܱ
�-�>��C���)=7�=fo��T���f���<�P�<���)b�=���<j!��v｢��7mV�sd��e'��n�����%Ϳ���9��5#<�cǽ��q<E������D0*<���<	�=Աz��Y=��;v�e�F�=�|t��F=�(=<�L�t@=�&�<�L��$�<H>�_]=�A;8*=Ǣ=�
#��N=��n�\>��6���ۼ1R�f�L=�U\�Z�'=}b���A1=�VL��[�=ſ�<�;8�ټ�=���=I~=Q�=NY<�Z=��<��b;�>?pn<�.�=�-��2
�Z��G=n�b=�7��m���ļ��w�����<ib�=��=�jJ=�i��|>�6ܼdY�<$~�Z�ۻE?�9�E�=��$�
a��H�=���կ��m�/��S��9�>��U=Ι�<b�8=�3�<�(\��P�=��>����t�����=_��Y�"��S>)�=�ڽTx>[m��N�=�*�=�p=;{>>�+��= ��=0t�~��<#����D�\'l� K���@��;j��=���= ����E��I8��=l������=���=��=fX�=���;£=��<���r��=�,>�{�����
����Q>��d��_6��e�>��=�w���=�;=�x��d�KI=�W��{�=�#ʽ��C�}��=�J=�:=�9�=(��Ee�<���ҕ,���<���=(TV� �����=ݦE��Z�=Z�+�Zx뻨Q�<ja:�p��n��=&n
��ѽ��'��c�c�:g� ��{�=�.!����=��ؽT�,=ט=I�::>�=$��[uN=1;�=7��Ā= ��=���<ٱ���_��஽U�"=:���
<�����<Ġ���,����܎���=����E���h�/� >��X<�	F�ͳ�����<qg���9�=V��=&��=��=�j��Z��:;�<��=ؼ*>4��<�ä�ť��:��=ĭR>i�
������c"�������N4����<�eٺo��%�<& ��}Q,>6�U�_����x=���x(D<i�4O�;s�%=��9<y�{�}�=  -=����)	>�j���0�%	>�.!������%=�T�<�����wĽẽ��t$�5�P�����!��:�����=LC��U˯�|��<��	=ꋖ��8�<�F+;y�=5��<H0�=���=��7=����ؽ.��=��=�o���Ć9"k�<�3�<uU���%J=�ӄ�S���[���E�V��<ͷ�=3�>��bI>�Ϝ���$=4��p��_�=���\�6�,��=e
�{ej���=|����c��Ua=)�-=���=���<P<�=F5��3�I=���$���<�y�=��e����=� Y>$e�=�ؼoϼ��o=W�2=bN�=�#�r+U�G�@=;*�o���-�U��=��H=0��<�3��4̭=�}��V������x弶�+=.�c=���=ܒ#>TU=���ɽQ�5<�-L�!��<��>�JX=+Eؽ��=}����9>D.\�X�\��>JԽ-���l?�=�`���`f=Lu{=&��;}ZĽ����=�J��������GV���=M��96a��$*=C�#>O�+�[~=a�>1=_U<��.0>*)�4��6�=���Q�*�����Y�t�k���a�=�-�����=R ���i<j�t�k:�<�	>P���[�!��ع=*3:�0=H��=����O:��q=I�]=�꡽��>ϖ��e����=�f+�<�=0�<ŵ�=}M�<��%�	��=��s<{Ca�!詽���=b�=��#=n!=X�����=�=�=Ϫ�<i�<�n�=�+����<��]=�z���C@=!��2{>c�ż�!�9���=|e�=L��=����VμM��=[�zr=w��
��<�C����;��VR<u�'��v�;���1߂��h���2,�8�<�r���-����M�=���/�`=�BS;���<t���r�u���n���W��Ľ����J�]켆�87N
�<,==R�<�'����A��v/�q�;�uu=>"}<M㖽ёٺ���W];8��!��=��ӽ����1=f�Ӏ=��L��FX��?�.��<?Wc��:�=q9����<���� >+�t=�޺�s�8C�%��"��h�=�&��{�=}Mz=�lZ>�T�;�6���XF�X���dl�<N����J=����=Z�U=��<?EM�A�����T=ǫy��#�=-����.�<����R.��;��߂�O���Y�i����;χ�=ڦK=��ǽA�=�D۽l���F6>}l����-:��,�w��"�?=�c���������ڡ�/��<��=�y@=�p �g�����=T�����; >�֞;�E��R�><D���	t=<:�=��Ƚ+Y�=@ZI;��=�|˽�S�꒛<�ö�!㻌ǽg]T=6 =�ݬ=3��g�;s>G� ;��W=j��=�Ц���'��y���2>%.p<��{���>��=���C�?���U=k&�=��c���Ͱ�Қ����P>���M-�=N=}i�bd4=O$���=�n><qp�Y�<��$;J���Kզ�)�=T�Լu�>�M�=!��>O�=�Ō��5>sp��@彖� ��0㽓I<���==�<��N�<p����ri�Jc�<bxm���k=6=钽����<!�����Թ=t�����,<�J �(!$��B���<ؼb�(=g3�=�>6����(����:=Pv�=U�
=
�$�ȩK=���=q0w=9������7�<�(��A���s��m�:�>����>��%�Ỡ��'�7=��h=�p���DŽHG�=�`�=�h�=hT>dQ>�-�=�}*=��=�l7<昽]��=��8��>߬}�<.S���=8x���Y�<���<��<L#����;�q�������xy�̌ >�.e��?��K�]��L��l�=y܂=7��=r�=E`��(�}�����>z�?=׳���Q��
�Q<�ҽ�d�=j�u=�Ľ�jr=�U����<r�<���ĽqH&�xz�=W����0��ϒ�0��<��h��="����й���a='W�=�y�=�65�e�=��h=�=�f�=5����K�6>���4U=��½4����$>�<R�=�S>��4��2C<����j�v����7T��}�<GG��M��;�!������Z������ូ}��=9�>&���A.�nކ����=���=ߜ����=�};=ת��̽~=�V����=3��'��=g�ߺ������=�p>��=_L���3�=��˼C�p���=�1�����#v=��@�槮=��=�⥽�Խ��SR�q�ռ��b����= ���=��<�Ƹ=��~=���]��>�=&>c)�=���=��.�͛���Z���Ѷ�/�l=��ܽ�浼b��;��=8h���*=;U��.7=4k��t���x<!2U���:��>�>=���[�����0��c�3�m�<9@�=$�e=��߻ȇ�����<��Y=��==�=�y�<��P������$�
:��c��:Y�=�䋽�[ͼ �=��>;_e=��g=�Ѕ=��(<al�%L�W���,��=�;�c�Kऻ�|�<��L��4 ��)U���p=�͓�H�����\潿[�<I6=�����=�H=QV�<�W��WE=H���;=���:�ư=�WU���;�	*�|nֽ�=��n<�w� �=�b~��vB=�h�;@�<Kd!>���=0��"cA���;^QI<��=�q;=��M=* ��P?i7�l�����=�~�='�(f��Uъ�̤����G�;=���=�>lJ�3p�=oUҼ� <���=��M���_7v���N��ߊ�ek�=w6U=�y ��L�������J��9���%<]g0�`����'V�@v/�_�A��-\=�!��#��<"�����^y����Q>H��;��=�m�=`ŷ;J �=2����'Ӽ�l�=R��=_C����<6�<�z�K�����=nA���٨<�Y��Z�%=�d��c
>2ԩ<��:����<L	�=pp���q�����=t�<Aũ=���m,��Y��Lu���?���Խ�㢼�>Ƚ5LW�����ɋ˽=��&�����=��w=܊�=x�&>��9���2=�] >�e��=W�\���<k�h<���=��U��xj=��$��]��R�����b=%��#�=�2<x4�<][ѽi�����=�'�}A&���==�@�<i���c��6e��P��,��/ ��EAp<ĳ:Z)�| >�4>�z
�DS=��w=9��=�h�=��0�� �Gz�<��*����=�Fڽ������=���<M��,��=�2�=���=">��5�OH�$�=�O=�˽3����W��q�����++�=��<@������=�
�=�!�=K />�:�f*���>�ʅ���=��!����=c%>?=͂*=��>� =n!��4�KʽA�<���E�W��EH���"<""�>a��Z�=�˼=�\���=BLM�n�=p�z��s���1C�8O��K�=�~B�:�n��g>���<�v<>�&��	h>�TX=|���鍼�Ҥ�E�ǽO��=����y�W�-a%>�>�k���<Ƅ.�1ܣ�_��<"��=y�P<�Z�=F����E=��=�J9<�1S� ����]>4,)�tI��?�����a=���:H}�=R�zx������;'��Xѻ;{�v<
o�<�r=��=��0W�ڥ���<��_=S|=+�Y<���=�<(o��V>˃<�Î�7&W=w�J��,K=}�I���%;d���� ��>�~>��<S۽.?=�R=G2��c=+q�=�*d<�>O��kZ=��ؽV�n���">3�ɻ���=�=��Խ�c|=��=����xg=� �=�8=c���#�;@e�<��1���`����=�Ξ<��=��(J¼]섽夙�����!:>�*=f6�<�>��7�=c��=��=?ƽ2ON<�=�yֽ�,">d.=��=�!>����З=^C���Jʼݼ/���ἦ/M=s�=��R~��֕��>���B2=<�>-q�=	�=_�= ��m���f��H�=�bw�1�=�<�b���Ei3=N�=z���#��==�W:��(�n_>&�b<UM=�L�=��>��<Ħ=_E�ż���f;���b��0�ۿ;z�H=��ѽ�r<g����~<ܼ�=嵏�U�ڽĐ�<��ϼ�����e;4�=X�/��|�;�	�VQ�=��8	�J=+� �;�!mG=Ґ��Ҫ����='�;;[�����T`�=+;w������=	�=-�齛ȧ�La齃A=@6>αe=D��������<����)���2>�x�=�Z> ڼ�C���.>�u�v� �^��=�2�;��[��'�#x��u�F=3ہ���R�,��=������R�Q�U�h�������xs=ց�=�+��6���8�M=q��<d��K*��Lk�A�[=��w=?џ����e���»O�-=����{8
=���L�,�Ͻ�g�;Կ=?q�>5�z<$c����'�i�Z=��<���=�6r<Õ1��V
>�w�<�����p<;R��0�1����I���V=��s��5��������u�e�7���_�<�ݡ=��<�V��d��=��><�]�"�V�K�'<|�r>�7<;�*�r��=-��:��`������j���V�cڝ=�{�=�D�;��=��
��ŧ���=���w��<��<�r*��4>�&�=K�u��;�}��=\ =)P5<�����:=g��ۭ���鼛ϻw��=]Z&=� �<<�U��j�<~��������W�E>����O��NR��A��'d=c�=�^�+(Q��j�;6R�=e��[4���=�}ļB�����Ľ�Cֽ���=�{=(OP�&���<C�8��<��3�6�M=��I�״Ƚ���<Piߺ�_��.u@�e=\�1=FF=F�; A�=�����4>�4>����۳���ϙ���͆����=&�=�%�ɠ�<�6�A�=+S5>��м+�c=��<2" >��>��>-8�%zջ�yӽ=�y.��9<<��P=z��<��<�ɂ�~=d���	o;V��=*y>�3�;���=��<՞B���t��I=�r=&"_=1�=���*f;�H=`k�<K�Y=`��<�恽]U�=���<�}=y׶������=�K='�<D+۽�<>}5=���=P ����<�Y�pP��q�<(7=�[��,�V>Z�=���ԻL�*���$�=}��<��߽$@�=�c� �ʻ���41�,/���%=.����<z�����<��
�f��<iD��5m�;�ꓽ�S7�<<���^N=����_��z��=�=	��;U�#>�\/���<��:>�+�<����a=3C]�7���W.���1�'%c�/�ɽV�~Aļ�\y�d_�=����og���'��T>kų=���}���	����!�>/]�<NZ"��>>~��=]}E����<ɴ�=��=9������Y>�Xu�Zf�������&��_�=�),��£;Q�>��=�ٮ=���<fUl=K�=U��=0��tv+<�놽�E�V�=�.����c���Ǽ�8�= ̀��ӽ������ڼWP�1B�@BZ=<S|�3���MǼ1��=l 5��0���ӽH7�= F�Ka�=U�x���I=������4J{�|Ά=�
�U>�If=/�T=�i(���5�w=`0��?�=Xka�EW�<��x=���*������E��}�=��A=�=�D�=W(Խ`�=ٹ=�6���}��;|���y<����*��*����J�=��=��}<. ����<������'X>w���+�<@y�=7�i�]�|�'=�8=R%��2g=B!,=)�=ßE>�Ƃ�'}�=�>N/�=��=�U8���=�u�=�f�=���<��ڼ���;�"����A��^�<mH�����=fۮ�Da2=K�{=0�ǻY=����ºh�<(hH�9;>t�齝��e��`�;��=��0W=�%H����<{��<؇�=�6<vO=�7����=d�1�$�� ���$/����=%_��D6��9=����c=�����t���+�=��=�� >Ê��1�P=m�b���L�;n�<&O=+�>�*>��Z��[�{�=����-=t����=/��=�Q�j�
=���<�+�������=<(��Qߗ����=��F�2=Z�<8�<lxʽϨ��H=qR��`Ի�L���2��"5>�0�=��M�=<����n�ͼV1��Xt������=t�/=yY<3���		���=�߼=�e��g��E���<�g7=S��=�6���=Q���i(>���=��<�u<�b>��<�(=���=�8>�=��5���	>����&8=w����=C�>8Խ�!�=�����i�<9�=�����U�=���ZF=�����<�����<��B=x���(�⢜=/�)�>�$>�$�ow=��>=��<��/�񲇽f�;���fY��f�$��T=S��='hǽx�_��j>�t�<���<�X���F��2�w���3=s��b��=w�h=�v >������s�o� ��=�>k��%�="���~ٔ�~�;=��=E�J�1�P����=۶p��>�J����4�W�ѻd����<4��M�=�=b�e��=7	�<���;�9>(�m=����x��=��>�}s�� =�B�U˜��j[>򕎽l�̽��`9>1 �<O�-=�+Ľ+���(>N]��5j$�u.���=��C�*��;h7&�!�ür�>>�!5>�xW��3�=��m;�R��m#=�=�N<�uu��q�=�**��M���0���fZ��}���<��+�[/L<��T���l�񥌼hk/=Ģ
=xP)�˼=9��=t�;=v�ܹ��>�͓=��<�x�=�)=�OI=Z��;���;$�o=9p'�M�<��_�0n-��L�G��=�B��M�<��6�G.���<�D(�}�9��q`<�9��*��<���=M�:��'=�f�=]K�=C�<>���]��%��U�-=b�=:�I=5'>��i= �=�̼�A=a,�B-�=�+�=��=�56�MKZ�]<i�)���,�;M!�=�f�u&=W��=/=��=�<,�<7i����=�~�<1�=�4Y=�2h=_j3=Tf��ٖ�ձ��|M�<J��s�=���<�_���S���?:� _�=�>f�&=�"��Pȼ������:!9/�H��𩤽:(��� �Lܽ��b�#Q��s��:��=ŉ6�O>�=�i<���=g�ݻXν�M:>
����)d<��3>��g=�{�=%HƼT�=rX�� �(>���=���=��꺭B=BcĽA{½���<��=X��������-�=� ����=�������9�o=,�ֻ���=���`�>�==}��ܵ�r'�ŗ(����=p��9
�ur��.��m���E���1�KD�<�_��)���bF���;�\��h�����=�
���w!<�M=�W�a��=*�l=����r��N-�FF ��+ٻÙ="�t=���RL�yM�=�$;���>5�<i��=,a�<�ը=���Tᏽġ�9�=q��<I�?=6|=���n)�<�K0�r:=`�a=Z�l<�N��N����]=� ��Z΁�ЅK=�����r�=������qSI�G��<�I =e�=�̌�hw��{�$=N��<�.�d�u=�</s�=���<N��=6��:����||�=�D� |�=��x�Q�P��u��UＰ-�<J�̽B�����=��������Bj<q<����=u��c
�;��<j�N��P%=�=D��u�j����=�x=���W4=�<E�E\��k=q��7���!������Qq=�1=	�5;��=��=�f�<[��=X
��A%� �|��=r�$=pj�=&.=0&0�6�Y,��ҝ=y�<uY�<�t5��|ؼā���%
>,������=t�Q=���:�Ӽh�R�=|�>�qսˈ�=]?��-C.���<g�=��>�\�=Bb���#�<�z=�8>�)���=�ط=��C<�"�=�<��A>o����&?���̔=���B�=.��I��=� c��>�����;{Z�<O�.�:]F�>U	=>�@�����R��� >w�;����gY=! �=��<�	5<��">�$=����z�����<���D�=̖�=��o�q�Z�'��҂�M�E��p>��:Dz���{J�B3�t�����=V{�<��F=���=���l�4V�=�z�=� �a<�V�=�����(��� ����#�X�<=���= G�=p��<�6���'�*r�=�:�=��=rwc�c����x�<��=��ʽB����]=��>�=7R��yW=�5�@��g��U7>�5�=�<н*� >̡>�^s=��1�_e�Y�~�kf}=i�=i�ƽ����[�2��W=듽K��u�|=�h����	=��ԻD�:=>8+�����>	h�=���%�}Њ<��=KO=��ѽCaB���=�y"��2����a=�K=N�=����s��Z6��ܧU=��=r>h>�O >�l;�텽E��=,1��(/��i(�9*�=r(Ľ���<ST)�R��=}�D=���<�_�=?e�;�LS=ط'>�V7�̡���Ӽ���_��=�)�,���Ͱ�t\Z=�݃=�Ց����<6�=ߚF=�\r�����3	��P��I�F�CĿ=���=����OP>p���l\1>V�:)^O�);�=�����M���F�=~�1�<��<��*r��qN0���&�4Ƭ=R >ޟ��rf4=��=���=>m��8@=�J̽q�Z�N�;�J4�9ӌ=�|�=�����60����=�	��Ľ���<`����s4=*��;�qC���=��3��6�=W��<�H�>��=�J�:��^=���=���=9�U=�ؚ����s�=���c@��嬇���8>�ŽOP<c�)�=��=bx���B=�1�<�@�=b��<b����ҽ��<-�v�v��vx�O�<�چ�u�M<{��=�g>̂̽�A�=H���.u��i�=껼=X{=^�Ͻ!\<S{(�Y��<�>^ڽ<���+|�����<�IU=���wZ���k[:z6�=�X=X )����=uE�<.u>��J��Z�<w�ȽK�'��29�<���r<��v1�Z"�����=��"=Z?���:�=~�����S��[#}�����H�=�w��Ƅ<�W�=���	�@=
D4=�~�=�WD�PZ�=���=�%��c��.��;m|�=pl��_t �����ؽE3*��%"���<�:ֽ�>�}�8�!>�V�=�SI=b
e=B<�N��~�=]]��6��:q���=��+=#ûƣI�y�=3�=��(>7���Oh=Ú��)������=wm��F���&=eU½9��=�>�N<���=2¦������	�8�<=��J=­r��m�=nC�=��V<��$��d���99=j*=Ηƻ��
�*I>NF�o�e��w�=58
�Lq�<�.p=�� ��]�=\�m=,��=��<�Kv꽆-�<�M�ja��_=1i�����<��=D�l=�
ɻ�)<�i�=�]�|]����<��Y=O<�i�<�K�<� �A�>���-���;�|<�H򽃳ؽN�E=e]���2<X좽�=�a1<���=�'����=��-���;y|�=�i�<�6ȼCD�%����Z-[��{���,��!�-��=�[���������=kLW��%�<ݕ��D;{�:��U<[����=v�7�2wX<&N�F
�=�y��5��r�>z�G�W��������W>:��=>�1��v��*Ὀ�=6M=�8<��ü�7�v_�;��=�gü�E��3:N�W=
�=h��=�E��g	�u�a��b=����X��Q�q�B>E��=H8���1�=��=RPN<SR���uL>�>�]=��9>�ʅ��A@<c�=��;�C���>;f�n{>�v&�j�<?�=���<θ�<�`3=E�x󲽊 %>l�~<^���ś����=�m��"y��B˽!Jν�A�=�U�<�;I��d>K�=��Z>�G���̻��=�A�<a�4>��T��n�=�=h�&����=`7	���4���=���ǰ��W�0;i¹;ޑ�<���=;>��<L=y|>���cȯ��-ּh�x���F>��ɼ��I=;:���/=��� ��mV<Jb�=c�����ٽ(�ͽ�1�<B@����=n��<�>�f�>��ݼz��z#>���=h�J������,��qJ=�8���%>�_=�y������5!��$Q���C���>���;��S�х�;{��=������=p��q=m0����<�R>Y�G� �ս�����= �=�x�=NM�*F�=?ޔ��-=P}0�tj�<�o{�q"�= �һ���x<����� �׉ʽ�����;/��.=i�>5&>܂q<�����ʇ=�G9=��<ft�<x��:Q�#>A�o��q���ܽ(���<Q�<�۽��
>��=�!=���<�S�B��<s}�=6F߼�Ly��浽�I�J�V=G:�=�`�t^=�ˆ�=��ҽ��`�.��D�f�"eٽH�k��t=E'���ͻx�0�Hᏼǥ@�"���������;�=Ľ���<?�;1��Q=˽>q��<���<�}�� �6=��	=.��=b��=ѬԽ����$�X���̨���%���ie�<��q=*(�<��=I���α�삥�H=l����g�>ab��c�������K=i�Fck�ۛ3������-=�tI=	aI�:�=�K<����=۠�=-`=�8�>�=u��߁;�@��< �+���v=8�ټ��c�@�E�ꛙ=L��,`����#����P4��fI�cRZ���K=�>f�h�-�h��:�=5<�=��ڽ%�=�y�hh�=�-�<JN1�w�n�y���I �5�$=�2�<,�=~�ýzT�=�`ļ���=�����;����=����
>$.ϼ�`غ�X�=��{�� �=^�\<|��;��R�|�k;��R������<��+��K�o���Ѽ�b�=�=�j}�m�
=����)��,�mw6={wI��u�����<�x��v��<�g��Y�����=qI<�{۽ٸc��ѻT��<+߽*C���=��<��<�����E��߅=��?�Н=�f^�Q6����=�E
��/>����t�<b��;���=b�R>��d��j����[���J��>��=�`#=�5�<���<4�{=2'������I�=7	���E�>2Kɻ�j��=ع��Pa
>�[$<��"��c���U�=�\��@�6�h1�=��;�WP>q�~�F���=���煾jG�Z]��`��[��=����Xr=I���*��'�rt�<3$J=X�ܻ�t彙��<QE7=�.>I]:i�U=��&>%���&Ng=@�N�ԫ=F�h�һ>ȏ�=3qm<^ַ=#�̼���<����枤�j��;s�= =��:�;f����F=����x1���=���;g^�9��*��U�=j~��G<-�M��Y�=^����	��I�=ɪY�'��=6=*<L�=5�=��l�)j�=/u�=_JH<B\<%M=؈�������h=ݠA=Y�4<��˽ s?�|�=�'�#\	="�#=���<���[�=�2��.��S���q���b=�$>>�)��63� Q,�i���6���e�ޑ�=�@�#��������<��G=߽�#-�)ʣ�^������'N<��l�$5���W�$	=^�=�(<m�=���������a�@;.����l�=���������=(73:�Xi=I�Y��b3=��$=�8r��O�<�	{<1��=Q�=T��*��<��3���>�H{����I�f�fӴ=���=9�=9^�<?C=�Ÿ��<'��;�T]=io�=��ۼ�>�=ʉI:�G����:�Β��Kd=�x�ui=�����=��l<�.>�q��f*R=��[<m��=/c�=[�
J<:0�Ss]<�tt=�S�����=��k����=���=w��c	V��Ђ���<�p��г��>��b�K>�ȅ��꙼�}�������<i��=�3ż40��=�
��>�Az=LI�<,.=�I�=I��<\��;k�/�;̽8m�hA>��=,#�H�T>�95��2�=�O�<fuͽ���;R����
={�7��1D����~��ׄ7=Ԫ�=��۽���=W��=�鶽�ܼ��c=]['>�L;���4��<=c���1=ue���=��:��?*��<��d=��y%���Z_<�:����]��������=�>�
�clY��2��=2��g{<�K��8=�5=^+����<EƁ����=��:��c=B��=�n�=p�r�,��=�y�=Ꝯ��z$>ū-����=�F�<�ا=��=G��i���:�=���l��;b�����BM�����c �<d=b�>Tu$<섔<6 =�o=���P�<�T�2>�$>B=	]1=G��#�X�ϑ=��y=����=r�=�ܐ<+W="�;�0rû�:B=��^��ִ�8T�]�A=�v-�]"���S�=H5�<����d�=�B�6��W�����=�<�*�M�)��M��i=�?��D�d<ܥ���P=��ٺI�½XW>�j>��3� #ͼ^ͽ�!����#$ ���=(R��v�-���ս����k�u��ɨ=r�V�xM��]��>�����=A��)�=��;��w=�ȟ�4&)���ƻ���<�<Y��:=+"��x�<�j�<�nl�W�<QΝ�$�!��->D��=y���|�v��<���<*'w=�-½�t���j�<��<���=;rW;!��Qou�M�>S�E��yP=י
<ox>�n��m��<�⭺p��	��=>:	=��Q='+��v�>�����=�����7=��=�I���ۼ_i�<���c�~���l�ktq=崅<T�=9.��\��$g�:>��=��n�V
|=���=a�;y��4�T=br�<v�>������A=�S�S��;��;��=1�3=�#f�r��=D�X������}=@�=do�=0�%>����=�F��.\W�&��<� v�`���;`'>p�=�����������
�~������I�=�I�="�ʽ�Y�<��d�X�D=�HS��&h���6=��ٽ��=A�>凢���=z��D�s=1�D���,<A�>�����>�8I��B�������;=��=�g����=}� >i<:��&ս�l}2=��;P��>����r��=�=�q`t��O�=-3�ˑx=<�_��<�x <P$��b�1�������!>}��=��;�#��Ƿ<�Iν��8=5�K�����,n=t��=@ȯ��K�����o�nyD��"A=�w���Q���ʤ�<�<󘽷���jރ=��g>�?�<D�����;���@�<m)������s=��<�=wt><�4��S�-.��Q]��s��������,�)B�<�&>�Ү���i=�����=$��=v=��;Zـ=l�>�$�U=��<�R� ��=	�W=������=�6�����k���[>FU��̄X���/>}�;�ѕ�w�z<9Gr=R�Q�N}=7
��a� ��<f䅽��	1�v+R>�0>��=�@=t|�<im����}=��<vw�<b�>�����&=�q���&=�Z;=t�	;�赹��<<:ּ']o���wB�=�5F�X��=�4z<6hd�e�:W(��}��n;/�
<zO��v��=E4���=؄O<��ͽ��O�����;�3�=5���"2���kڽc2=����s���b��y�=H�=*]��>� =G���̊�Y�~=��&��s�=���=G�4���>�_=�
�!���� =xz�=#&��[�=���<�ˍ��K=wz�:^�	��X������Z��=�ٽ(�����:we�/G=j���<�>=�;>�"d�ԭ�<4�8=��=�<���<Xx����=��0�]�F��e�=ʕ̽��'�ɥ*=�l<.�����c=K�Q����<t��� ;����Ж=˸,<��5����&��=Y(�;��=oq=�×=��Y����<M�<��ϼ	V>8��5y�'�>���=�f\>xX:��E�����=aP�={�=[�=��Q=7�	=d�=>�C=������=��>�'�<'�󼭜k��h1:�ۃ=�7�<�><t��6�.�K!���>�=�7�<޾,=~*�;�cV= �:��w=dn;�[aʽ)�����=ex=�B(=>���m�=)T#=���=��=���<ׁ�@��=�*�=��X<�<T���}=�5Q=�Ї=�ه=���5��=��o=_?���b㼊�>kǺA���1�L��Š�̸X>�a����<�v��}���>��=&�'>������=��=Y[�'<�Ӂ�A��=�潡4�=�<�a�JO
��]�<�;=�0�
=|<?�>��=�����8���=���o@�e���*aB����Ƶ���μ�Vb�wM�=J�>h�;K��=e�=Ta>PK>�y��W�=^q�=�1=\�<W3ۼ[����T��KF��R�����z';��k޽��#�pR�0{���d���u�7���\�=��N=	8�p��f���)��t��t#���G�	��=`�#>G��)�\=8��;".�=c�煽�1��&uW:�Pսu��<=.ֽa&��ef�;��=V=���t�=[;=�Br�#B>�r�=�s�`�=���=Ju��6��Oc�����&���V=��r=ukM=�G;;�������<�Ǽ�lE<�8��Ƚ��>�`3�DA�<�7!=H+(=��|$���>���=�b="�B=CRY=t���<=�B;YUr��	&=,����>g���?�=<@�g���ؼCLν�d�=tH=�E�}m_=~e��b�=
0�9���g�=����4��l�g<�>��=�v��c��=ݖ��
�<u�^>a� =*�@=��i�9�=�;�,�=�,�8�S=Ǔ4����=@&��G��<x�>�����Z=%�9�Lx!�<>(,���(>W?2>�,���=7=�u+��J=�2.=�	)=6#���9=�E����q�{��=7ὠ�=D}b<�+�=tş<	�l�a��<�=�=hی�2��GJ>T��=���=Fz�3�D����<�6��D�����~�=�\�=*�<;_�n<�4~�Y([>C�[;�y�=���=��y�(ռN㔽�q(=�/���a�z����g���K�q���0�=�xs=@p=��+>X�@=�ʽ�F�<B����6=�g��[A��տ�=�&�=B3��v�
=]C�=����m=�[�7�5=�'Q��N��u�ý
L��z�ʽ�=�WM��ŽNk��#c��k�3>�$G���<"�߽��N=Ԏ<ڨ)<� z��e���E�S�1�)޽C��=��/�f�b<�Ņ�e-�����=�"�AB��
 �=1���Ҿ=��ӼPׅ<����'?=+i���6�:�M>+�->��<jԠ�_`%�|�<���������G����=bl��>�<�$+=q�=�0���1���<Pd��޹=-{��S�	>����(����,"��e��X��`�=��A=.x=��8���F�:��=@�����$=1_=�W�=���;��.��-	=r��=j�)�Pl<1l�<�&�=8��,=;_��<m�<����A=wy�=d3d���H�|_
>�%�(�J�b��;���=@ݼ�1�=�H=��>c��A�1����y�<���MZ�}<��r=�#��*��'��D�=�/�<<.�tf�=�L�=4%=�>u�x=�����=��5=Kϼ��5�=}�>�'w=�N�7;��Zk��O�;�����<�N0>�7��}��_`�<���<�Uw��~��sY+=a>`_ɼ}�z�c/�G�ٽ�2��A�Q�H�=��=��a�2�C<��=w>�d�=��N� �w=�o$=�:>羽=8�K��H�:/n�=��<� ��r���#$>�|�=p�<��r���Ƚ�ݶ;)鐽��v=�}Z=B�L�t=	z����=�>׃;۬��DK�=���`׼7�N�u8��$.��>s彞���Py��2ѻLxf��=�H>J�F=��<]��,҄<"Ƚ�U<�'<�T�=u�`���<[;=�@�=����o���<�)���;>���&6��O�$= ��<5���.�;3d�=��+>} a����6BI<�?��>\��N�=�t=M����g=>��>�L��1y���=�u�<ӽ�-�l<l���o=�{�J�=�M�<��<ॽ-�>r����=C�=`�<������3=�cr����=lnz�������<�#'��� ������J����=��ӼGQ��u<�3�<S��@��;�d;��Hq���ռG�����=��$�C���=�����;�_=Jٽ�v�=��h=Шؽ��=�C�;�ʽ��'����=�L���=�(H��5T=YQ����=�ꞽ�At�)���#�z�:�<��������<t;���[@�௼=Mz<�_@��~�A>����<�Ƚ;�R�=��)>*$��U_=5Ґ:Z�N;���<��+��=:=��?W=�=��	=��Q����>�l=�w<�ۯ=��!��Z
�<N��=���Wg%����=B�==�����;0=4��H��mʼ��T�<�ڽs��Uf=��<Z\(<����8��=�n�
k=�R�<7cx�X�=n{?�^�=.������$&R�}6����r�mn�� ��F��=M�=In[<1bG�d{��y��;�q���>8m����Z�>�=h|�=rV�ɽ�U�ý}ᙼ⎣<��q=�u>��X��,��!h��ӱ=m B�3����;G��k�t�&���u^=�\�����;.R_��Y8=���u���&�\��c���~!=6�Z=��?=���=(��ß�=�>�o������tļh�2>uyN����v����=\H�<��=�h�9=��=�6\���8>7!��\Zc����<=2�=+�3��a����=3ǽ,wݽx2�Q0˽��>���Y�4�N;���:7���Pŋ���C�W>����0,�Zj)=�C�Vb>��>��"��^�='��=���<NF��[��;�<n=�9�N�W=�w&�Е8=�G��{����;=�;N���Y>�XM��K����<Sk�=�>���+=�X�<���rr�94��]"�T�ļ��b����ny����=o����ؽ�h�<��λOD�!a�=�ǽ1�]�  ��=��9>`=�=�G�;�#�=q���=[f�=SK7=��S=�ֻ��=��=�&�<�����=/��^A>w��=[uJ=���<N��AE�<�����H=2$8�O��H=>�-�r?!>�l<~�/���=!AֽǼ�=z�<C��u����T�=4 >�`*�<k=�d�E'�g��9z���ߦ=
DԽ�^�=.�=Ț>�w�=���}�<>ܠ=庘=��Wz�Ʉ�=wW�K�=K��R��<����/)���>�ȼ�]�=��\�i����"޷<_"�@r=-1ߺ�#�=l8)�u�Y�� ��SH�<��Ƚ��<o�<*�D�U�½)Y޽>�=cM�<�u�=�݉=*/q��q���3<�US��J�=���=�����?R=��L-�F�>���	�ʅ=�ɴ߽Eh=%��p�O=�i8�D�0>O�I��e�<;N: � =��e=`�]��D�=٧�=WL�;$�=�q%�����ּw2����9����<m�����ㆽկ�=Lu?>"?ݼ;%X�oO�BSb>r\��2�#�^�L�� ��O��J{�G�=T �<�����=>�L���˼��I��뉽#p�A�'>S�=F��=����+;���I��>�zZ=��<���<^c�;Ց@=�]�<��;��=d� ����I�Z.j=����/>c�G�JSo<�0= ���Z���/ֽF(<d���yk�U;����S�?>x������<�G��P>5H��~7=��>�
j�� >7�=:=��H6^=-��y�_;f�<�j���R6�tG�Hz!�Q����=Т�=1�7=t�<�c=5p`��༭Y�,X,����=��Ͻ�L�=��>h��;>�C���y�?f)��dV���D<C��T�=�{<S�����^=�l�����=�?��6�=�`ͽ��#����=;E�<J�����4h�0�n<2o.�E�<籷=@�q=�U�ImI�#�X�P�"=��=*��Ǥ���;��y=k8����_���F=y*�<��y=���=��=��v=��=G,�=�=��=-��j���=�=q��B�����O�<>�\�<�{�&i��9~�ד�<F��<���=�E�=j�=�-�����<�r�<�5'�\�Ӽ���<�C,��T=�ǽ7��=��W;6S&=��;�X�0\q=v*>�[��dpL=��o�2ڲ��1���1�����pv)=)�d�w<�b�q`����{���AB��/E=c��Z��V*<��Y>���i2=|�=�ل=U�<��<�"+��K�=�c#>E7���o<�D*�	л�W=y��ա�?�.=FcA�����>*J=+Ϣ=�������=�`=�b���<7�6���=�e<>��Z=��@����<���<��<��M��-�+��=�U���X�=l����i�=���=���=�����s�e�C:���=m}�S⋼+I�<@�=����=�m<=�f�<(n�<�l�=�����<�$�\��>"Љ���ۼќ=��:��3���w�<�mN>��?��{>����c$<����f��	��>Z�0�#=�?=�돽r�o������8�N���/��܉=��7�}v�=N�=�9�:$�������|�H9�������=4��;�>�=4>IF����L,��Ƽ��=���<G�4��=ޠL���>=��=F4>EEw�M�����8S�=Uu��\d�����=���)z�=Q>T� �@*>"���28�>Q���/�=��S��d4=�Rq���(>���=�m�<Fb�0�
=��=����X�=���|�ʻ9��=RIS��*����=P�(=l�!`�=�C�=����	���DU��=I�=¯R�-�<����r��=���]�?=o�=�%�Θ=���=7�l��[��«��UU=��9̖���0�(QZ=�?�=U�(>U���@����A��G>���:l=���x��<0I�C��`�ٽ/�O�_=&.>��Y;xp��7�=��X<��=Uu��Nfd=T瓺�_�=i��=ű��}�＀��<���3�e�sR=���/�z�4t-��%<�љ�jG¼��V=��g=AF�-�н6�Ѽ{i�=��D<g�:ތ=+��>x�彇��=�=���<�z�=�@�k�,�K�=c7W��3��|�=��-=r�4=�U�kH*=nu=K�=p=Ž��n<˹�@뜽��{�Ɖ��Q�<S�=I�>V>�Fq��I l;L��;�9���=��Ǽ�'���h�iJ�H򉽥J�=]j>s�ǽO��xs�;�Ӏ�F���@e��;�Lm�=Ң���H�=~'>��(=}��;;.Ͻʆ� ��<�Y�<���=���=V�={�J�[,@�H���<�M���.��,�<���=�t=�!��?L�<
�2��;h���ݽ>�Z�N�ν���=�G��i�9S�>���=�i���d�<���&�=�IV��l�<+)?=�ǌ;�u<kx��h����=j�����<fBL�����V��~�ԻOY����K=���;J>Q��<��������eٰ<�^����Y=�v��i�ƽ�M_�]���<6=�w�;�#Ļ�];
�༰�,=T�=	[m=b��=�Q*>Ƭ[=���=4�m��5�Z�=��7��(��K�>��J�=�圽�׬����C\ɽ~n��C㽮]ü��1�".�<.�<���=e1����=�U=�����.>ZƄ==�:�=�v=lߧ��Jѽ��$�(4�K�=�<3XS=�� =��=��=B�V�r=�=���ϩ-<���u���=Z9�=o��;b��=#�I>}�>K���¸�=w��=/����=9~j;qe�8�6�a�Ӽ�`�
��u
ս��T;��<�(B�FD7�"�=�N�<@�ιI�������3>G<����xս�7!="�1�⩄='�h=�?�=���J��\n�;�[����;i�=�����v�<�������<7�b���?��7⻕Aټ���`��l���7o��"�=xꖽԶK�w�j�\y�=M!=��f=��=l�*�gO-<H�=�=Yܻ���b�<Q���=�F�<q��=5E�]�ݼ���=3�P��l�<F8>�$�=-��^��{��U�<�&�t3�<h�|��aj�K���ʉ<񡍼L|)���L����<ь�=#�">���<��<_\=U�=�2ʘ�N��=KW�=���<�e��Ɂ�f�>�C��ɋ�=�7v�
�u=�:�=���=y
�=F����5=���=�ⲻ�ƽ!QK��h3=�B=�[�=�=Ž#3�=��a=/A)���=8����=~{��^x=Q,3��.�<!p�=�g=<d�=�����d	�~35��X�2������=�D?�[��<�Y�<v;�E$>��]�<�����c;M+:���<I�+�XF<|a�^�ཾ�8>&�}�v0l=PhT�G��<"۾���q������W���>b�=q� ;�'=�����5=��$�c|��k{��J���2������R{�=x�,�.��-����=4=�s =��<�E��:�; �q=���=�_���7�<���y!|�&������WZ�`�l$p��@T=#�&<�ᑽ��;�2Kw<�}h�r��=p�k/�=]ٻ=QzD�3=�f���<�w�V�=)
�=[P\���ѽ���!熽v�=h�?>G��=���<k�V�����zE=��<���)���c=�e�=�р�ko<V  ;Q��<��=.M�<'��<�P��m%]�o𙽐jM�㡢; Ni�K6n����=v��ԗ<�J�<'7�gd<-I�&��<�8��[��˄=�A�>{J3����=޿=)mW>U���~ ��I=�PP�x�%>����~2='䕽Ǿw���=cp=j3�=A��
��v���۽���<��<_8=�{c��{�=y��Au��q��fx=C����>{<R��h����=ޠ�<�ă=:,���)*���==��<��H>x�=�$ =0���F�3�>e�_?�<���= /J<Ý>�O��f�=p<=�7=�'<T�D=�={M����=�����<^&����2�<ө�=౽�M�P^��m>ѓ\=I�<��U �W������
���z��f�<A�=��a��U�?=[�<>�ڽS��=��@=�����<�P�=E���5L=�i�?q<g�>�l�����	�Ͻ��C���=�m���ws=�,=<ԩ=��^��
�|/?=����=w*&=n��<t��=�x�#d�9>�=�C��������S�=�XQ�7�|��_�<���<q�(�@}�<P�=�c=�x��iW=\���x�x=>��0c��S	���c<�<�y]���=�v>/�=x�h��ֵ�L:=7��<�Z*���h>�0�E)�=u��=]z���O=�f�=�x<��=4�=��<)��}�	=�rؽ��;­,��7�;��vP	���һ7�=�gg��Z����ؼ�=�=���P��.'1����=�>���$<�$���<��U=��e�wX�=@^꼠QF�)���"�=�mN=��<����SM�=���=�E��+!�=��4>���;(�=�;�V�=��u�����=���������4����=,ܰ�yn�� �> �Լ��B��i�=��=�
9�iz|=h�<��ִ���= wI;�:|;�l-�LY=��>5���ۗ����=�d
=p�=2p�=��y�5�O����1�c��\�=w���c��=3���ή�=K���ɡ��\�=�c]�)~�<]����}�	��=-f=VI�<;?�<X>�����rŎ�i�������h�q��>P$;�|���w��Ͻ��=��3>c\S��c=YR<�X>�U�=�+&�����b7��;������VV�=�t�=0�˽�Y=:l��w��q�#��gN<��v�>0���h�=���	�=|���%	=�I����<�۽�q�=��B=���;W<6;Z�=�J�!&#�A���) ���N�<>f޽�ri=tym=ؾ������?��S��<Ԕ�="=)	R<x/��|�#>��<d�=�]����=�^=`E��z��=I�G>YQ� �= �<ǆK�'�>W��=.�>u��-����=�b=�ŽԊ<�w�x^��9�>`�>J(�=��Ѽ0�G��7�����h�=��b=����->/�=c�=>����d��ZY��"�L=�6��Cm���NC���=��=�s�=#�<���e�;'KF>��=�|�<�03�V؏��\�R�M=�h8<sq����t<l4�=�
{=)�黊nu���>�,X�� u�3vY<�����>�0�=�ĵ�j��=��=W��=�_���$��(ǧ<<浽ڑ�=��˽8�"�`��������k�7��v=)1�����<�^��e�;�	�=�l=��p�T'�=N(�>5>���S8�<��û.�.�6�=�X��� =hpH= )=�4a�S][�^zY��$��o�f=m�����佯�b<w�{��;��=ѓ'=d�^�J6�=���9���R����<%@�=���t'�<����r�=��B=*ܼr�ɼ�~m=� �=Pm�=�<������b�">�f �;u(<�b=��9<x:�=9���Ѐ<+��]�=��������P�]�_�҃�;<�|=�E,<��!>��=��=�"=����>��9=��
=+�0>�;��R>=�K�)P�;�g�=n��=@%�o���ʲ�9� ���0=������n�z��1
<�6P=<�d���>�Rr�zC��fd��t���>cK���7��j�H<~X��v�*��ؼ�/=��=>|�<-�v>N�U����=�ө=z��= {�t|w=�==���<�qD�M�<��X��D�=m�%��r�zӴ���z=�c<�g����캣�=x��<(�J�q|j<\Dk����=nl������L�9G̽���=�J�=\X��*��t�z<�+�;�]q<���S��=���=Ŏ���m6<�����x��!cP�f���C��G�;?<X=����h<I_�<�lB�ȱQ=_�:ҽ]���<�����b1<�=T�r��&7�D���	�p=���4��=C�,����Qw��,g=�(=V�h=�J�<tR����=n*1������<2�=7�=x$#<�*�#^�=�N��<��۽�IQ�*��ڬ�6V�֣��2=���H4=��=�����2>�Ɂ�+���N!���(="쏼U��=�k�=�>>mL<�pB��:\�x��<͵��>g�=ܻ�=��w�	��=��
���E���?={��<��=4�<�N޽;�7�sA��F��"D��U�=ĉ=��8�+��=�ͽ����z�Ͻ"%>�[=.q�=7ղ=t��֛����<H��=���<T��vG�$c~�yc�<�	�(��t=� a<ab���ûdx�m��=9{�<,W��-V>$X���� �]>��½a��<ZS�T;>l�<2�Ƚ�����1�=Z�=&f�	i<4����= =:��8����=~�I��<�,8�R}=�#�=f~
>V��`�=e�=�[���=�EM=Ʀ�
����x��M�>ԭ�=�����=R�'�j��}��<;=��	=c �;a�<���Я'�?��XI�^~����μu&h��䰽@�7=��!>���<�t��^���Q�����>*�+<,X����>)W�9�>�M'�̝
�s*��fI�����=z�뽁�=9䍻b+�S޽���=+Ls=����`����C`>,�x��`�}��=�(�:�t��ך���s;��~�Yw!>�y!�ַ�4�<���=f3����<�μ����� �=_8��O-��)#>�W��n�=�2۽��;��#��e��$ؽ�y=�ԉ=�Di�$`���l���R��q'��&��*�[<���^O�<�����G�<E">] =�Z8=�g�=B~$=��r<�_�ս�������>�<i�<_�6>�C=cã����=�4����@m>��;�Z�x�ҽjC&�t��=�X��܇V� o�~���{��{==��j=��=��g<���~b{=�,�����r�=�=��<��ܼ�����`�J�xu�$^�efu=14=��=Y5��M;�<�K�<�u�3�c��/=
�:=m�<���r�=��`=e�F=)Nl=������6�<:<7� ��c�=ߪ=�5�hZ��eL�����h���0����"�g�)�.�ݽ�e�;#�߻4�C��6>��/�>"��N�=3.�=�A.�"C��c�=��h��μ��= ��=����G��"?O���v=:��;�9C=4���&�<����㙈<���=�\e��62=��ݽߚJ���<0��=qi̼;��:�=�a�=]�G��q >x��:`l�<�#�=�oƼ�M=��?��e����<߰�;�Q��A�=N����>�=Y6�=�:�V@"=����Yϛ��jۼN��={]����-> �$����=��3�4�=�:>~q�<�%���$�;5�W=]f<�{C=xs��r;�����ğ>�_��v�=��=H�>�f�=)����L\<�(>�>>���c���vs��(L==�	=v��rz���|��Y(�����<h�S<$Y�<�QȽb4W�[>-:�;����I*�<��>����5O>�;��=n9�=�#�ὔ\�<d�����=�z�T/%>�����A�Z)?��nڽ���< M*��˘�ᔯ9�H`���|�*���?$=�>=��R=-���G��żj4�<���3u>��<δ�:|�=s���^,%=oE�=&>�Y��<R����=o��=B��<�\�=[����������<��˽�����2�=��X=p��=��H�>�1���GV�TH�<�؉�MA=�T���H=�X"<���;�]����)��7�Z�̻6���W�]=~�h=j�3���x��=��n=�C>z���<��I�K��g�=��m��u=j�=�T�=��ܽ���<�g<ϼ+����2�Z[S��)=�� <�໼9"��6�w�=A3�<T��<Mh=e��=iB�<�r+�{�)�4��@5��b��tO��2"	�dԶ<V��=X� =(-/���c����հ�����<��;=�4�<6=�_~;�Yh=2Rx:�T<g�ȼ&Ve��;��l�W<R�"��4>����/e���ǵ=hI|=��>R����:���q߽��h=h�v=Zo�gO�=�����%���Y�=�ګ=D�<��ڽ�"=��a���W���:`�����p=��=P��=ü8�5��=t�>,��<'�����\Q=K9_���Y�I�<o����W=͂�<hdŽPA�<U);ϑ�t�!>�J4:�>+��=�N�<��=��=�7ݽ'����=*C7=�ϡ<(��=ԩ���=�7�n��MNF���=٪H;e_->6
>Pd�^�����L��j����o�-*=�;�¢��]�<�ۜ��H0>S����/��b#>����d��Ӌ�%͌;>'>�䇽 Z#�L'b��j�=����.��=ܣ���q��� =��׽0F	�/�<=_��;�1��K�=��>��<%��;#�>r�p=�.=6"T��-̺S��=N��=��e==xѻ�j=f;�e��k�Y�*�`�;�R���%=Ʌ0���E��� �T��=9=��;R�=��n�[E�=�>,�>J΢�0|	��>QN�,��=���m�"c�=%4�<r>=�*=��Ƽ���N)�o�<L\��}�=�܁�7'<m�M�D��d-V�@D	����G�;��=K�J���=-��5��=��*��tO�N�μ���<8B|<��H�(=���J;���L+<=��D=o�<�?�&����<� '��v�=r'&<Ҽ�=�=ۂ�<�=|�>�u<x�����ql�k�=�=>����r�=0b
<��=�¹=��=��=�=l�U�c����;-x�=,|r<#,��]�<3�Q=B�+>Kv<k7a��ND=b�=�Z<>` �+�>ͅ=<6=���<��t�;=�ν�O<:��=��=��Ľ��c=yfҽ�X�<*G
�����=%�X=�_Ƚ[=����:ý�>�Y�<s0�<��=]�A��F�=��=�z!�j�<�� <x==4J��K�Bj��ݹ�<	�#=��U"�=PN[>��x��}Ľ�eT9�>�5>a˽�0��5�m=.�=�xۼ�`�=����U�=��<Χ�<D�R�b<��<W1Ž �Q�0c߼��Y>RD�=�d�;q��=d��=��+>��!>���=&�׽���=�v,>K�.��%��\>�m�=���ʅt=p	�=>5a�	>2
%<F�=��车}T�Ѯ�;߂J��զ=�P<�㡽��	�^��f�=��0=*E0���=�}�7S���U��>����Ɇ3��_f<�����s|�� �=���#Ѽ%��=��N�D�`=�*�<���<�:~�<��hz=V> uļS]�=�^��¼�Ђ=�B�;u���u�XǢ��ʼsH�=0�6�������\�=��	=�=��>�&�����=L&{�1_�=?�>w�r;�<�׽�	�<`�<gŐ��>B<��~;T��=)��<��{=V�T>�=��>�m�B�,�-�<T�պ��;=Bw�<jU:=3����=�9�=A���U���u�,��h =HQ�=�|�0�<<�0�;}�=��+=e�5�B,'=yE�؝=N�۽�%R���<&,�^N>��u;i�4��J滾�����<�E
��[��41�<�N�=e��=�8���h<������1=�R�<K�5��϶=�$>>�0��]��{�;
�I��q����8��g=\�<o�6�C�e=+h���=��.<j��������A����\>���t�r�=US�=U�<\]���e�<��{��ۼ3�\>Y�Y�=_����`�=�Gǽk踽����G��{�x���=*��==�%<U(���+)<,ʏ��~1���;��=�ڽ��=�U$=6��Y�!>�a�U,��!����<D���=ွ�h��J�T�.�yF�<�U>X���#>���߰��U95=�'=�y��V�������p��wɽ�b0�=�H�����&@�<�<��K�f�Y���w=}�2=�M�;�]> ��N����邼��ǽ=(=`��=v戽�*���&�+��������������_س=��<_��=s��>�%<��;�ü�=7}>�W`�6=fն���=Ft�=�6��h>�C�=Bg�=���:h�<��=a�'��=��<)l�=�ͽT_��a`�<�w*��J���'���n��y޽�~�=`�=���3�<=�{ּHc<������ʻr��=�1�vu����������%>��p�
�$�Խ� �����P&��|?����'=��=;a�=.}7���J=��=���<�=#��?�8�;��>=��=9e��N�<o4���=%��>�=��+=��s���Y�^�/=��
=	m�=Q68��9��7��d�ѽE�*�5_A>j���N6>Ӷ]=��Q=Ҿ-�W�)�8L��Xz�=k��=7��=#���q���z��dx1=� ��Z)D<�p=��=����z�=))V���;��=W�>��=#J�+в=K�ٽ�&=T>������R>Kj��q�J��>�˅=�_�=|����=����MB]�r�D>g�@�tӽP@}=W�=4�s=��=���=�=H�F���8���f=D����(>%�i��4>�|c<��վG=�Ȗ=�Q?��).=�Tڽ�z.=�u�����=؁J��	�<��>ي�=��=�;G<�n>A<�e�;��� =��;�����=�:>����
�Q=B�����7���j�@����:�� ��E���L�o6����y���=b�ȼo�H<n4���񣽡ƺ<���dWB��ɚ:�7ĸ@��=�a6���?�V)�<��='�ּ򇼷Z�;&
�;T�-��Y��?L?=}��C>(x=9dE���y=Z�=��E=��=�[{=ij3�;zV�I �=h�0�'�Z�乛<��%��<�&�=�>7ɮ</?���I̘��'�=39�-�(>�N>�v=_�=��Q��n�<��=���"(�=җ�<m@�=YY�R�>l���1�4���(0;#=�м��K�6=�s�=	�3�*��<��6=#C��Ś�=P,
��Ơ��k�=�$o:��I=G��=�-=eQ=�U=���� Ѽ ��=_��F:@�=���@���/��oE==�6���	<���;�S]�1��=.��<Z���Й�=#y뼟q?�ݦY<o7�8�{��P��������N�f=N�=1Sʼ򖧽@{�< ��4c= 	�=��p�����/��=��u=�@��G<߃.�O��<�#ŻBP=y��=�D�͘�;����'�=�>��"O=���;��=�=c~o=2O�=+ߴ;$+{<Ia>"�%<M�=��=*W�s�;�i>�숼�Ѽ=���=_[��`�=ќ���5��
L�ri���L�_<»N2=~0�<��<�`�=e0�Sqн>{���ռӖZ<��.=,{=h=M/�<`wd�/+�_Z�3�_�s��=�s���Ƚ@q_=йƼ��$�>Zؠ��-�;a�>^�߽�z��*H<!�<م�����~D�=|j����>�w=c�=�����1����� l=�+�<��R� �ü��Dg�;��g�A=�ő��}�=�[��#S6�=�2�=�ݠ�%��=������n�9�����'��N=h�����;|�;P�;��S���<1����=���غ�/i�=�Π;=<�;Xi��jɽ���=+�ϻ�w����ν\�>����;�y��YV���\=uvi�� '�׆��	V�EP&��ٗ;�
�=uP��&*�w�ý��1���]�����/X��BĻ��A���=R�@���=�N�;��=>���I���@V�ь=��=�I�<���=#蹽#�<�f��SS=��=�[�=�&k<Z�>=D
=��5�=k� �Z��<����`�=�Xp=��;F�+��!�B�?=	�=�1"� ��<�M�=@�Ƚ�2D�*4�t0	��jV=&�=^zD��8A�t4y;	=S�=�r�=/]�;V2�=�I��H<�=�M����#<�)o�G�<���;�0����J�*:��<�TZ�B���7��8��ჽ���=u?ս���c~�=~x���=O!�<ys3=��}��(�=�_=��/=\aT=Ͻ.<ߕ��ɖ�_����>�HZ�k�<�H�� ��<.�q=��>X����@�=*��=ViS�i�->[`=yG�<\̼�6��8��<#?G�~~�;{��<���t� ��b=x�^=��-=��˽1�=��21���>===�/>��˽T�I=zyu<��|��F����Z�xJ=�=s�����=g���#� >B�<��S��<�6�����dzK�'�:������==?Ӽ��=Q���=��$>�� >� �<rdڻIJ1���ٻ9�,=pj�:E6��翽���<=�<�8��r<�m�<s��=��}���۽i�)<��=��=�D\�hNC=�e��LL�;�sI���:=��<�Q%����N<�J�=g<<�|@=*�ܽfjD>�����E��x=�Q�>#��<Qn�<��O��ca9����</=!�ݨ���>ɠ�=أ�(� ���Y>�ީ���V<ꩽ_�V�J�k�iی<��0��Q�=�eR��"���a�x�w�{a�=���W�Hy=t�"�=hԼ_�=l��p�=ϣ�=����G�����<onۻX�<��6=��w�c���M�=KjX:�!;>�e
>R=�o=q��5��i�=֌=�02�ó���Խ�=¾�=�A��d��:��8+X�m�����=ef���:)���P<ў����$�R�@�z?��ޣ��@Ľ��=0�>
�6�����Z��B����<��=�8ٻ>�P�H����<ǽ����<�f0=�/���C>$@�<�e`�}E>��	�0dK�b'*���Z;CAQ��|=9hy����a�b=y��(���'�< U�;�F��#/>�����;�W<�<����=��=ј4<"}���e �稅=(D��?�L�ս�p�=7쀼�i!>���[-��O�<{�
�~䖼����6���,�-=�����	V�<!���Z甽�ݜ<qv<U3��C��*O_=b��:8�"�����f��*�R>��߽�����=x����ا�<�?l��|u;�н
��i���׼�����%��Dkh=���=fϯ;Ő=��]�CZ�<Ա�� �;�N<O�=7={��	Խ��1>�q��T_�-٨=����P��g�=�"=��=;Pn��E�<���=�l}=>�c=P�=9.���̽R�=�)�_0>-�=�3���Z��mý���=�~��YL��w���K��m�84�9A/��<�f=����򔕼3o >����`�n}����<|½A}��!���>���<'��q����w=Z��=[�=@�=7x�=�$<�GA;��<	�D=b�ν�j���f���=k%����!�v��'
=+��<z�?��=�.�������9�O�Y��=�/�>�>���=z��#ɑ<yy=�>Ih9=H(�\F^�o,�=��w;�xƽ�=���dH��P2�=����`Խ캍=�q�=���=�f$��=�X�=�_ý��>�<"=9��=����F�ཚ�)>�Ɯ=��=Ś���.�FK.��W���=�B%=e�=Q����ɽld\��y��Ƚ��==�r��y>�� ������/�=J,U����<��>S�C�b%=�������=�5�<RPe�WB>��ؼč<�X5��F<����k����}���)"��E�<��b�X޽쒝=���=W�=���=��=\7�<Q3o=��M=4��z�3>S����;�$��y��Zd�=�/�����듽)	=Y�����e�$��<�/��i���g�=��R������a��=?<`�T�=KFt<�*���<����Х=�Hq=�+>j��=V�<���p�A<is�=R>}ǌ=�߽�����p���z`�B�c=p=>��y=1��=����(���ۼ|G�=Z"6>��=�=)=�:��<�os=D�N�fB=q��]�>��=�e�Q ��9����=���<��=�Q��yR)>�|�<�6���p�=��<�l�=cr�=�_�=��C=c�����~=[p>��J�ؚG<�s�;�.H��.�$D �.Tj���Ͻ�>�<*5�\S=��Ľ�%�<�DS<�U��8y�=쭽�~=���=/�>޺B�����R?<�8k<?">Ľ[<iA��[��`m��^�<�$�=����b�N�ҍ�L�輈_>_�=�M����=?����ɜ=�>�=�ߤ��>�=
I�;}��=�ǟ=����%�⼈����= ���<Q��T��UWP��ۊ<��]��u�������p9��7�=t�R���u;Ԡ��U%=s]�=�LL>������a�4�\��b5��H#<�h<�k=��>���!Ln<� �:�+:�'��M!<��G�V�U�me��`ſ�pZ�:����t>6iڼS�K>����W��M�i=>���(-��$Q�w���L�y� I�W㓼ݴϼ禵������'��Q�y��&�=$��2{=� ^����Dq�=-��V}���$�<�.���$=Kov=�v���U����>�4M��#��tl=g� �t=t@���v=Hhӽ�ԽЧ�=T�=;���E=p=�P���=���n<��ýb{�=q�=��ͽ8�]=D/=��=�P0�+U�ƚM�z]�����=�����=�/�<v���#�ٺ�=�<�� ��k,=r5�;$y(�➽���=3��=�9��{�Ͻp.s=��ɽ=ܯ�V��<�%;�v�����sy���>�q���&(���9=��	>�Ѻ�f�=:cٻ�:޽M�e:��=6�d�r��<5s1�MB�=��;=�4=��*������!{��ܷ�6��<s�:����3����<�+=# �<g�T��ȫ�W�i�e�X�Z���0y�!�=��:=�67=� <�b����H.<NV�=���7�";S:=���B���Y��*�<���x���:"�=R�P=�n>�)�<�!>������쐪�VTE=:�=ƍ=w硽fZ�<��=�$=�7>2!	�_)�;O>[=�Ƃ<�,�<��<=_J������(�=�4R:�S�=�c���O�;o��=��X�Q|/>��=�S��+�=e2�=yg=[�����=�� �] p<מ==�=�o�� $�U�=�[J=��
��e���=��s��G��l�<�OԼCy=��=K�i<?2A=i�Ľ*j=.nE=햤;��<�@��h�-T�� �����;L�=���<�hӽ�6̽*	�=3> =�/*��+>5_�ᔉ=G�3��
W;v�����=��=����ND�<�->�
=�r�<���=l)�=�g�<S�X>
>�=�9�7�>K�=
�a��i>��]�U-���)�=�����M�=�H[�6C�<�T=V�<��8��P����=*`�a��K=<�ɼ�׽���=D"G��ӼO2�=WN�=���;��=�'�>����=(�#��h7<���=�AR��ҽ�h�����Z�<S��=���a�=�G���,>��=�t>�
=��}\<
�=>�N�<���n�=F��<>Q�=ʰ�;{�[�%4>�ý�VǼ��O���R���ӻ1���>4�<�u�=p����ȷ::H����=��h�=�0�<,k�;��;1$o�}�=;���0=��1=Y�<R�(�q��=!�$�OB���U��70��H >��V;!h�=�m�=�.=n�e�Ƹ=���?���?�^��;�;�=?�=c��=:��<�G�lD�=�v�:H_ǽ�%<��?=���=�L�=X��8�==G�>�[=y����߽(I�=���d���=�_�=���<tSA�f��L	=��<_��k����'�<#NI<I�<�`�����=Z���'�K=��Ž�|���c�=D�>؋��ͅ�</�l�t�/�2��=��=��G�ۂ����=S�`=�����2�+�T<�(k=y75:c`�=�l���V��	UٽsGr=�>L(�����c�=��<������;ji�:r�qN<��ռś�;|1�<�����jb=`��=�Z>�Yջ�rf����=3?'�_L=?�v=�v���ł=�� >%���P����*��tF=ؚ�<�_���"�="ᎽS������&�ǽ^���&j���`�=�i=4��;p�ͼ�S��lK�g�==t=�<�����q����=�	=X�A�Tm
�:�g�<`鼿J��j�<&D�:��<5f�=��I�O1��+N6=Xi�^3�=������=�2�<wuy�lK<�e��`C����YQ?��&�<�3�=�Ъ<��<~�i���%>�F׼��޽���j�<��<N�=K�=�T=����G�݂1�K����2�;qC�����=��<��}=�s����=.�����K=`.Ľ����=T.>Y�>�S={��:�<�w� <�Ԏ������8>`%=�|�I�����<\l�=�I����g$�=��U<(��g���,7��?�ǈ�=Ԁ<s����>0�&�^��=�cC=��b���
>��F�4�=H~������p��=�WA�@��AG"���ż�=}���D��K��=�>��;ݫ��-��=q�N₼���$�;��<�vc����<8�9=+��������f��{Z���o>|LD����P����Č���8�?A�<*�=;k�=q�<�Hp<Z�v��GŽG	�L=+�G��>Us�=�3��N�<vm	����b��<:�w�4�O=�$�<L�����=��^=�*�=�Oʼ,>�=/KA>kGM�l�� l�=�b6���m<Y��=�&�=j����*>X��=r>3%h���F>i�ӽ<��������=
U<�Z��J�e(F<�;��9�=f�E�K�������Z��;�d =�_��9�� m|;M\�;� ��fű=��:1�>~�Ƚ�c�<�r>�mC�La6=S�=�e=���Ț?=ĐĽ{��=*�
>)ɢ<UȮ�_��ż����<1Ο<XI�=+a��w��x�=���<h��=(U[��ؓ=��˽)�B�����<!i<�F<���q�=1�%��;*0?>��<��e�d����=��=�����(=��+�G*	��#=<��Z��#�D��=� >M���̰=�P=���=,}�<3��=1=���<$��L�3=#z�<�1>�o�=�HؼϬ�<����n^5>�H¼I�%�z̪���>�Q?�ƅ��>~�>F�q=#6=��C7]=*�b>��`=  m=-�1�H�=*k�<�_��7�=�����ͼ"A�<Z.�=@�Ƚ�	7>��?=J'O;&�\��l������^m�<:6>k7��ݨZ=Q���}�v>��4<K|�=�|�:����F�A�]���̽rֽ��g=}�ּXg���M���c>����α��,#:��0>PC�=��Q<����ig;� >{(>5���m�.����=�'�<P^x�揺=fۊ>��=���<���8�� ��)&��[�:���=��7�._�Y���v��:ͽL�#��d���d<Hޞ���2=�J����<0�۽��;{։<p����q4>(�*=�*�=c�	=�F�&>*�T�>�v�=�>]A=�f>3==*�ǻ������q�>�h=��@���:��8���f��<� =�Cͽ��J=��t����;�I���l!=�Si=yj�=�U =�.�^����[>RK�=?Ȧ�uά=&ـ= s\�<8�=��]��NW���L=��P=��>����;�y��Ѷ�<�Z��sM��}�!;N����<�*�;�p�֖>���<֬=���=\/h;�C`<�5>/]�:�!�	=�߽<߽t��@>!o�=�=�|�=e�B�7i6���#�l��=�������[��)[>��(н�9J=�p�;
t=  m=R+=�Sv�ގt���=�E�;Qj�=��!��lR< ��
��_@~<�C-=t�>���=K�3�mWҽui;�X�Yp��n�=��=A<����{��b��q=��ٽ���=[�>���= ��<����<��ǮI�zn=k��=<l�I+���=_�Ľ��Uk�=���Bz>�G�=�^���׻=H¾��Q=e?����=.9��7��L=-�>"��=~���9���co<E�S��/>�;(=�W`=?��=1������2�=F�?>��K=�">D��*<��=5p�Ӝ��z�T�S����L�]Ꮍ
�>0�?����=��½��=�]�=˵U�FO�����I��o;h��<Rk�<R�4~�:�v'��L=����������2=޽OѾ����=�ѱ=K֪���Q=}�W>6�=D�W<���Z;m=�b<���=�����>�lo=��J=�I �Bͽ,�ɽt䢽��=$j��|o�����P��1>��ѽ�<�g >�(��`��AO>]>'	=��r��n=�"h>)�2���;�i�=Ʒ�=,"d�3E=錧<���=���:�e�H�;a��
��<.�����K=�Ҫ���)>S����м7]��jb�=�_�>ŗ�<�|=n�`=8����ޒ=j�T��"��M,��%�=b���������<�JS=a�	>�uz>8R��Zu>�X=��m�<�8L<�k�<�p.>�F�<|h��<8=�7�=7	��i�(�ZN�h��|�<z#=���V���$=!>t;i���#=��*�����E齈:��z��4mo��=�<�F+��p=�v� b��:�=��޽�(�=�j�=!y=-4ܽ���<r�h >��)�Of*>����<�:b>���	�J=�IE��(�;(�l����=u���[�=��c=�l8�K>޼"�W=�=͟��������KV�<͞I�ro|=�f�=��>�7=��,�}5b�Qa����=Lo=?~=��|=�)f=1O&9Oe�=��=�䮽�� >�㽊"p=/M�=����&�=�z�<�go����=b�=
<$�'Z�;g�һ{^D:�k�;� /=8����N�?P4=O�C=*����=ş�;�ռ���u(�<������=>u�<nT1����7��>p{y�f�f=t�Z���,=c�B�,Q�=��:�),�����i1����=Nf��=}v�����=���=v�k��Z׼���]�=ڦ1�O�8�-à��y<��C=�5>�f�=B�<�8x=y�f���<Ė�ۡ�=q&� ')���0=��j�S��=�k�=T��<�Ϛ=�H�<��`=���=縼]��~v�Kou=��;��F=�ګ<`�;�!x�5x<ț޽�'=,��<챫=j��`�9�iI�;*G��~u%>9��<���<Z��jY}�~��=z�:<Bӛ=M�=7A#<�� >��&�Xs*=��J&5=�f=��}>_=��(����Yۈ=��,:��{���<l��h0B=>�L=w`_=��b�X��=���.�c���0�6
�=5�;�✽.�h�H�ƽ����{���%6�<�a =�����`=<ٺ=����i(=��<f�=Մ�=a��=��v=Jl���?=�P��ܡ=K�<=����+���l������;4`<���<��D����H
= ={�d����%����?���ƽc�'���"=�; �h�;���Q;�d=Ns��V3W��Sp=q ��R{>� ���Y<��&>��{��G=}�K=�>M<�i<3:�<�M���A��Ϡ�'<�ػ=���������k��Sa�R��
8{��+v�����>є�=i]��XQ�����Q�=<�=lC�<�T!���L>�M�=��/=��OٽE��<�֮=�E�<�7�=���=�T=
��:��l��=�CA��mѼ����=O=�u5=,s⼗
���~�=�ϊ=�"U��K�q�P>?���=)�ў0�@)����j�Y f���ؼq��=m�}�Dt�=��d�=i�a=��'-��-���6U�<������%���
>W��������,m<Ӻ�=$�2�5��du꽫��=L�>� �z/���e�����0�:L��]�'�/Qe�Z�=މ�=��|=k��<���=Eh�<*|�=�ۍ=�<Y�ؽxD����<������T>R�<��#���V<�t�����/��)Yۻ��|SH���O��(-��F�=�D=�o$�g�:w�v<+=;=�jɽ�(���A=���=C�=ʶ2��慻��p��);�a�=W�=[b����1�?��=�ጼ)9�7
����h=&�F�<	'��R<��=N>��r��X<B1t=���=T`=A�2��ν�H���8�=v!Լ�1=q.<z�ݼ�{=�;�$Dt��c���+��n.�u�=�:�i�w=��;M���9����=@j=�E�<���:3?�<�'1�r�B=:�>;��Gj`=�7�B����I�U��k����=�����U<p��H�Ľ���	�ؽ �f=*�̽q�<�ƽ�J:	�%yl<5�">C{u�7j��	�"�cS�=Tg���=>2�/�
�9��_>5[�=o8�=GT?�R	i��J�=i�@��D�=�C.����<�����-�;�9��><@ͻ���`��=(J�<%�)>���#��=;rs�K�H��`�<������<��м\�Y=��<�-��<>G�J=,m�|2b�n)> �=�c=��:<�Q=�;�<r�(��<���=�7���[����=�b==�O˽����
ʞ=�=*�w=&*�=;��=���7���轠��S�Mܽ�t/�㉄��/�=���=r������;�4=��̽�6U�I1ĽAO�� j���=�`�=۶A������=~�=SK�E��=���Kt�6�=�=�,�n5�4\M��W=�v-��U���R���)����/��
�=��	�Cf�<�L�=�+�]r�=��3>,= HH=O���}�;���s�C^<�l �
ݓ�Z`n;�ҽ���Y��;7e=lD=nE��N>?V�񔄽lF�T��@�Q>B2��S5�<s��=��\���>Э�.��<Y������5 d<����u�#��<s��9��<�Nf=�K	�H�=$��=W��%�=j� ;�o����^=	N�=8&��$�����;�Xt���W=��P=���=���<��ؽ���=�E�=��|��?���xk=cx�<a�=��c=�Q=��<�.�=�h�.k=�j<�=�=	�<H�>)
�=Y��<V�=��=Z|7�g�:$�	=�i�=�b9>d-�=)���=>G�»DW>�ƽ��'=�D�������<>j����=G��Nf�)O�t=�:�=B�=��������?�'�V�u��=w��=�ӻ=�i���#�X@=�+н���<9$�= gV��]߼��н�0��=|�[�F�	I�<	���%��ЁU������ >fr�Q��=&T�=�&>w�4=��:��>>\�H<7�=���=і���=;��>�>�4l;R�����<��<@�<��=�|+���>�̚�yY$>3`Ľ,���v>_0y<C�i�,���&[��ZP�4�q������oM�5��=�'=�Q=M<�����O'��=��<*�=�ڙ�����AK�Ł=g�<��	�rm=��<���=�}p=�d	�J^;��2�<�#l��}��x��;�=���=��d="`V�H�J>�E1<��Y=�z�=���S
�=I>���=_茽V��>Sr����R={��=���=�#`���">Dz<��S��ش���>�Z�dl�=�co����=j�=�4=��<��=bx�=h��=��)>*�=Wa�[���=*�;΢o�jc<�{n�Ԋ&>8Nϻw��=�+�=�G��BrU���=;��<�=1���}w=�u?=���=��мx�:�<����H��B��ż	�>�켕�>=��R=l�����=9l<��=?�=	�(�'G)��θ=�곽}�K�	n����=�e�=2D�=}�=��3=���e�D�.��=���=V=�� =����%�=�w�<u�$>���<��=7�a��=��=��A%�< C=���<F�>�e��i��kV<��"����;Al�a��uQ=��������n�������<�(���s=R�=�5�=?���(Թ<��=zD��[G��&;3�� >��_��.ӽ���=r�x�E=�Z��j����z=G]<���J=��<'m����Ѽ'�,��%Ҽ�s�<~^�<M�<��O=]:<5����Ԉ��H=�O�x~�<�3	=x��^>�=N;��J/�<q�<���<�/�=�ID�R~ս�麼08�s�=�
>��"�������=L�m<&�%����X[=�;�<L���ܓ;(0�=���=���<J�==�X=AO�<₽��껑��<���<�ɽ�ݾ���8T�I==if�=2v�=:$$���&���߽�=�r6)���1�Q^p�<���/E=�a<��*>=�h�L��G"d;��=qw}�.O����3Mɽ�=�;�MٽW����E>�s�J�:���=�#�c�׽��'�x�h=/�=4wY=<L���
>3%�:�ν��b=��8�L@���8�=�s˽��_�G�������<ϥ���*��<(n���bV>d��<4#�<���8�2��=��;�B�~��=�vw=��Q=��G<�`�<���=#����2��`��Ўc=��~=U�:�P<���=�^=��Ƽ�y���=�A�=��;��];[�>���=z'=��-=�b<=�e���%Q<0���a$j��}ϼē1=�����=�#>Tn>��x�:5^�=�0�:ូ	�>W�]=�ܽ?�Q�����=�"=��;gD��T����i�n֡�nw_=����E��qOY=߰���_�<����Ë;���=g��<�g��IM�F���>��27�=�M�ʷ=+ 
>v�����swý.�b���!��:�=����eΎ�B���9���>=H�Ap1>��Z�y�E�Q�O=�D(�'��<������R<��=�?��u����z콘�v>(�����F���;CK�=X:=޲ݽP�:����h���+>�=�O���R��ꊼ,=Ny����_�fH<�0���J�=V(��<ݽ#N�<�=��Y=v�='�>M�0=��j={��3>�������̽ɍ�=�*g<og��Kv^=��8=
�R<6��: <,�=w�=d�=G�=�����v��V*<�d<𼰑-=�h*�H�Y��Y����<L�����?��♽1k<��E<1I�W#�=����:��W�(�=ȓ�<S��{�<�P<�nɻ泧<�cc�<�=J�L���!=��!�7�	=`�=�'N���˽��뽈���t��屯=3��=W{*>L;�=T��=�쐽A�ս�S�=`�=ܲ/����<��k>ʴ�=V*-=���=�۝=P�Q��=�����e�=QoL��g= oR�C�
="!�=1<>��T�;�D(=���=���=�j%�j>>��=\lм�g�=�<Jۼ#2ѽ\qg>���F>+k�;�K9��ij=��\���$�h��;�����=�?�`%�ە-�#F>1���~#<?J�»�� �=�2�<w+��̶=������=�>߼���=iP�=�J^=��������>(���x=�<!�|=��:B+�<m�x���!�1��=A=��Y=EL�j��6ģ����j<�=��<�j���R	=Bݥ=�P��m��.�5Wӽev>%$��t�=}��-\<9*�<�e=�J==�#�=̍=y�>N�b=�˽6�?��l#=�ϴ<�==�@{;t�&�v����S�~��<&<ڽ3��:����P�<1�I=Y�Q�>��Z������j�<c����?�=�
��˽<%sԽQ�3��㷽2�޼���+�d=#�ʅ1=Y:Ľi�2>Jc���<�/v=B��=�DB�$Q���<��{<�h���R�=4��=��3��x�;��<�pG=1�=tǭ=bQ��45��c�������%\�=z���k�<�H��$��<�}ͽ0�����X=:0ֽz�
>�O�����2�[��F������u	�<�_>��1;=&�d��9�=�eb��]{��z>>���%���n=���<�<�Y=1�1<ϐ�=�i=��v�=+�)�s���ݞ=��p�����B6�#��=���=�'$�X	�<��=r�սM�ǻ�L6=�a�s$���n=&>��RC�=j��'�<9׋�@=S���]6�p����F�=FG���q�ք�=OB>[fh���<�P���<���<m¼8��=��+=侑�:�>����dB)=���=�M�=���[ݽo�=�� =<o��?ڽ����O,V�q�A����M�=�!ݽ?�s<��>N�=���6�p�<L�v�%>80
��~�=ҕ���=4_���\���;,���U;-���]wN���=��G<b�ýcXG�Ak=��=m`5�|m!�w̞�{v�<�
"�����jw�/��=�t�=�,v���ǼX�J�<�X�;m"����=T��==�8�(�=���R��=Q[��ӱ�rh����=S�½�z�<�Q0>�����<�_�<9�h>��[>v52��=W\F<Բ=�B>01>��<7�1=i'���V��s
=1��<��=���=T���bG=��7=a
X<�V�=,�%����=fU�
 =��4�'f����=�&�=p9���q`=��-��E>�"żqp=|�R<a+Q�Gڶ�ކ�<6�(��L�������=>.�<�EY<�hK=e%=�{e<�����Uy�if=,�p��4;�S=:�s�_f��<���W`Z���C���4< z>IR�:��<.K�<�͒=�?=@s:�Į<Y���H�=}�������9	��vI���
<�߫�=�-�;��=^��=Ѵ�=	P?��Y =��p����l�;>��ͼ�.��q�����M�a=��=���<�����W=�<��%E����=9��Wp�=�EＦ�����*�(ʽ��<.(B��½A���c������I<�����=��)\ ����<���l�=PG���Ӛ��ǵ�6b�<#s�����޽ٵ�=�%���<BA����>>�ȑ�*S<�=�<���$;��!=�C=<�0=�B�=�s�=�|��y�=��<Ox��E�D=&���A�O�����$n�;4�
=!��☽�@��G��=0�}=q>���j&<����=�x�<o=��w=!">Է�y{�5掼�Y%���=���<'�U=.֖=O�g>�
���!��,��X:�=��>RZ�O�=�G�K/��ϽQb�=�4;>a�>��Ľ�q7�*>�=0�`�|�o����=げ=�\��������=�ګ��_轑��<%BH�u9ý4=>��=w��T�2=�,�=YÅ�苏������N�çֻആ���.��+��A>��G=�5I>2<ʻ�u2>sL�=�~����m=�ā<�zK=�r�;���A��=f\�=F������;2Y	=�=����Q=��ڼ�>ټP���>�0����=��P=�I�=���:>�����y9v̓���N��ýx4�= ϰ;(�%��3�=nK��s_<h'�� @-��S.<�?$��==H_d=��ݽB㍽>�����m<���G>R;�=�9�8�g=�� �e3�=T����$=`��V�=���e�޽�/i��tݻ�K�<s��v�P�(���o��z���ż'˽I�U4=@�&����Y��=޷轷��=-��0"ֽ�Y�=�p��<N �<����N�M=&?��&X=A�ԽV�����O�_��=A�������N�w#V<����GJ�� ���*�Y�ӽ�%(���<���T�>t�=�'�c3�d�<Ir<$h�F])>Y��U�n�b\���v�l�Aֽ�Z�:��<�U�=/@�<X�;��b������;i���K=�7)>�x�=�@z=��=7���l4-��=�4�=�[��,V���0>�]��&��\L �t:�=�=�Z������$�=��=�H�="��9���=�������><�����i{���;�] ���<s����&���=l�H<�]%��W���8=�l�="|{<F�� �=m�'<��ǘ�=�<=��=�\ݽ���=O���gf=����`�=����轂{=�<�	b�$c%>t숽B˿=-L:���"�!>�G�=����=
[�=pI��g���%�)�v@�=.1����j��.:��
�<�@��宽�W=�������V�;�_���ν�i�=�]սq����>� �ʎ�=�iu=ذ~���T�⹼��@�����=,>]O�����<�\C���Z=�U9��Y��)U�=�������_�={/��#��R�ý׻��U�ƼG�<k���SV|�vI��R�� �k96��z���>"?��h[N=��:>��=�=��=�ϼ��=e���z7�1��=�=�3 ��1=4x�=��=�w`=M�O<,��<�e�=�핽pg��=������ٽ ��;�P�M���� ;<��U==���̃=�ӄ=�p�<���<ju��,[�=k+�<�<f��<3>7=���=��I��9.��=K^Y=����\�<�?�|��=�q<�Z�<@-=�dv�~|
>M=�<�B=8�^>�/�<c�
�چ9�;��1n�=1��=��<��(�e,>��_;���Wm=25�?"��/�=��=hWJ>������@</�=f�3��V��F��:���<!�-= �N��ƍ=�E=7i�=��;"����Ͻ��F��=�}�=H����L�<�Z�콇�a�=n����<N�S=<ㅻѱ���2����X�<�r=7�R<�V�<ͽ��b=��K�v4��R��"���o���f<�� �����m2=I��<��=f�<�`�=�=t�׽s�=���=�|>�F=
���4�K���9�0��z����E�j���=ޖ�uK!=ȗ�=4:�v��<�!��\�:�j0�w�l�G�+;���=��s=��-��31������<�<����=���"v�<��<���<=�?�Oq=ʯ�=ʧy=(�Խ��}���;�l�=dY��b���#�����˔=�$��{�k����@=<����r�=�Ȩ�Hx$>@�'��)%=bh�����=�t��:4�o�2>�(�"�	>ĥ���Ƽf=�!>�hh=쌉�$t�;+�=�$=c�6��ؽ�!���Z]��?�<�*����x���K��Z=l�ҽq�K���<�m�{p���5�2�o=��=f�V�%�=���t  �\��=�߼�A>,�����{H�5��=��>�H�df��p�޼���/�Q>䳠�v�b�P@�W/�= 8�;Mⶽ�@.;\�="�� >�=ď4�v2ԼN,=�lx<��<�%>S�#�jdG=~;z=���;���z+�<�|��VP�����8�D=��½��q��<"�=b�P>��鼄�=2��[���U�>>�"�=~�=y��;�*����1��3��g��=�����<#�=�F<��=<0_����<_*<~=�=�� <8>���<�*�"M=��3�5�]=+�%�X����y>�n��<r�<�A=��g�ǽ�4�<��+=�J��~ɽjJ��O�:=gQ�=A�@<����SS=��4>�=%N���]~>2�c?�+����J=��<�C��<�R�����C4��8�=�Ѽw%=;��<r����kQ=qQ}�W��9����G�)��P�9E�=����I]I�f�&�Xފ�f�\=F������=yڼ��
��f����=����lE%>��C����<=�<�{�<D����Q�*ꇽ���u��<W��K�=�(��"9=�!>��?��-	=�%�fA<�=�;�#e�4Ӧ�S�>\9���̊=�<�0���(�<X(껆��=6��=̩G=����"g<��=��p!=���<�8�=Ӥ?�T��=�Y@��J�<�"�a�>�]������~<ju��(]>�'�=�$�<��-��Cϼz���h�<��a<�j���<"��='�n;,}�4�i=µ�=)[��ɽ��'��������E�=-�_>��;�<;�.ɼ�L1>k�M��5����B=5w�D�=�r�2˼���>'������T������o�/�'V�;a����F_=�G�<4�ǽ�G��9.�=�:~�<����,P=0�"�lm�=t���:W�;��=�������=�U��ˊ�YR�d��o�˽��d,s=��=��d��t=�vX��oC�f�	=&���z=�:#��f����=��<�>`O*���S=m�.=��*=�!��={<s)>�Ry=V� ��<[�P;��!��M�����B:>�T>w���6��l:�:J��Dٺ�Q�/=�l`��0�=��=�e,=�ٗ��V=qM���Z=;C�=Q:>d^=����@�=��=������<��9�(:"��=�.���8<��]�����I�c��땼�~�V,_=�㚽~�>f�q��	�Ɲ���WP���Y=:=n=P��e�=�(�<�K�����<(]�<����(<J��9�l=�Y�=]�C���=뻝=��<�.�����5���|^���Ľ����W�<L��=l�?� ��=̾=��/�=���y�<pټ�K �W���48�|,Žj�e>�_1=���_�=���=S�=�T��K�����
��%oT�*Pڼ��0<�x����<�ط�Hs�=�Z����A�jꇽP�Ѳ=�>��	<x�~>�~��F��=\�����B�e2���¼�ǽ3XN�{ړ�c�d��6��O�����=��[�6ס�;+>=�սA��=��='��k�4���{=�	���:�8=�:�塇�{�̼�����a���\P=F��=�e�=�p�{(>��=;c�=���#�<~4.=��$� �>��Ӽdֽ��#=:�=�����9�a-=�Jz;'����R���WH�����0�</�=�"%<$��=g2����>�T�=zX/�vK�<��<��<ۆL=%�'�,�'XG��ۼ�9���~�"ͼ��=S��<�!��EE�<��8��:ذ��=�	=�S�	�n>�J8=�ʰ�tҍ= ��0ea�2��=�d����P=��=]��=�B��N�4=kn=y虽��=��6������#���p�'> ^�H���`U=� s���M�<k�=�'M=�1$>/�i=��>	ٞ=��,�����=�=2Rj=2��=�*<ԉ=o&�=wA��g(�;o�=�N���=?4��� ���4�}b�=�ᙼa���AP�=5�f�Wܽ������=����(�;��O����_�	�[�>��#=�V&>_<���=q��<<�5��>�̂=�4���=�;#j�=��Ҽ��3>���_��<؝R���=��㌗=j�P=��������J��mN�݂��>���I6����%=И4����=U�->���=��<�����<ۥ,���)=��7��_�:�[>�(0=/c0=J��=Ղ4��-Y��=;g5�	M���u8�Q�E=Atp=֘=;�=2Y`=���=�[�<��e�co<v�=�t��)�=�9��|撼�q�<�^h<O\=�,�,��B_l��2����=:���V>�h�<j�Ǽ�<>��i>���=մ�:t���,�=ˋ*=���;�T�=�YҺ;�k�&F��)>�=#�]Ľ���= �;k8��#����e_ɼ�=�=y���Ǯ���=^�N=�ڑ=;ż; �=���=�<���=1G���B��ڗ����Nѽz��=�=(��=Nu�<�%����=���=��<�:0=�꥽2A�����=�����=��N=j�*<
~<�B�<q
s=�2��D��;����
>K^-�T�@;C�=��!>/`0��<aa�<�P*>�t��y��4�s�w�����S���Vm�f�l<�@��i��=�c��$i�;��<
#ü0v=����"�B�ý��8<��=�ez�>�[���<1	�=���=酱�Ñ���H�JQ�;Ql�v]�<9�(��I>��=��/���m�:��<��:���n�FN��'3
<�J�Sq�C=�S��d��=���<�N��Tv�vK�@�C���T= �m<�e��I���@>�k�=_�ż���<$���ꊍ=-��=ͤ
=,�*=�9 ��=e17��ɧ�����=�={�k=('ϼ��u=�t��f>�����5�~�
�>D��=�l
��y���~f=)8p��c�=Fu�<��#>,��= /��,��P��;��=74�<4�>l�p=Џw��M�=���=ˋ�=�=5�=�0=<��<��!=6I��Z��@��<�Em=�ȩ<S���î�����<W��=��>���=!F-�h�=}H<�-��mA�����=��s=Ɇe��N�=�#>~���&b7�z>�M%>�؜�?"��$ì�~E=Yag=�i�Y:5�=��`��<u�z=S�=<H��<-��=ttp=�ׁ=;�8<D�M�4�b�=���=�=���1�{#'=֭��N�=r����=�F�=��<�
��-�D<6',����<,*�=�| >n�BW�=�Qڽ��G�	�Ǽ�U>{n[<��r��Q,�zJ8����� >�,K��2��0_�>��=�pJ�ced����=6b^�����8�>C�<�G�J�T㯼�l�=�}<��;��֘
��
����=���<-�$=�p��H�����;:wn�c`��Z��=�F�=Kˆ=���=��Y��EW�=$D>dw�=����8�D7�P�˽�p�=ӫ����9;��缔ch����<�Q<�<���"��z��Wx����g���=���t?<�
>=���=�ѽ��=sH�<Y<P��=���+=�����=�Vr=LZ=�"�h���k����=�Q�<��ݽ�SĽ��=`Y��K=$Vмa)>�#�&�)Ⓗ���<�A=��|�*���@�=D߳�4�޼�!��}��rh�<�%�=x����)�-�/�����~��=re�<�=�:>(������<�d��Ug)=Z���g~�=ރ�=Ϥ���S;����Z'�����<4�=�t�<����.�=�7=ZA	=y�g=�o�;ບI�=������<1��#g��(zU���S�����D!���q�=N8��약�?K=��=~��=]�=(�{�\�,=��l�v���g���tW�!7"��𣽡%���=I�g��������Ѷ;��i��vD��:>I�����=a��==��NcP�8&�=鴝<(�=z��=��ڽ3�M�3m<qX	>�*#=P��=�7��f�ϼ#L+>�� �+�ͻ�O*>��=�$6=��x���=�F=!��=�)��򰮽��~��R
>�l�<��1��x�=Wk$>�����=�s=FΗ�R�	��ɖ��>_�>E��=�}<�9=�o=�V=�1>*�
�e=��|<�d��N�<�u<��9�=�/�����Ĩf�_���:tp!�L~����M�;3>)��ȩ����hd=">���<�"=#DX��4>qV�=�4=;����?�~H���׽�:���7��~*��Q�a��8�=`����4;���=L�=V!���ˁ�!�Y�ieK��xܽw5�=Āp��<�ߊ�>�5<���</)�=ܻ��@��=_��<�>�	�<��T=^݂=K)��?��=�'��7ۻ^<=�,b��t�k�<j�S>�ȽA��:_>[�?<VW��a�=�<�S���e0=z--�b/�!����۽�.���c=-�>�P�=Ej=�ݟ=��=Pj=�=���o�<��K=�*��L�=*�
��=��<��7���,�񺂽���=S�p�/�r=8���O>�G׽���9�=���ƭ��\��=y|Ǽ?E7�)J=�4���ϰ=`0>9�=�Ky<��G��.���^0=mp%;Ŗ�3�>L�=���MR�<zG����<���=�����Z/�N�<|�=�j�i׻=�ỌY�=u#���{>�=sh!��䄽�����;|��<c��=��
�ȼ\�<��;.j�=/|�=��ֽ�;�=�Ws=G��=ǧ���37=�B	���Z�M(�=�=Y�S�K<6���\�M�=�윺ե��պ��ZM>�˺�F��<���=��%��j�����:K�=�v����=��{�+�;9
�=�[��="j��
�j�\�Q��.<�̧=���mIF=w'�=l�
���>%�ڽ.���r �O�7=+S=��$=1�&=�eٽ�Յ���">�
>����>��H� y��I�.c�<�j8�� ���LI>�R>��4>7Q&<�Ԧ<_�=����l�=e&��W>�s���=�&�'�����=�.�~.�>C��������G�=�D�<��	=�a�=�=~����(��b=˙=f>���I=i�>Rh��%�<9����ϧ=F�J�p�=���;�vн]�R��'>������=1]�=�~�<ѡ4=�A��j���G=��3�H�?<�T>���=�v��Ӌ9=��<	`�Zn�=��;u2f�,4�;P\����3'���x�`�e=sp�==�Ʈ=.`f�"3=��Ľ ����=�qj=��@��n��WV=h�ེ��]��=R>B=6L���c=�����=v�t��p��xZ;�I<{V=��=H�\�z�=�q6=8� ��=���
OƽS���=94�<{���W���ͽ��ýॆ;�h.�6�=ѷl��1�=�vJ��vʼ< ��� <D"����FXw=0�2�D(O=P���don>(<����<O쩽)!�`3z��9˽F�;��<������=^�>�=�����~�f��=5Qʽ%����/,�����+���,�LJ�=d�=�*��˽	av=x�P<b���d�@=�N=���<�<<R���(L��g��=�g{�gf��- �<�#�=Y*��ȗ��D�⽮)���=�J����p��Ul��P�{���ȯ��������d��?:
=�U�'5����L<,�����E�� >�7�=g�&��<�/=1Ja���=@��="�>>���Oy��)������I�=�3$=��B=�Sb=��>��=Ķ���=�<n�����=]A���]�=.�=��=ZG��l�b�\��=-X�8,=��=r�׼kv<��k���̽=b��O��=4r�
;<�իR=����2�����u�����=LS<S"&��H>�r���[ȼY�Ľ��]=�2a�I��<��L>��a=���<}�X=�3�:���<�����>�6�v_=�̱�	��=܅�����=:��='E��oV�<��>$4J�>�k�/��a�=9v�K_G=s�}����D���Z������=��=��;�z<�펽z���=�D�h�=>�D�=�&;=h�f=Ѐҽ�0�=,�i���Y=�����Ƚ��t�P|�=���/����ͼVӵ=.Ϝ�(��l���s���4><'�������<2�@�0�v��:Z=�����	�����<v��<wl1�TZǼ��A<>؟��a>���E>Bw<IN�==��:)�=��'�����=�ɹ�Wv2�J�>IN��n!�{@���佼��=F��=�LT=�Ń����=�F�=��ν�ӽv����g�#�����½��v=ݮ4=�ƌ��2=T.���<�=>���ἤ=Q�H�zUϽ�֊�<>�HW<�B�<�"6�\D=�|���W=�+�|5�<�5�;�rҼUS�<�ƻ�׏=)ǥ=�5>�_c=�@��9#{���7�=+5�� �����=c�����<=*rؽ�Vi��D_:z���>2�c=G��'��9���V���=��Z<��G��J��큟�8d&�p	$=
׋��M�<m�0=�1w>a(�s��3�=%��:�[�=��&���p=�F�<C�N�c��=T&=�	�!�->��<��=_�>�����`=`7��I<:5�t@A=��)�xX�<�+��S�=���e=:L��˼�5�~<�qƽӁ>�����:�"�g#f��/��½ $ｼ�7>/'��K��=�`��{�H˻���=-�=�%������'��R�v=�$>�ԇ��]���k�<�Q�=4c==�
>�ʭ�.�];�ټ�0��=^�:�+n��s>��=pQ+�v2��P���Ӥ<�%A>��J��;'�p��<�����½�e�NZ>��>����Խ�h��n�=��_=��#>K��& �<�y��y����">��������񏻭�K=��=y�%>k�=U�V�BF�=�<p�AT�q6�=UT,�b��!~>�=�L�;��>����='�M>�.= �}=:�=~@Ӽ�=#dӽq�=�|�=I|��*�=ka0=ш�=ob�=w`�;&-�=�ˍ���ؽ�3�}���.�=�T=7��=UZ�<F¾����<�C%�C���\G�E��zՍ�i�z=f��=��k��3����?;󼋾켟�;]G�=C.�<��=��3>�;q��!�=O�<�&B<���<}�������Om<�+���w=��=�	l���묽�Iy=�Q>c0�/�i��w~��!s�%���<Ӵn�"r�����=�w�<˃=Od�
�ҽk�ؽ����z��=�>�<0���A�J<���ݐ�������="�+=7]~�����=�H�����:k�=w�f�	���<���<��a�2Տ�!ay< �纳�<�	8��h���<��=u\��N���&���������S�=��[=�{�9^�>�
���G�w8O<������.=���)�=a~½t =���=|��=���='D�;Y���D���ݿ�w����=, �����=|��������j� ��<{�'=��q�+�5���˽��g���=����a���[0>�D=�ͽ*�Ӽ��.��sҼ3φ=�`�=.��<���!J�?���I^�p <�Q�<Ə��� >�ӽ'����� �=#���O<�Q���<qз��%=�z1=x��*�;�s�%�/=%a�=P��'��=�	>�\,�*y=�t�����-T=��˽o/ɽ!��<ɝ�=1N�=�U?��~T��p�]p�<��=��żc��=#�-�}��=�<
��<�c@<N��<4ja=6�����<��,�~=�=��>���jo>�����6��d_>W��<P��=��=�T�=Μ=��=��L_�=7�뽏Ϥ���=7z�=~��=��-�z��=�&>�z�i?�,�z�t�ٽ�䲽w�=̾+=�&��%0>�w�7(�=���=��6��'��U�=�-A���˽ ��(Ҋ<2�Y=���=�#=���M�h=�,e=��Ӽc�=@�=�ř=B������L@����)�<ǡ�<��>��>F)ٽ@DT�����JMZ��,˽ކ=���q��V���,=(�ǽ�t��pѽ��wV�=3O���r����3�V�Z=��R�T>y���-���p���l�֦[=�9�<�=0=G�;>�������<g�\��5�=�vQ=GB��+��< ��=KK��H�ɽN�<�Sǻ��EԨ=�sĽGp2>����0^<[��Gy��+?����=�4��4=�,�4ʹ=Z|� Y޽
B>�Ii�*=?�O���*��˼R�ֽ/�8�s�=��T=Z�Ž�Bs=w<�Ʊ<=$	� \;�d�8Vu<g>I����:��M�F"��h���l�,��;�b�=g b<q��Z޶���=̺/=�==��<X��޼/����Ľ�OA=�4�=N�;���=.�>Z�$T�:�bֽt��;g=��G:,>%�=���=ȭ�<�/���H����<)�f=S�=�'7=r�����x=^���!��<.>ȦԽ_-��˽���Z�#�ǽ��=���xn=fA���@A�^=�=I�T=m�<{(�׉5����Vס�pq=b�k>�"���<@*?��#�;68�=m���1�},�=q��<�l'�k��=��f=��뽜�#=G,=/i���~�����=��=�
�=b�=r
���;�NA��	>%s�:>��<r��=~�;���񍉽���=�мo~�=� �=�-�=�	��<��->��<�����G�u��<U|�=���<Uٛ<܋#�=��=���=\���<?�G<
}�<��4��i	��{=���=8$�=q�R<�T=t"=�/	>6���'�;���胲<��ڻC�=���<],��+φ=:��olѽrՖ=HO]=^*�=_<��f��I�U�b�8>��n��!�<�w=4�=���=�ﻺ�$=���<wƄ��}<�2�r�=�;�,P<o�=a�	�-��=��B����� �=0Z�=K������xL��i�4>���=�勼����,:<����=�^X� t������(n���3=�7�=C�޽��q�+��<���<Kkh;L�X�15�=�����!�3},� ��">>H[�:D�>���k�=/�=��l�r����=9,�=�8꺆`��Z,��1~��H佒�=[���~�ح�=DZ��xS9��%=��=%bI=�а����;��<�O��D��=gI�<$����~�T�4=*��<�g<Te[=���=]5��mI>�3O=Y��=c�	���=W5���1�=�m���]��G�"<欽
bs<C3=��=ㅋ�G
��c4�y�=l�H;�����= u8=�>=�p=ɻ(��<*N,>�����[K��b�Q=]�M<ǣ۽��=_���8�5�fݒ�g47<'�3�����ʛ="�6�g���j�=N���=<=!��=���"H=_#�=+��<��= �[����ŏ<��<��	=��b���u"=p,]="�=�ض<�f��f>��<���=1�f����<�����D=A�����g�J�/N$�,M*>���2����+��G	��8佫-(�_.���Ƚ����!=X=c��e�<��ڼ�꘽v7���%��;�9^Z�<�J�=�߽
��<6���9H9<j�����=�d�=�����S��%����; ��\����=��G��8���Z��nm='o�\k�<#������L��<���:�s;#N�=�w_�Y��U��;��ý���=�V���W�=�w���='۽N��Ɖ=F��=����A�'=�r�Ɛ߼����"w�a���s7=mc����=��E>O>�'�=>�y�<H�>=�ɽ$%��z��1Sh=>��o�=���=�ӽ*��=��A�_=�o>h�����Ţ�=�2�=�����ȼ�=���p-�=h	 �c�=�T>
X>�D=`��=KP8>lՊ��A7=��=JR��|��[�=��S>�>O=� 8�^���~z>�:�+�ڼ9��<2��=NMP=TGa�P����;h����=�2~�� >��Z=��r=�?<�s"���=��K�=��L���)=�
���;�Z�fN��`�=E�=.������i�>���=�]�<� -�����[=(�`�#��<�U�����#>�n�=�b��3j��W<��=3�}�If�h���M�=�=���C���=*Ʒ�ۈ<́+<���==�!�=���=��=�v> ��=��=b^�;0��l[;-�/��#<�K�7�le�=�=�=�ɻ�N: ���=O:�=; ����;n������3P��]5��v�=��@��kC��Ia�٦��ݣ��{�	^Ż�a�|�b=ݼ��QB��t�=8�<=IJ0��!n<$/B=^�=�=��=���=ǧk=a�6�%�	;Qy��л�*�����ebJ����U>ٟ�~���������~��D��d�=]�;i��􇠼�� >R7;��<�',>�==��=�WA��K��T[�=�{n=a��=U�G�����ꎦ�w��̘<���;��</D�<(�E�N�p<� :"�ý��<=�b���<�=�����h��N�=�\�=�-=0n�=�>:j���@N�($=����l�p=ܼ�=�%�<�*�=mt�=�D?�)̀�J�)��I�<���X
^�6I�=+���.�<�{�:�=T{�2O���>�gǽX=�׬<<��=��Ž������"���==I��=:C���%>�N�}���۶����o>�)#=)뷼(zV�{��=�T=�䧽K�=C�*������M��}|�=�h������������=��:=-$��/>R��lC�3��=�ڽ����;<�ѝ;��������/��|�%ٻ����o�<��>�"����]k��k�R�Z��=�帽�������\#=�v���/�<�r<���ɧ��u�=�E�=�FU�+��=�\�r�<D���W�=�=�D >�l�=>8i�ƹ�=5�q;PKړ�� �  � PK                       checkpoint/data/39FB ZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�G5=�W>��=�~��j2L��o`<P��<d�f=Y|�:;�=��a��>��1<�L��=�sݽ��=5�4��IQ�+��Y;������s̽���=�	>��=���S�>��T=�)�<����,>����-��l�}�m)>��=g��=�ڊ�����M=��udm��q��ļֈi=eB5��Y>� ޽�5%=�<=�7���<JYz==��Kc4=�*�=��4�Q�޽�.��:�k����=�'�=��=�i<yl�1��7!<�������Y#�EY�<��>b,�=��=3OI<���< v�<��(�!�I>i��<6(h=���~A�Y��B�==��=䩞��/�<�=�r��9��=��g<��X=���#�_�����]��1�����a�5�귂=�!>K��=ȝۼ��S��]#=��~���ɽX�==+�<�"� b6�(�=4(�7���r�� 8��E=<7�=���;A���M>P��=��g=e6�:g�ƻ�Z��5����=��\�Am���ق�WW�=�g�^�	=��L=�V��=>��;uR/=s��C��:�Ž�I����^���+����=��~=q�/;^l�J=����-q;+�h�(� 7�<�Tͽ�T�=���<^]��D�=Ȧ�3Q8����-=i�>Մ��!ܬ��1>�_�M�=�ɖ��D>����Xv�=^�=�l��=�?5�Y��;���l�������(D�h�f��]a>2֠;��>l�B��6f��6�=-�>��>/�W�9Ƿ=��(�m� ��A���>�x��ݤ=�D=�����_�����=��g=}�=K��tA>i������<B���,�A=^<��7�d��̳=Go��Pa�=���;�����<�?����=k�=��=ˤW<Q��=c�ݽ�����ý�z�=_~9v����j=���\�_����=�xR�ή�������"=8��<C����P�������'��=^�<焻��*���n<>���=ǡ�=�M�=;
���=�����S�,�+=���cr���^޽������>r�½��׽�@޽������罯�J=*L(��<�=�rx=��=��m=	��=����WM>0 >rz>�д=��O��<��%>��t��Kp���R>{�����(ս3!:=���=d��Q�<%̃��O >߻w�g[���n=JQ��=��[=G����~�����=��=fj���gm=?~>=
o��>L^���^�=��=4i�=�yK=@��<��$�~����=����q;Z2>w�=��̽m�;��~5>ѓ�<�k��?	�0Պ���f>b��=��=���=�!�����:���<�x5>�����r2ǽ��=�Ժ��~
=Mnt=�q�<u�.=׮�A�z�Ȩ��c�:]�M=Lm>� �
%d=a��u"�9�"=;�o7 �2Ϲ�2���,���KZ=�>�ʽt@�<,͂�lH�=s�����2N)�1 >k�.>1��<qV=^:0����=����Yq>�"Q���=yж<w��;��ۼ`��=N�=e�&<��j=XJ)��a彅��;�?���+I����<輠����N
��a�=�Q��0��_CT���=+�b�I��R��<h���;%�JL>���=�c�x��<�y�0J��rn�� >BN��k>����c�=r�^����=��=^�s�l�<�60�/��=�`�	p>�B��H_'�и�xd�=�f=sM1>�5�<\�ݽh�<�o��_>��;�	|�=>ʽ��2�E��=��4��!x=#�>)w�=�J��^��>��{<:%&�/Q����+=�O�	�|�ܚ|�^#>.�ܽ?QýCrQ=�$���>�z���a>���®=�[�=c�3==�л ꬺ�������E�#=O ����<Z�=���=p���z�=�̕=�.`��C�<4�=2!���<��=���)<PK">�o�  �  PK                     1 checkpoint/data/4FB- ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��46g6H��5{NU6�е�v궚�\�'�5�,c�5���m���A���?�6���ت��%�}��_��x�����A�4' �
5��T"�5�tĶ��'��6��R5�6>y˶�='7�T���-��(L�k�6,[�ՂV6�#�v26*��`r�'<7��uS�"'7�P��𶚷p5�6m���öZb���6���uy���	�{6�[�6��z���D^���GH��z�'j.��87�yM��J"�6Bh��7P�m3ൃ4h��5]�6�Ǵ� Q�5h ڵL�=5�����5��25�x�6ز��3����u6\��5��6\�]�̨5PG��?p6L�6��46�!6��6���5���U!�6uG��X��D��6��ڳf5�A'��/h��5๋�"��	��PVж�<6���5��5\8�6�w��r�c�����$��	J��m�6�`w� ���m&�6�]��� ���6D�I��@���Y�6fG6���8-6�d�5I�B6����M6a�Ŷ�-�5���5�����SV�µ�Wߵ���p ��SV5v�Ѷ�˵��q�w����ĵ4狶)��d5�*��`εO�6�5����5��i��0�5��׵�#�L]��懭��.�5
�ص4{ ��J]�ÌO6�i����n�0673��kǶ �j�h�s��2A���z6����Y.7 ��2��5�g�6Ͻ���)7 "4/p���~5s޻6<��6 ���<k6�Y�6�Ū�ԮZ6�[�5�`	7L�,��h�6ք6�P7����T�,������w�5�?7X���3*���j�ݧ����������6%�n<N�r������ ;�4�b�յ?�a� �R��j�����e�?%W��A@�:��5^	�6�xǶ��d7j:�6���
W)7 ��:cP74�6Nȕ���m6�f�6ŏe6�sn6��M�XD�6�MZ��nl5Z��5�qk7��L6F�M7E��6^�D7�뵆b�������	6��7��[6N��5���6/��6��b4��5���6i}�6���4_6S�pqd7�^S6&�P6��7���D�`6�P5 St6l��5���.��~c36�j6"\���5�]D�t�6D������Ӷ�;7@
�@n����T(4�o��Qe������M5W+���oݶ"�׶��~6Z�6䱵h��6,������Z���"�7 �6&�7\��<�6B�·	S�7��7@�6�+��{6� �B�ٵ$Qn��/���7��e4�5��`̈�4:�5�����5px}�:F�5�5"� �5���߃�w56�Ҭ����gĴ�˞��i�쮃��� 6u#��
�7�_�/)ҵ�m16V*6Pߏ�*琵�s��6͗ɶZ���B]6Qr�6�����p6D_�춓��}G�~S6�B6���6`���̶x�6,u�4C�7���6�	�������H'6Lg�6��6��5�y�?�o�,�$6�[��A�4��K64FصZ������|�A&�;3�6����~�5�1T61>y���36���57���6�`G�N�"�{�?��ߡ�ฟ6��6�c6���6x��6�gV6���5��Q5��T�WH�6z���T�E6,f���f�6��	���7阨5�uV5���3�$�,�6�Q6  ���I6(ǶK�U7�|�య4 ��68�J6���5fP�6j���5,4�6�� 5d7$�Z6��H7:�K6��6�x�6�X�6䋜��t�6�`���l7�X��׃7�͈5�;7���>���"��Ͷ�R$�����~,�����F��^5��n��60�(5~���&3d��Z]�x��5�6M6`I�5�� )޴�_f���7��Ӵ�.7haL� y4�$״3-6//6�� H3�;�6��SZ�6h��Z��� ������86��ܢ5�r��;��e�����25��5l��5�ۣ���A��.�6f��ry��``¶�ʳ�W1�5�!���Zk��L
�k�5m����������P 6��1�♏��wڶ������&a>5~L��U!�N?ٶ��33�m�6�Y0��z��;6(2���5\��Bx�������!�5 `�R/5:j#��#��V�¶`*�H����6Я��A㶪�5�@��3�4��7�W���no7�R��׶P�ۅ7��7b�\6������t7��7�zB7<��5��V6�Z6��7�bʶ=J7�E�6z�6�;�6��ල'7 ��3�G�4�X��������5�m�5 ��4�����<� 퀶DXG5���T㘶Fn�5�+��42�����>�u�l��?���ꊶ��N��Wɶ��`��(�gL5]I�6Ԓ�6 �I�6�H;�5���6� � ��1�17��ܶ��`6l$�5|{�6oٻ��������6��m�X���:LŶY$!�$K�6��5�ʵ0���($�6_A�5T���:��6^�$6��s�`<5�`�`6�`1�.c�6����\%6��3�S׵t�Y�V�dv66H�,��à����5�\ȶ���6�b�Xq�52j�5�O27ׅ޶0���p��A��|l��'�f<6�\��ht���c���5i蘶B~��5M�6l��������5?K޶�u��bF7������������L6��^�����m�4I�6�-�6Ew5k	��d��T=6����!�40`5`~�5RX��z1�6�D���n���ȶ�������N��*���,�6`<7@%B6���t�5G�6�
� p��#������eK��
���j6�I6ŀ6�����y6���nr��8H��$�v�ex�6�*�5?��x9u6�P��FM<��ݶ���Jn���v78�	6�5�y��o��ҩ�6	`���`������7$K��5z6�'��q���(���丵V�Y� �ж�ʿ�y����6Bܡ�x�Q�H���.=6�� 6&D��{�6(㜵����K`6�;��Ϻ�FX����4�_U5��Z5\X�5ܣ��%���=4�@6ę�_|����G���837�D�6���6 Ot� �6�T�l��w�6o64(�(SҴo�	����6�"�6�&$���\�6J�!��d$��i��������6�jQ�"QF6�o6	��6�7� �0��5yv6���x1Q5rA�6̘�6n���y
��競����(�~5���4���DZH6�U���(���������D���0�5Pݏ4$��6����2;����I��|�6����5h6%j��L���uY�6��ӵ�p��!�*^�5 -%5�?�69�බ(�5�G���	�4���6���|l������6����L{�60���l��6_Vp��i�5x)�5<��x^�6�дF�f�\k���2��˂5l��I26��5[�M6 �5*l)6]�5��W��I�6��5�S"�@��4f$���6j���ݶ��>�VF�5i���2"�6��
4W56�����{�61��6O�6H��5�Q����6|:�5�W6��F5�x3�
㶔{�<͵	ж���4�j�5IK��J����b���Զ��d��ƣ6��4���4��7��]�?.����5��F7"妷��b7�蠶�cy��+[7�k�7�QV��;87��5����6|���(�@*�p�7�z�66����K7��u��L���a�@sz7�jW3R�v7x��6+�����6���68��4�Oo��� �Ll�Q<��߀E�h����������;�7Su17|�t�1�D6��7=���Q7�FY���v�ZN���7j�rf_�z�u7�$^���-6Nؖ7�3����)7U���U� ���]5ֶb���Ե�ϸ6���`�84�g���6rW~�t.��̞�\�-���g��]����A�ö܅	��w��Rf6�w6J��t-��h}.4�j�0�K�h�X5��L�K�06���
*6P4�6T,5h�6�|��'
��8.�5(6�$+6 ��2���K��T�6L"ص_0�5�$>�5.���76�^�6n��10Զ���BQƶ����2%\5VG�5�˧������\6�-��1���k6� ��"��58\s6
���I�ŶS�6��3��,6N�6��f����5���5�����KpU��m^6\�X6P�|/]6AD4�\�`+����������N6l��6��d�495�����i�4�,ٵ�lI6��ȵJ�V��/��b
�5Ȓ��NȵTA��U69|H��h6�õ8�k��7�X6���T�7�t�5� �8�%����6<x5���2�5*-7�G��$�5X�����@P�6����
Y.���2�B1,6�I��8ʵpM��#@��V�6N�dٗ60��4P���6�
���5H�\6�����%��6�6���,6 ȴ(������5��m2j��50�ȴ��j���O�k661��6�r.�b3�5���66ֶ�	�(6����5Z��6�T,6��>6�d�� �۵I��&1�����6H��1U�ȃ 6.$����L��q��\57���8 -6�ڎ��䦶p�q4�ۅ5�䄶���7aj�6)En6!�J� G�5w�X�vK}�T�5����
7T$�6�n�qQ7���H�X5~ֶ�؜6Vݐ�l���-6�wj������?�60`5�D�� Ժ�Pg,����6����5'�6�Fi�dq�6y��6 �6*R�5�F�5.����b6�'��g4�ZE�6I��6@�!� ��PD��`f5����g+6�[=6K�5��U�u���<�W6�S�Lg�6�t9�ޟG6�U_���3�T�5��6�,��Z�9o:7D~u6�Ӷ2>6t.�� �Ƶ��6���6���6�c��~n����5{\6]��hpE6{��D6�,6�*�kE�,����j
7�V6���5���2�"-��#�6�u��}8e�7	8O�8��g8�7Ʒ2-8�̧�[�%8�����7�r�J:8��+8^7V7��7�?T8��
��8�2�7�{�7H�6��M��g�6��\��2��/P7"?�N&�7�е-��ш87x���3 7}�϶�"�6�&��JY67X��6���5I��6tf�7@I�4~Y�7x�T��➵��]7��c7� �6�4	8��6�5�:��6k���Y:�0����Q������퓷2��6�L�4	��u�6�_�4�@ѷ�y7�٩�
"��i��x����׶̡@6���7�2��9�7�8�7����6�`d� ˩�Z޽�h� �5>��b`7�E7i�D�.�˶Աu7�l�[��6 �϶��6�e�����������4����,㐷�g�7�`��2��c�ж�
��r���p�7��ݷ��޵��
tG7�z?��F���?.��O;���4�Q��ܟ?7�J�R�M�!􅷨�0�'��6ߨN7{�Α�74@�5���4���7l#�6W~���_17���5怽7���7
�;7��Ķ��97��7��6�6*���6��7��ŵ�6(�R6��x7όB��V��u��7�Z̶���7p4b�K�8�?/�����Xi7|պ7`��5�7��g7֚6w)�7����j���;7��<��s�6���7�\w��D�7x�����5t^(���74��q�5��q7�� 2}�҈7���6ڌS7�+7���H65�7\�O|7���j��55J�7s7�\I7h7	��}76�+��^�7���74zm��>u7�"�5�6�(u����5L:}6�,K7� I6Ą;� U7��6�m$7P޵�Q+7�7@�&4�O�5� �6���6f�@�X4dj�L)7��7���`��&��������d�w���Z��`�6��k��u�X�\7_?��0g6�ն�乞6j�;��Tض��׵�ݚ6���4�U�ꢊ7<���l��71d7&ն��ķ��8��M���&�ҧ��Tn�6蹕�B�⶞�P��˷���uZ.�x9������~��^�C���ٖ�7��-a���7��S��7tz8|HB��&�6���|�&7����Zs��$Ѵ����ȑ��5YV�����X�6.��4��6�1��c��X�7k�7��6x⻵.�7 ���68��7
�����^������Y6,��,�t�x=�,֘7��w���ط���g���]L��٦��X�ߜ�7L����f���e	��y�4dY7tq�j7�?��D���7z7pz\6pY�_�7����Z�6�q�6���6n�7���7T̶��+7�<��@�"��67��27����Ġ�62�6h��"�7�0q��-����7\�"�"��7�7༎�=��7(��5��8�Ғ���Y7�A�|��6�|�7�8��6R��7"�:�o�7O"7���7S�q�7޵�7j�)6|������7�F�7�R�7H[8H/�Dy7(^�5s�-8�wT7"Q�7X�"7�8��`7��84��7v%�7w���n'8�I7�#8b*�q7k8jg̵�
�7�� ��y�6@;`4��.6"���"�6䁴�H�f7:)��e��6������7}D�L7xz���Rf7���6��5K5�0,=7��A7�z���輷H�U�!���\6�����t����0���� F��M7>�ط	8�6�'~��&��e�@nJ�xʷ�e�.,Ƿ�.b6��-��47�ڷ CC� ms����6�[���ƺ6r"���F��EX����b�綼XB�p�56V-����W���QE�ao�$�� %Q�(A2�Q�n���7�3з��k7X�W��G7�:�@�4p�-6 �o�A�?7p�����7s=7����`i7�I[69�7�A5��[��m�5��0��/7�C�6ya��)7��2����6�_27 7��gw�Us07��7�_���6��_5�}L7a��7��7���6ǲ_��;�����7lN7p�ڶ&�6h�17kq���7 �x���7Թ׶!�7^�>7@.�5v�-�,T5w�7|Y7���7�Y���Ŷ�+G�R��U�'?,6hJµ���x���?�1"���.���-�L91��"d�`��5�u�7��q��6�q]���6k�S7�����h7V
B��c�6,%��h�Y�8z���6UΖ6T*7���L;��Eq�@h���)�E�8�b�Ï?��ȶHWZ7�D�6	5ڶ�.���"66ሷ�<3��H�`f�2f�����"7��4�Ey�7�+��\6/���u!6
RQ�n:�7
�z�`96�ݵ�Z*7q�F��W�8�"��q����·g�8�"���ȵ+�_���䋶�;6��7<�����6.�h7.�\��h�H�6$�6�'6z#Y7h<�6��6qn�7���64X�|�O�� e���е�v6PK�gHL  L  PK                     4 checkpoint/data/40FB0 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��@q�@0e�@u܅@��@n��@?d@1��@@��@}�{@���@�`�@m!�@{̅@L�@�ы@AS�@�Ɋ@m�@� �@F��@�?�@2��@-~@M6�@�Ǉ@��@͵�@o��@��@�@���@��|@!�@V@�ˋ@g!�@���@rf�@S �@灂@�v@�b�@�:�@���@�v�@���@���@
e�@|9�@i0�@0��@��@)��@L��@�}�@Ê@�F|@���@�*�@���@�z�@z@[$x@���@�@/��@u
�@��@���@$0|@�=�@���@C��@��|@�\�@ɗ�@���@�&�@�e�@T��@e�@e��@ؕ�@Y�y@�4}@��@�N�@
�@"/�@��@M�@�@�.�@��@��@)*�@ �~@(�@U[�@v�@:u�@lz@��@���@_��@ٍ@hۅ@)�@+��@!�@F�@$G�@�Ӊ@��@���@;L�@�x�@ؚ�@\B�@Em�@�͉@���@�߁@���@��@ Ί@䕇@O��@'4�@F�@q��@5�@���@ق@?#�@߆@	��@�t@*��@[��@8�@���@��@�с@,`�@`�s@�ǂ@�W�@?�@-A~@u �@�̋@�~�@���@��@9�@㾂@8ӈ@���@Q`|@W�@Gm�@ɥ�@HI�@+��@���@�`�@gހ@s��@���@�.�@���@���@��@|Q�@�.|@
�|@��@�É@�k�@d��@�[�@
v�@_�@���@c�@~�{@�s�@)��@o�@��@�b�@&�@Z
�@��}@�'@D��@�g|@@_�@�&�@���@���@Ň�@zY�@ ��@ܙ�@F_�@9�z@@�{@���@zt�@2�@ȅ@Y�@|E�@i;�@�q}@�T�@,�@磊@��@ꭊ@�-�@�(�@��@^Ë@�#�@�r�@�ƃ@��@�~@@�@
�@���@���@��@���@9+�@,n�@r3�@*�@�Y�@=�@��@u	�@|L�@[h�@�}�@t~@���@~݁@��@�Nm@M�@my�@7gx@~��@=��@��@�܊@���@h��@4�@H��@?}}@��@y��@$�@<��@:��@_��@���@"߀@�[�@1ي@�ۄ@���@�w�@�4�@g�@*qr@���@��~@i��@'�@�@�m�@^�y@��|@�~�@�=s@d
�@
�@H�@9�@�'t@���@��@P�q@�1�@y�@��@�U�@�z@�p}@)6�@}}@f��@"'�@�{@�x@�a�@ݢ�@���@aV}@�E�@#�@ �@tt�@���@�@�d�@�U�@�"�@���@�n�@���@�ω@�،@B�@1�@�f�@�@�y�@r^�@}m�@���@���@�Z�@��r@5��@��@�߅@� �@���@�(�@/w�@��@���@e΄@�ߋ@]��@*�@�7�@�@4�@��@A؅@��@��@H\�@b�@T׈@#�@�P�@
Ȑ@� �@.U�@�M�@��@>��@f��@8��@�؆@Z��@\�@�ۆ@�V�@ф@�Gy@n�@ -�@V�@$��@o�@���@8z�@p�@Fޅ@��@�݉@x��@��@�Sz@��u@�2�@`{�@g�@�9�@6�@�K�@��o@;�q@�(�@���@�T{@*��@`�@�n�@!�@h�n@�	�@&x{@�&�@�>�@���@-��@�
�@�@Ю�@�	�@5$�@�e�@��u@ <~@�y�@�S�@^��@���@��@�j�@�k@e;�@퇈@�Ƈ@�6�@o��@B��@M��@%��@�rz@�^�@}�@]��@H�{@�)�@�h�@��@��@�@�7|@0 �@��@���@��|@j�k@�p�@�*�@���@d?�@	1w@[��@��@�y@dp�@�"�@���@�8�@+�@�ˍ@毄@hV�@�@�
�@At�@�&|@*�@&A�@��@��@�ׄ@J|z@� �@��t@/X�@�o�@�x�@`�@�2�@��@	p@�T�@�R�@J#�@y9�@�x�@�v�@�	�@�y�@PKl���  �  PK                     0 checkpoint/data/41FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ��?�@.?�(>(W��>P��d4�x��!�m>�O��P� ���I1?-��=D�	?����h='X�<�հ����*o���N�%�n`��7��>��L?��=Ⱦ�>��>5F�>4����9O?�yv���"?f|���>�>Q�?C"�>����O���si>4L⽧����W=ͱ�>i�ԼS^m?�>��,?<�?:Ι�5u#?��:>;!�	��>�o�>lE6���"k�7��t�>x��>61?���-�+���x�sJV���ʾ�b�=��-�A�=�\>?��?��*=# ?k6=��?Σ-�ޝV?��8>|�_=�����R3�̆h�W�E?/^�=�v龦��o}�9��ݾ�u?] 8��$V�;�Ҿ�Ɋ>�Z���4���)=_~�Γ_�/��=7��>y<2>��<�=�{E��+�;m�C��L>��=j5��P�������vF?�݌�}+>`��,����O>�}�>_�Ծ�ɝ���#?/7�=���=�U����4��*���j.>���>˲�����>�_�uW;?=��ӝ�>	�>s� >��>�F8��l?\]����%��h�嵦��F}�)df�fR%��s�>rQ�>tB��`	��g�>�= �g���C�?�,�/�>������?/���	�ý(�G�T�E��c>����l?U�(?�˄�]>y�?n/>]/?đ����?�H0��c?�@>� �D��>�F>�7�>��G>�=7�&�7P=+S�s���0>]��7�?��R�p���>kR?�H&?*la���N?������?�7�?�?�>Ũ�>�1?�+��澯QM��>K�-��� >��"�G�G>��վ�����>�F=>�/1?<$��!�Z�?�Ⱦ�-�=L������U�O+��c���%�>9 ?��?�x�>f?��@�\��>��;��>c���Gl�9�E?	;5���L�"�X>����R!��9�8�.>D�?���64����>�ㇿ�I?��0�?���Hb>?�?�$�>��J>�����<�=��v8 �>�*?k�t>n���i�����,�%ML?��tH���/|�V��>�E�4Rn>�����T?SK�>f�;?9�h>�E/?D0���>"V�>��r?ē�=Yl�46��e�?�*h�kad=�?(�|��H�����A? z?09���W?�I�>�?׭g�&�>�*�=�d�¥N?A���I$�U�9��3)?Т�>S������>!C?�ea�E	�>j6��˯>UA'?]ҏ>�N��ۡ?����,�9
?J�%����'?]�-����
4���?���i~߽Sn��¨��4g�>!+?���>n�����ҽ�?�>p��=r�>�w��s��������C?�E�=4˴>�
?		*?	n����,��վ)^>��Q>��?��d>���E%�>` 뾃:����:��q>�?>�U��t('�/XR>8m½���>�c���ڻ����>�_ؼ��ؾ�,O��Fu�?"�>ͬu?��ξ�ǽ�e�=�!?�Qg���?��C�)Y�>����1�����b�a7?q?�����<������V�=�55?��>��T��F���eI�B8C�Z>>e��|�G�n�=?do��J��Q�>Q#����x�զG?�Q>{߾���`�}��Ѐ��fs��U�/?3���u�>�T��>�����x>�d<����	?�d�%Z>�' ����>��t�.�(����WP!?�C=L�>ڡ��j�2�c�>M���8?���>��8�xI0>ˉ�S�$�j#?���XZ?�O0?��?�]սw�4?���,l�-����,?S�����Y��CW?I��u	>��>n�ɾ�?t���am>R��>�]?�H�>�n�>���U����־X[澎+&?W���{�I���>?t@G?{@���?wJ�>P�����D>?(��yn~���8>Q�m>,�a͚>PKP+���  �  PK                     0 checkpoint/data/42FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ>Sa;��N>Ll��G>��ƽ?�!=�s=>�;3��ꑼ!A�<�,��$N�R��,��<��V>^��=L��K'+>�]�����=C%���9����<�,��q�>8��=��>���>��Ѿa?
=�I��>�4�,Pþ��սՎl>
{��y�(z
=��k�Gb����>f�>b'5==t>�[ >Aぽ�>	;P>v���#���i|<ظe��{�=ͨ׽�>WcX������������-޽��U��� ��6 ��r�>΃9>�ѥ�$e<��ƽ�b�>�{�<<���ś���D\>�X>O����>z{�0�۽h�eBs�����S4��a~��9�;�݈������V�,���)�m�^!>I�<���=2�@=�
>|�ܽ���p�j=+�o��2ͼ��>�ޠ=ۏw��D'�/e�>��>�c>"�ʽ��P=�N�=�\�=b6>�ɾ"dp=��P>BG=�5��	 ���%����<�Y�R�!=+�/��R׾?/=���c� ���n>�e��mTF>�3�=6�̼�
&>�~>�Yz�cA>����y���1�M>�A�O,H=�ۡ��@)�V�����=�v���қ>���귶�ZQ�>pI>��!�>�<Q�<���>@L�>�T>�u�=O��>�����%���v�#�>�y�= ��=1B���>��ž%�<�¹>��<=Ҥ>��C>����ɾ��l��"�=4�d=ͭ����������ˡ����E����?W�7�]�>e�B�|�e�[#�_�J��{(�a��=��G>�>l��������~��C�'�7��Z7� ��ɲ���z�>�;�>�Y�ɹ�f4X=�廆F\�5���J�ֽ���I_>�N>��P�p��K���T<]��7��5Ҋ����=�3-=���>��>�B���T=a�h>r��>���}�M��s�<�K\��S>��=��;���S>w:�>xX�>��=>��=3,z�/�>�c/=�V>pf�>]1�������>��>����ЍR>��>��=�"� )�=�>�kx>]6Q���>�	�>�m�n"q>ZkN�O��=�> ��>G(��d�=��ھ����M�>tr��y=�D>�y��it�EF���3>/W��k��=29������R>�`����>oL�=�X_>G�9>�pU>�]ƽelK>�{�C�V��F��8�#�X�$����>�$>rr��i��E�OZ>UM�>���s��"�=�@����=��4��C<.�g���3����>k*F>C��>�1-�wZ�=Ցf�\�T�%bh�]�>�0&�e򽬃��K����P+>��>{�>�����:9>���<:�>�I=nH����D�)����Y��=�_=�Ȕ=)�A�X��:t�> b�0�X='�>�Ͻ�{m=�(׽،u��н�����R��r|��V>�>�Ҫ>�t`>i�˾�z>��c�����U-n>�8<��=���9Fo>�:�>��b�8�Jc�>g�>�o���>Q��<�c>>*%�>	/�>�����!'>!�ʾIfI=9�>×��y��>�hx>���|�k�Ҥ���>#�_<��K>�o�=��i=j��;X�-�j(�>hH>l�|��H�����RU3=5@����jJ =��^>_	S���=���="X�=�����g�=�W���������>[#$>�w�����<
`��}���@��yO�[�8=O�/�߷�R���j<A��=O�g�9�|>����/|>�<����F���.�::c>�n��ʻ>��<��	�o;=�K5=/�]=h��=Q�Ǿ+�� �)>2��=_��=Bkd�|Mj�
�P<oo��976��'��`������K�`b�=�_��^����<��*���4����=}g�>���=�X��6�>C��8*==A=�׌>��v<��˼m��>��1W�d�L>��>��p�R�/>����u ���6>T���t�=�����*>�l=�b�>Uy��f�>X�>�l��eK�>E$Ծ���=dfp>�8M�)��>���>�m��0��>���wœ�=>��^��>1�>���`�*���>�L��5׶>z}b>��0�==Ll+�b�ǽQ�`=c��Z��"�=g�6>�h�0gr>P>>�=�Y����\>O��_���(>V�&���������#>�ET���$>I�ڽ�`>LXk>cƾAr.�����*u��;�>U�I��Cq�Iũ><�>�Ϩ>�2a��"s=��V>.M������jx���ľ���� �Q4(�qS��%>��B�˚�������>��i=�E.�@���?8Z�	�=56>�6��a>u���e�%�]��>�v��B��@��>&�x�'f>��>��>K<�>	�W>���m�>V`>��Y�0����3�>m�=��S��`�>��=i�>����?^
>-���4�A�>Ab���}<��>�Q><t�>�p�=�V��Im���<ˍ��>��$��yQ>�����#=�3��;n>׼�>���=ʄ+���>gE>Θ�x:�>��<P�~�}�׽�$d��y&>�E�,0>�q;=�>�����ʽ�U򽰊��9��>-��.��><<�+�=Ko>�S>�,׾ǣ��]�>On>���>)�=^؇�����l�E��C7=�e�<}p<H�I�ڴ�=�0�>��/����M0���V��g�μj��>��>k�>��>1~`���G>.5>�I�>�m>���z�پ��>�IY��� �+�Žؽ+�诓�'0�>Ξ>�p�bm��w:�B�n�}q�>à>g�����F�F6��~M�<1����\>)ϲ���I�#>��x=uG����=r�=���=�9�Ӈ5�C|�>An7�X C�
x��qY>*�;q޶�d=����<�o>I�?�Ϯ���\�a�;0������C>U�$>l�w>�>�f�>����{�>#�;���m��>!*6���>���#�˾���>��
?l1a=t�������	�ƽ�4<?⇾�������Z
>��>�>�m�=�|>�(>31��[{R<��;)�ؽ������Y���ӽS#�8�N��0 ��Ϝ��\>���=���ky��y<[s۾Ac��e~>�K�/D�X�x>D1�;��<W����>��>�=� �>F�>BS���N=%Y��n!���ɸ=v��>.t>:��G��>��U�v��=v��O��>f�L���>���k�=�R��W���]Z��^�>�uh�t>��y��֫>��/�Eq3>C22�V{�>_{�>�2<�J�=>4N>�M���Ͼ�U�>���=��r=4�=N��=���)�=
��>ꨉ<̈�z��>%�6�"g�����"��\pѽKY�je}>q���p >}��>��]>��>�M�=l->,�����=�O>�Dľ:|����;�2����B��$8�g;����P��^��{�=z�W�E>\���9zY���x���McI��5�����r���M�<��U:>�ɣ��Y�q�1�u�6>/)0>s�����u��	0>��;>�-�o���f��9f6���q�#C�>�rs��f?>dms��c=�<>X>,c/>�VK��yG>:$[>T�5�m��=c�>.��2۽�}���4��TO<X1|<������>E�f>ӝ�>B(>�V�=4�0>h =7(w�U�;>�F�>��k��d�>G�S��MB��L)>��Ҽ%B��Dֳ� '>}#�������Ѷ<N�{T��c��7M��t5�qJ#>JwU���+�-0��žҘ�>c��=�=}�μіl>�̹��+,>��z>y��<P�\���m����>�J>�8�y�4>�ݽ��P����pg>z~��u�f=��\���2� �諍>��-��cU�c���ї��X=�٪>{�B=�܁�8�>>������>���>=Iۼ%D�=K�n}$���K�G�t=8uI=t���r����Ύ�+D�>Q�>�	�>?�9�ϡ����>�����A>�=,��=�nh�<|ͽ��X>X��>�$>{�P>zZ�>��>������;hV=�7�<ޟ�=���=g�@=�U�����8�='"�<ȅ����=��=e��=��z����=YnZ��1e�E>�}�]U����<�D!>A��<���<��_�t�>��/����_xJ��>΋��W�������p=(iԽj���Z=��8-��̳=,k�=&~<yA�������5���@0�=�9��� �=0�#���ս}�:KJ��n�j�i�s��=Q��=��)>�Q,�\��od�>���^n���}�<9��<�`��n�_�a5�=EV4���.>�.<��4F��^)>���1}�=`��=��<���:�<�>g_�=ܷ�8�W��������;�㮽������4=ˆ�=)�<�	ν-��<ss>N}Q��u$���>$:=x|'=�x�ND���<�!>1�=l��=(>w��=�^l�$W�����3�=�SH>�0�����M!>)�=6���7=�Y����Z<�:�=�l,�~~�<�#�<$a��}$�9Bw>1!�>/d��t,��;�4>�eؼa �v|>���l<�k:>�Ƥ�'bȽ���D�$���ɼ@�?=��=KVS>̼�g,>j�Y��o�=�.l��]�h���w�.�Q[ܽ�Uv;��=����>�M��ȩ<vR����<Xt=7�)<���<'��>�?�s����:�>�߁>�й���F>?�t=*��=�,�=p����_�[��K��.�}<�E<�Z �Ğ�b�!�e�S>g�w���-�(���ڼ7������=#>�=pU�=>�< [�4�j>����[��=�:�;�Ο���=9��l���`���"=��%>��!��̤�6���>�zH���%=��>#h+>ƿ����=��m�����J�i��v�<�^7��� ��Ns�{2�=b]U=gY'>��=q_1�z�=�e<.[=#G>%}�<�"8�p���.���2�5_"��=B<@5>�ac��ea=a�ؽ ��=>"WU=��3=���=�;B�,;=<�>t�F;��u=n�>�������=/���K<-J��Q ����=��4>d���F-j>�焾,i?�K>���=�)>[�>�=�=XW�������'>��>�;9�>n]��=b&>:\=r�L>���P���+��6#>�#4�6Y�=�ܗ�8;�=�����ĽɄ�>tHR�n�(>�8C�K\۽W�¼u�-��TG<i=��W>�-��	���+h���>GC=�}M�=Վ�=
��<�܂=�k >�Г=�7R���=sA=�mY=�-�=K�>�Č=̄�o���F�=׽��=i/��
9�>vN�=���EY��'�<4�o����<��w>��<v#=!0�=T����h=G=D�������?M�<Y�=z�6�>qB�mR��r����|��?p>�r>�A���k����I=Y��>�1K>�=)�x��?=�I,=��<�5>�\|=��=	����&N=���B�޼k�U�5� >i	>�,��|���MyP=V*�`����Y&� �d=Q2�<K���;a >�	����=V4��9v���?��Y;�P=E��<;R> #�AU�=o��<�?�=�X*>lq�=�oB��S��[�=)�D>�Y?���:�E�
>���5>�RE>�K�<d��>�c=0l���f�$p=��=K�O*��Q�=�F(�HS��w�簬<��x�U�h��j��0�=��+��2d��� �ex�;r��=}� >�I_=(>,2R:,��=7b�[��<&j>���={7>pCB��ӛ����=p]_>w�(�M9���=׽Z ;=�w��ȟ��9%>�9���!�<r�����=�"�=�3R=���#�ʽ$�@=�-1>�:н��/�X� >d�<BռS�W�-Qf�G��sO�k��Ľ��>���M�;�@�<3��=_` ��&>���{M�=�^l>� �H �=tT��b��+>��Ƚ;H<����Y;2Z�z6�>ӯ�>�dO>������F��7�=$����Y�<���<�44>��>��>`R�=�R�;�!>��(>�>�=���|)��~��>h�=�j�=H㠻��. K�	�>z��h�ڽ�P�=U����>�����	5��{���E��8��;�t�g�e�=��E���"�<�������A>	$��F��=Be�5�=�i�<�f�no�D]��̕��zi>�%��9:=�X>����Ay_>>������~�=��/>�f>�����<����E���|%�*��<�i>S���QS>U:I��N�=9�o��
��'�~��>�J��M�>�R꽟e�=E�W�=0�>o�<c��<y����3��5V����k=�kS��9��M�Z>��B>G^�>�&ɼ�lx���G��)�;�&=��K>]�>x�N��+��n��<p\>�\���r>�3�>O�����>��r>��>�pU$�=p�:�^�<�fv>�d1��Sk��}�Anp>�뽊6�>|�Ⱦ[�J>����%��u>�P��u��4>��|���>��<ZEs>�Z@=�񴽨�ŽK�ҽo�վi� >�l�>�������v׽A�>D�x=7E���[=N �<k9]�t�9=A��=�G�<=�b>�k�>��/>�(��$=]\g�b9=�z����X�J&�����	�=�v>����P�k>Q'����=IL=)��=�^=\v��� ���Ζ<�>P`�:�}1�aB��+蟾�I�<Hh>u�A�Y�2���=�^=_=0��<;��=����==�/�<gJ����=��$=c���>Y��U�(�=[Rq�n�5���c�A�Z��>��s��\4���V����m^��o�=�x�dE=N8=縗�fP��̸=�qǽ�y�k��ki����=�*��<@�L=�C:�ϊ=��n>��ѽ�s>XW���=�8�|;
��r�>��)>3W>=D$u=����Q�y�ƽ�i�<�/;���S�O!���>����V<��C��"�>�|
����Ԡ�>6y�=������k�i�>y3>��f���x>�"=�>q��O����>�v.��-�=�M���8��J-�>�^Ѽ[��cݓ<�]�(�vW>q��
$�a#>�3��m>;���5�;��=�J�>m�ݽ�$��� >���=�)���R�=p�������eD�#�40=>S>81Ѿ�=#�-�p�'���>9J�=��>z	�>�v�>	-ѽN\=�%�V ��E>�Ј�磵��� >�O=�1>�:�>*�5�5����
���S�=PhD:�m�-�b>_Of=u��=13=�1#>���=#��%�����S>�����1��C>��a>�������U"�=���>� ۽�`Ҽ �># Y=P�!���=oF���2�.���=��>������=���=f�;L޳9![R���=�x���s>wv)= k�����>���@�<{r�=��]=��8=!�:>��>L�'Ē��L�����=��A=�n�<-*׽�S�>��Ľ=.�:G�>�;{��t4���`����=��h��+v� �F>T�#�2홽V|�@��<;ゼ������<�Y�2��O��<dA=��^���=wό>���=� 
>:�d>q8��P.���Ƚ��=s���#�_�<�>LBC�1S#��=���=M5%�eo<�(]���A����=��>�~f>�`Q>����z>a�>��;�RR��� >����t>1��p9>Z��=��]=;нv�W�j�B=(�뼰�����*�ڱ`>��>��B>!lZ; z�>�臽��C�f�I>�����=���>����?3��J>Ņ�������>_t<��=>�s�_K��!=���[>aJ�=Y���{�^R>���^�W��K]=�)s�F�f�"�z�'{�>@��QPi���7�UMս�k)>f#d��r�=Bܓ>ؼ��i�>�Ch=_޽��>#�L�&gʾ�t>�Ԅ��G�<&>�>��  >SO>[T��Eӽ=�!���`�j���BI>����6�r�1�Ƽ[Mὶ�>X�=�����,S�=��=qu�A�c�&ռ=٣�<j7�	����E�C�Z����=	��ݜ�<��>��>�����#>�E��m�L>��Aq�*�q>8F�>&�&�K�Y>$wF:3[����i���ܽo�� �=1��>_	��1h>|<r;��>r�{�.Z�+��>4�>�+���+�?>���U!�>�%�����_�=h�)=�>ֹ@��b���b��d���¾ޒ>��Y��+��T.��FR��w���]>--�>(=
=��=57ý9f�>kT�<��Q��2>ҕ/>Ɇ�=����ԽX)�=�j��1D>UU8>I�.>��y��渽���P�e=��=�mv���ʽۙ>�ս��>a����/S��߀��Z����<��<�܆>��&��>���A��v�:�;L��u�7>~O��t.�>6��=�����+>�qݽs*�>�`��q�w�3��=�e�=��<�3�}S}��*ֽ�MľW{ �U4!�p��>��=�����n>�;�&�r=�lȽҞ�>���>�C�:�a=hS��!�=�K;>c�y��S)����y����/>	�(<�����><#y,��.?=�>q<��C0=�%���< �>�����P=�搾�Y6>4P�:�Y��y�<�>���>�,¼B���&��&)<�E��>5��<��w>�?��ܡ>�T�@m׼�l�=�͘�VM�<�g��[j=Us����&��Z#�8_T����>�����u=��N�o�z��EL>瑥����=n�Q>��z=�M|����>��d>�e�=p�j��a�I�A=��>;f���=D�"�!9�=�0���>��~�"ʔ>��c�a�h��M>�	>�e�=�!�>�?3>�Ӽ��6���D> x�><\��+'ž�=˯]>ռ�=�#�����<�{Y�-
>E�����I=�+>W��>@��>	�x�w�߾��=:R�=��=7PD=!�>��
���������eD�=S0t�R�n>��=��s>y6!>�e>ҺW����<r#s>������]�M�>+A�t�h>G�0<`�<�=�f�>x�޽�=_��=���=&��]'�=�)�=��?��4�=Z=�T>ʍ����jC&>yk�=Pt������0>]�s��=⓴�d�=�r4=�?�=avg>��=?�>�):>�J>��=�B>�;�ӽ�>�s(�i:�=���=�&��R5>HI6��A�=dH���L>��=��a�����BN=k�o��a��dz>�i�޴�=�a�>}W->�>Dܜ� ���"4 ����>�=f�= � ��,>�à>�L<>��<�3N<�r޽�+1�L>>XQ���-��TxT>�/�� �=e��>L�>�>.�j���`�Ʈڽ]i�
؀>^L>}�==�m�=n��= �-�+��=a�k>�8�]�N�D��=><->��5>9>��R�ݕ5>��n>W)C�h�����=�w�=�A=�o�����B>�m�;�?s�C3.=G ���=��A��>>��� �E=�H�=!�>��ľ�M�>Wn�wK����U=��#���>����Z>ǘ�=ۨ�=�K9>�Wk=-L=�X�>wW��3{ͽ6:���<����Ŭ[=5�<ܱ6��~;����<����Eɽ�Z��ٻ=�xk�d�,>x��>혱��|k=���>!�@���|��.��(���\�>�KH�N2��M=D�a>�~W�2�+�î
�����̊
>���_�y�F�Z>��S>�aB�iS�,�*>4\�Q9��f[=�>�@���=�K�W� �)��=���>u��rD>���j�=�&=�Gt�^�5�&<���|��Ԫ>��>��>鞔��㕽1=�Qً>#=n>}�{>}�O>��>�����Q�F>��>����Gc��8�)]��\^��3>���=	!���:9����v�U��A�=+�[> ����Z>��!�<��<Y+q�Y)5���=�� �h�j=˪�>_�$<Yh�=��<�U�;D�x�?Ͻ�=�[��~���ޫ�����-�����=Ē/>��̽�S�=Z����=�Y��[�Q'm���.>%E����"�k<� �4��kH�voe��q>
ˬ���:=��(�����B�*7�>�>>A=A�ܹ�b��=̋�>�q@��?(�x�=~ǽ��f��@X��F�8u�wn�;�א>07>��F>kM����<~�4>��,=�Y�A��=pe�:@^�n� �?�=>�N�f��<"�F�����w��h�{�	n��ul�>�(�R�=ׂ>�Y���_�=��V=Ų>>�l�eRۻ��=f�>y��=%�<#+e>vZ>h�={m��j%�=��|=�P�i�<�}C>&h	>+�>&-R��[>!�>4=>���ȥ=�LS>�.��#����u<ypf<E�ѽ��E>��Ͻh�T>W8����=#�=�)>�R=&a���<�e�;/_�wp潅SȾ���=��I��Z����"=��>���<��)���"r�=n�=�Q���<G]�=!�1>GO��!*�C᜾Ӽ��)����>�׻=mQ��z��>v��$M�a����=3ٰ<C0k>�i��n(���I
=�*>$y���x>G>��h���ý�u��0�=������c>0�z=J1>|{>*i�=.$�=q"�Hك��	�=&:���=��#=[)��9q=z��>W�ʻ�9�<�`"���=>�w-=��>N�,�@ס=6\�����<��=5;:(�l����B�H��˼����
�3��C<�� �̱>�������>���<��f�t7B����>&ý��>*�c�G>e�s>vT�<Uh>ޑ�;c���w�=->
�ڽ�PC�l �=�%��ko�>d�=#؛=aE��I.N���Ѻ�>A%�� ���������;xؽ=:�x>T��<��W��k����>�Oǽ�Q��%>��n=�*�=D���=4-q>k@I=w�V= ڀ<1�,=ӄ�>�.6�;�L>�gC��n�=a�O�vF�t�#>|�%�+�}��ې>���<���>�s��I� >U��=*��=��>�#>ڱF��Ĥ=�ϻ�#�	>��P˽xU�;+b��o[�<�0N>g�0�h�k��B��^��Mf=K�=>��s�>���=,�>��>�}Y:�z]>d��=�i�Z�>lIY>�w�<#9�?�����=f�Q����q_>k)>>�?�+��=�>���=���`�U�f!��� �̔���=�C��o����=��̽C�=�S����<D���a�b>A녽���j�=<�W=nP+���i��Ȩ���:_@ >�ؾry�=N��I���A��>UֽiZ;�lX>� m��)>u��<�v����@�n5X�H��;'n���/���Յ���l�,�l��e�=��R>�3x��f�0�T>͑�=;K��)����=����k��<vr7��k����2>)(?>p=��`>�'.����=?=%>���Tr��S�>Y�e=j땾�.$���	=��=S�:>A&8=��=mS>��`<�,����=�\/�-2����=t��=u�g>?R������y>��{��������=�ua>q�#�����7�
������C;%0���UX>�!C>}^2>P��W"�\#����t��!�=�y�򊁽�K&�y�	��,�<L�
>��=�I�=�>J��=�O���Rz;��|7�_��Q%>�N��t�>�Hm���Y���%>�1>>$����hF��f����>*�s��=�����ԽR�%���ܽ.Gp�������<
>}�;���o>��x>U��=V���T����>Hq⽍�	��b�J��=?f��\�{>�F�;[~k=Z�^=c/����:A����n�<?ʚ���7=_z�=�����8�β;���+=�Tu���p>��g�wq=dH�>���=b1/�A��=B��=�����=i6�>��=�M����)>�!J��*���S�N��=Rj&>z/t���þ�/F��@ʽp=�<��=������5�X��>¾j�k��=e��=6�����3<���tb�=I��O����<h�>=6d<���Wv��8 <�=%ט������}�=_�������>5ӳ�)��=��J�S��\�=ܠ�=V8]>_c>X*>��|�G>pT>��=@
\� Y�y��� � >B+�������Q��4�)�,������9>��i=���;�:�>�I=��~`�>�e���n=}%ν���=�\E��G���_�=4S�=�M����7�^!�>Ɩ�>{�e=�p\��¼C�=���J{��>띣��9���j�>@��=7�S>CV!����<��=��N>�ul>p�=�g�=e�E=�|�=��<=y�=Q�Ͻ;ƈ;n�>�_>ݸY=��<��]=pj������iH>is=��=l���s��K�l��]��Ҿ%H�����=V�뽰�>K��-Đ��������v�c������Y���5Z����d���=4��	�=C�X>��Ͻ[e�<�5m>$��N~p>?� ����<03%�&t����=��=SpP��G*>���=�M>�a��=)֏=}��*�=Nf9= VM>�v�C�5����+�����<��ټ�V�ʀ"�TYQ�����2>>^6�1��=�9���˽�^>���<���=L|���5��Q>�9���X���W�P�y�X�>��j�1���֟���>��>�����=��&�������1��d���f,=C�^>�(K>�*�I�����c4Z�"�c>���=��~�k�ܽ����Az�;�M�=�����\>� �>x!<���"n����>xͨ�2>eh����½��<��V��!z�]���Ǚ=�f
��7������f�<�(�;V:�>=u������"=��P=�K��+�m|���N=���[Y�<��T����Aݴ>��&�o�{��>j<K7���Q�=u>�t��nƻ��g�o˭���;dT�>�W��<���Һ�Ⲽ�ξ�l<�$��>3&�=g$���|=Ӱ�"U�<�$n>3_P>*�=�O�4�N��0��]2=I���/��)����x>V�9��9W��q>?����Z���;ɰ~�gq0����=#l"=�d�����=��Z<�%=�W�=f�q>�W>F��g��>�*�=�#�=�:=Yܘ���B���=O_�=��U%�>{끽�����_���W>�;9_�|�S:-�O��,�=��>�I7�dSD<D�C>q�����=9s8�� �zȾ��;�&9=Yq=�Z>2/�Y�D>&]F>|c��iP$�q5�=�>�?D��\[��\[>\6=>�>��:�\>�g*��qѽ��I����A�=L`켅�=�ڦ�U�u���r>�?$;��ý�+�=U�j��t�>��=3e$���I>��R>D�7<-��� >ST�=�����4Z�]�x�]s����#>�=>V��
$���⽑��=� >�1�����>~�����0;�P,��S>|즽��ӽ�Qv>��	>{�<�c#�1%�V|�<��C>�kz���>z�V�B��[>:�)�=%| ��g�L�>=�V<��ǽ��S>�=�N���=О�<�U�=��c<���=�넾H��y?=�B��7���-��=k�*>�ō�=��<��q�����w��� �p�>p�C�3�\>�|�=�!��8�Y���>��=��k>������Ͻ�A>�ů=wvʾ�>��T��f��������v���o��쐾�%�bPI>�
!<��k���>��K�>�M�=t���� �I?,���=��>8��=�$3>�f�<?f�>E�� K=��<ç�<UXY�e��>_F >��@����׈��"���&�t=y�=� �=��M�Pz>��x����SW�=�䚾�����P=Y=�W�
�I=�n����=��:|b*��*X�C�=ȝ��:�=l�Q>F�;�c�h���C�>�D�Қ>~@���g���.�J�I>���> �=�>i�=�O�><�o=�>{�h� j�W�X>\��+�=,^*��R�l�=	�ź�{���/,��$=G�;%�=���!Q�>�`�r�Ľ�~E�{#>�q�<��y����$��Ih-�%��<��e>t.�=�`��=�H�=�͘>���='9p�O���ۋ�J ���`I>��>qN�2�������e>/���R�=�qP���*��z3>�3o>/�u>��p����<K���e>`e�=GR�>�&=���=�%��~�=��J>u��=�>)�Խ��P>�ߓ=�~~�����j+->�e:>�}�����>}�c��~N��Pܼ�ݓ<�^��#�=��>�=��=Z�8>�k>g�:>�����P����h>Vf]��v�=3�=6�N>�dL=�iȾ�ez�O.>�x=����������.4>��j�u�]��=zս�L0ֽ�ݽgS�<��=�Y�� ��<I
ʽ5@��H�=���ט<��=�a=!�̽� �=��n�Zzd=%�<����)ֈ<�K/>���%=��"�~%���{ʽ/�F>����LE>u#>��<=�\\�<�����</������<X=	Q>�<��-$���3C�k^�=���&
���:=>�'P=�������֓�L�h��S�i��=_��>1?5=�츽�S>�]
�T(M>�?�>��>%)���=}󽦶�>�j��OZ>��n>{�*�����'�����꽍���F��~k�mL��-�=�o��>yɻ��#<�r>�/�-� �|������y�=�7<{�>���=��;C��>����pc?�R�-��;�>߯�=<�Z���ͼ��I���Y>%ٳ8��@��<!o�=vG����ѽ�o=��=�V��0��<c�)�Kx��2ֽ�Q>�E���Ľ{$��.�!=��B���<�Q9��'>�����>Q$E��?>���=��ɽ��򼽟>�tT�=v��i2�t���2>�-�=��:>3�>��*>r�>r� >�_������Jݼ/~p=�%�>�E�=���=!��}��5���_NV��*l��!'���;�B2�'EP���l�zj���^I� �,��lj>CBY���=�K�9#N��d�=z�=e��}6�PJ�iW��A�n�1C����Խ�~|=�.�s��=��ɽm!�=0��;����2ZF�@<��>�J�%��P>Z�%��ؤ�-�a:,�Ӽ���^�����轖���	
��/缯�޽������=wT>b�ӽowĽ�F>A�8>��`>9}�:B�1>�zC>I�>�Ē�wa��%ـ�"��=!����=��i
C>AZ	>=0�=�
T>oK�0+8��S<�I~�������=?�>a�X��:����m>$��;GLϽh�z�@�>>��=�/�G��ȶ�=K�v>���=���<���2M>`���&CU=�_��g>�$>���=��E>~�����=����N=�ϧ����������r==�t�,ߕ��`>��޽6�ýk�ӽ$̐��,��¾�]
�D+�������@=�ٶ=�)Ž� P�'"J>�!o������o>�=L����o>�W>*��=���=�h|=3-l>�=��>�T��BV��'��۽�>����<���j�>��>5�z�=�`��f��n������<Jc�>��=�̫���^�3��=K�K�'�=+��<�Dл�F�=i:@���>�A����a���C���=����FI���xk����>,��>�����Q>�G�<a���Z�X>��ƻ�=�m>�N�>O:=jO�<��=�nj���N���νY�>�w#��\>����8���0�ܴ�=4y=����	�W�����>���� �ǽX���f��=R6߽*E;�w+�������V=�E�Ή�=���c~���p�=�Z� �i��%�<>}��8��vǼq�l=
��'N>�)>-�P>؊�> �>�$�>˟�;�>cu��p��=b�=&�~>�P�=:w޽E">6��<��>A�ڽ^����<6�Ӽذ>�`���\�-���X
=;&W=of�=��_>��~���W���+>0����'���&�Ah>	��=��=�X<�DD�= �ֽ<|�<:>xD1�����_}���	<x�'�ǂ�=~��_p���<�y�<"�d>>8�>�AսG�����<��G��qW�?.F>D]�?AO>���!��eĴ�f棽�,(>�z߽�je>�ٽ;oὊ���
�;��2>�쐽��0>i��<'�=�o�=I��=�遼�9�=�bp>�A=����
�<%y�c��ִ�?}
=�=���5��Xs�AJ1>�3�>wT2> �P�U��=�V=���9uF��N���M
>*�ʽ9��=8t���`�=�����'<���<�Bѽ<>=w	�=�h<�2��.�>�'���=�^�=�g>��'�Z7�%�V���S�<����=�½>����=�+�=�xɾlt��>�P����"����=ݮ8��J\<�>�[�=���=G���3G=s��=�E����e="�\<���#D>�"�={d�=7��W�=q!:��~ŽL�=I�����y���O>����>�|J���<ݻ���_>�ļ} =I�;e�#!,�-�	�0��GI=���>5� >��>L�b=���	��=WB�=���r�B�FWH>�ӄ���^��>�� CN<*]!>V�罺r=Mh5>4I�Sgz=j `>�	�=��(��T�=?�h��0_�2}�=�0y=��=>� �;�_��!d������:������<Qw>��>�cb=F�,��Ê��M�>Rx<�^�>��v��o�>�<�=&�s�t���p�{�I;R�<�0F�+��bAD��_𽸺I=�g�<%�[���'�ZrU>[d�;�3ҽ�`<d�<�#R=�պ=ʹ
�!M�=��c=���.f6>��0cT=�ٽ�� ��+=�=��ƽ<:+�p�X;V<��>���c>@w>��=���M��>'/>H�/>�XR����=�](��g�=6�i���,=�!�=��K��)�=�W <�'����/>G��D�Tp�<��K=w�>��$�h�3>�k=�R >��d=T����� �Qၽ�o��G��=�ͺ
_�=� ��Yû��j����Y��;��2����=綅>y�d>���=�ϙ=� ���	>��\��	�=�F>�����;���}v\� ��=B��Z�[,"<��=U��<�N=Ϳ=ң>b���r:$��p�v��=Q�>�瀽��y�ti�U�6����=�<=����dG������Ai��)��B a>�p��;�r�6�9<�0>8k�;��(>_f�<	b=��8�������=?I⼑e>�y�>��K=#_>�u�N�Ľ�1��I> ��=�c�<�D�=?l�=��*�wd8=�Y&>Ξ�=��6=	yt�.��=
h=EqB=������=�J�<�5
�u��>���w��=���'r������<�� <k=�=�����c��c�Ž������6�Z=<�ue=��<߬=��}>Muz�V$���[+��c�e6�=H���ꅾy+3=���>?��H�=M �=��<z� =k�	>d�`>��oC�=�*��r���O�گU�-=�.�>i�B><�=�Z��>�G>*�2����	��=�$M��2����t=��>>n�%��𑾒p�=8�>�gl>��@��zA���R>'p<xuM�h4T���<�t��n4�V���N�=VyW>�d���Q/�m��Q.�8G7=w~����M�ݥ�����=!�V�;�^#�|#�/a����K�;�a�}=/Ǡ�@Jѽ��,�T�\<1�(��]̼Tνa\e�6����a�=��>�����>�fA�c�W>�aE>��=�Y��kC(>$I���]=Q >х<y1��H�ؽ��������� ><q�=L)O=�F�=j�;jҮ>��(=6��=�X�;2�=�^=���/A�=S��<&���3��:���3�0e�=��=��$>�C�c�+�>����=$�@�8a�=CZ�YD����\,��T�@C��}��=?��08�=�cd��z�=�����6<,���Y>�h#�_�<d|���K>�4�<PX�������<�c=�Dx��Ό<V��<U��=�˜=��=QB�=�q��K�׽�l���jK��@V���a��n	���=��->'��=1p>�/C��ѣ��+>A�Y>1��;Q�Y�>u��+�=�u�<�K齙ys��������>3=n�خ��� >?����>���⼕>m����>�@ؼ���=Ko�>Z��=+N�_��=�|�<?W>@�=��P<��*=#&t��e>8��=���T�ȼ��Ƚ��=p�T=Q�\>".I=͆Q����=<�n��~�<���y�=��8�g��=E :��;'>�Qe�"5�.��=<W>dsz��&���<��.��閽3l;q� �?�ٽ@z���>+{�=1>���K=��*�_�&������LԽ�1w��3���[C���<�|8��62�j�%�����Q��r=>��O���-�w�(>3nG=�K>��+���ʐ>Ü[> ����">q�_>V�d�{@뽊��<�>���������)��o7=�d>Z�~>�c>�Z =5ܲ��>՝M>ϢX����;�gh��}>�}>��'�f��>H�B�t3$����<N�=����P ���/6>/����������:�0E�y�#�w�>���<�X>�:>>�i<�^��P>���O�>�4μPT8�C^�>Xh?���j�P�a=��=P5<,c>%><��h��
���=f��=P�װR>#<[��U޼$<��h7ڽ��<�v=�;�{h߻�==�c>b#]>�� �=�`�ܽ���=.);:�t�L����*_*����=���y���\V��� J<���=�J@���_�R��(��
M>5����S���=D�V�<Di<�.>(:����=��)�����N+>_d���o�=�a><.�=��9=�q>�p6>�>7�>���=�=F��!G�k�>K�����
,>�� ��}8�M~���&>6�d>07���g=�բ;��m���0������!��f�5h��=��n� p�=�T����U�=� =�����ET�yO ;��Լ��|U_<���=[�B>�\">-�d���=>�P��Ƶ<]R �K�a���|�6׼m�c���A�ﺑ�+�h��U=�\4=�� >~��?��8�&d�������Z<�n;>�?h=(`�=��л=|�7V�U' �_�=�#r�=�j�=U=�����=���;˧�<A��<����p	<R�<�,<j ��]�=��=��F���>q�>�l<I勽ܠm�WS<.�{�k[�<Q>��=> ?=U���MJ<�"�YiP=f4�=\c[�8ƽh�g��3>dk��!��"N�k3 >��<�=���=,�>@��.T�=>��<�`<Ă�<+�7�=�m�^�<�H��A�;�@�=TwU=��>�k�=�.�A��=����X'����=�f��<���>5M^>�#=�#��W>����p�S=����	�<Q�g��_�=��!�M<�#�D=U�*>s��u�;_AK�(�A=T��<#����i�X9��$��3t���c=6�i�KL<�h�pp��QZx=Qܳ�P��:��=��̽�==)>~T��	)��`��_>���������N>�;����r:>�3��%�˽@o�=ڠ��@'��\�=)�ļ�L >B
q=�qh�|��= f�=�ች�<��K�>3?4����<f�]������)S�r�g�@#<J�G�6:>��V�B1��g<�VC>�h<�޽�'O>/%�j�/����>�=��轷�U=�۽�qX�CgݼCi�V�7A�=4�<��+<4��4�Y>�#=%����_=��=A�=�JԽQB=��<J�m:A�̽i�>�<~��='"1=z��=���&>�T>��.���J=Z6L>>�5>�r�6�����>��a �=�I��B*��jj�K�c=²<�Y�=�9���=V�J<�Om�q�=�<D�>LL>>s�=�7�=�������=,;�ך�3����ڼ�P�=�����=FΝ��jk�}.�>�`\>�*>��Ľlu;>v$=k�X=\_�<�袽u�b=��>Y���7�=�;��k;�;�+��������=�)�_��>�H�e�+=V��<=q�=���=D�M>�ۉ>Hv>��u���P�wS�=gu��pG:���=f���^��94�Ek�u=��>�;c�*>��>���=|�������^�Nv=��=��v>�	�܈D��=Cͻ��)>�i��N�]>"���k��-F���E>;��=��>8~t>�N���Q�<ZA��^R=*Gn�cy�m_�x`>�k)>K���j{�>�8����1�=�~Y>k������	W������'>�$�~�=�L5��<=T�?�\j¼~J޽\�>�R����>p9��]�������c%>9�����	�x��>7ݽc��aP���7+>�P�^:l==^��C�o�C)<J~��i-��n2���0=�����#����<ه(=8�Y�;�=L;��ZO8���E<a���tN	�-���y��Z�+�>_��`�>B�hn=.w�=EF۽��Y>�<��kL�=�Ò�mn�����<�� R>lA<�,��Ij�<WK����,>>�q��<�����#��o���V���*Z���<Kֽ^�q=��#<	�U��3���l���>�A��Ჿ�ȶQ>#����=��=��=W^|>-�:;6į�/�C=|[d�(/����̼�|�>q �<��!�m�/=���=�R���[��>Z��;Fm�.O �~j�Jʤ�?�<�� >U�<8!¼m ��`�1��?�������<� �����&��G@��'�`֝<�7=ow<,�<�7�,���
��;a$>�=��>� �h���=�����z!>���.�]�.
>W�=@<���������8��Z�l>^��=�W���Cs��x���_��g:��&2>v���5Q7=��>ߋ>��>��?�F� �=t�˽�򽛜�=��%=�#=}�&�V	y=5w���&�&�<�������:>�4=��$��6��#�0>��->���Tlg�Ʊc�0�&��>.>�b�<�= �M>脢�����Ҷ=-�ӽ���<����#�=�=5r�=��W=<Y�=�c,��E-=��ᇾd4#�������j�ʯ�/�=Է�=p&���>�a��ڀ��զ=Z������=ԯ�=@ZŽ�[=��a������Z��н�=d������%�x>Z��=C�-��'�;�)>�aH���t=#c��2�<}+<��	>jk�=�?�9���=�k=P�->�o��dP>꯻=Yߕ>M�<�8�f�%=^>�4>��c���ȼ
9�=�>ә���X���)���=E��={��:��="�Y�_���b�k���!�7��=>��=����޽X�*>#���VEj�����o<���v� =V�|���H�
��^Q����j���N�sڇ����=Q� �]��)a��7��T\�=���=�;
>;��������I�=�a��(����i�<��=�)�=�a=�@j�j�=�,>��>j=}>��'<���<��=�X�Lo>��=�� <�����l���@>D�=�Ą�=Ɉ�i`:�B�=bPx=A]j>C�R��H>���=�>`Y���$>��<��:��u>�P�=�|���ᆽ��-��}[�
x���#>X���ġ�oFS>���=�F�Y p��{��	�=�D�>�T����у9�i��<��(�Q[�=����{��<c��=R"<w)��`�<�f>�x����=+��=T*=�����0�X��=@�<w7>7�ٽ>]�<�L��[D>�M2>�j>>,�<@!�=�x�=�==�����=��,>`�f����/=Ȥ��@!�S���S ���:>5�<��=]e=ZV=Q�	=<9s�T�3�K�<[��=�y+=�ɀ��z
��h&>�t���=1��\K>��'�o����5�7kb=˲����߽�'�=��=�R9=(���!漣~��E���n�=��d='����B�<��	>��=D
>KA���{�<��f��^Z����Ž�	>��
�= ��� ����ր��=Z�<%��=���[�~��=Uý���?��=��>ԑ�M,0�m=��t�:F>[l=T��<l�<>�h=xڮ�n$J��W�=��>2�>�]�z�Y>�}�<��>����=L�><�>�{I�@��<IK�P=�=�<��Z�)�=2�ѼIk�=[g���%>����!�=�r�O ֽ�ʃ�T$��%�>Ю�'�Z��-��k�= �ӽ�^Q��,㽃~�<�Q~�a61=�%��vH���|>�y���>�F�����=$,n=�,.�4$7>k��<��ɽ87=F�r=��̼�7m��i2��q��7轄.%>���= �=`1j=+fͽ9!:�*�����;��=c�=N.���v�@>M��>+Û���rx�}�<r�>pZ>噱=@�x��83>{t�=]�=B3'����a=�5~���
������e����:��?= �*��nZ=t����I������=䲋=��z� ǽ��>���;�>mbD��8=��nk����*�1�>��߽�Q�=ˬ{>�)���=Ԏ>���#�4��y(�->�4�<��=e��<F漻#�n=�m�0O뽬�q�R�A��8μ /�=���>,$���	=�.�=�^�#�<h�]�ï����A=����: >��;=�v�=�Qk�����1<�)�=�'=?�b>8��+��<>7�=��<���_?.>�@��^ⅽ+�m=Tk�<�-ӽ<J0�=��;*�q=�=�=)d��}�<�%=��ؼ�j�<�<��R=�-��6T>{�Q��n>�n�=���<�+���:�2���1��Ž��U��.�-w����<ɡ$=���WA=Ԋ�C��m'�=郒���`=�,>���,������üېO��w=Ε�ZA�)�=
-�ݯ=�<�=�9�=�"=8�<����2>�=����N�]Ͳ=Fx=g愽Ţ���ڽ����B��� �=����÷=�M����=``>��=q\	>D���=.�%�>6��/`>���j>�:�����=�禽Y��}\]�����b�$���,�=�c��D4>���=y<T>'ݽӱ���E�=-][�
���1[�4�>s^��_�.W�!�==���n`:>�(1> ��a��l�'<n��;H�=��0��׽Ƿ��P,�=J��\�$��'�;"e=iIO>�w3>��ܼ��������Z��>e8k=�{��o&=��k� �L=�`;M�>
[�=�`�ݛ��U�+��Ь<%��^<ӲJ>e�[�,*X=
�=����V>GH=��>ZL4<|<�<�(�;8�=[���)�1J>�� ��0˽�=���� ��pļ��%��t½�v_=�M�=�]�u�=�,��{W�=�,����T8=6�,=��=6��<נ�0��<��սBJ<n���o�X>�F>_R%�˷`�%ļ�y=�mF>贄=���=ŵ4����=���j-��I�=?���
~�=_(>[==G7��u½/Z�=x|��7>�½=��L<sJX��IȽ�5��i>"X߽U/[=��>���e
>�J�0Kk�m<����1��貽���<�+>]EY>�ZM>an=��=��v�-�=�=[=@���7I�{��=�I:\-��+ӕ<-�pG>� ���>=���(���P����=t+_�^��=����{N<��^=*l��KU�<Bf-�MV�<�i��4?��

��u�<"1	�I!�=�y�<E�<,&>�s��d���
��s�nh=78�����=�ν~N>R������;�>)r��DX�=ڳ=,��=��">{	����;���Kf>�� =ٍK�cv>�� ������; ��;4r >g����5���==SD=�����/��#[���<�R�=~�a;sCQ�R�>�_ٽtn�����҇�`t�.�]�KRl>��1>�ܝ���>@aF�_f�=a=��ԧ�K~�=�.�,�E���!>��4�)�>>*�
��o��>�'��Y���];�K X�4�̽8�=�y�=��S,B>�0�=]*�����>v�=s4c>��<�q>��3>�ҋ<�ݭ�f�ؽ���=B���Q�%��=�n���=�D��:%��ȏ���7<�=��>Nt_>�+�=�P�=�u��o�"2{�U����i�<̟�=��o�:�8g�	>�p����=r�=�ּ���;��=�I�=7����,��;6��0��
�;*��{�J��d����=�1M>�S�����ϋ���Pg�T�=ڪ��F!���XV=۰�=�셽�����3=�q�<3�����n�>>m)���(e���1�-+3>G$�?b�@�̼�#��z�K�t�:>R<K< ��B�GG���=��߼��>�?W��x#=��;27��ý).��6�н��=w��=�����n>H�>2>����w��'�=�O��d�:�>G瀾x<�=7B��̻�=�n���=�,�;������b��.�=�c=�6��t\����A�� >Q���P>�U�<A4>`�����=�`��������`Q��'�'�׆�=�i->z�e==��=���=���cm�j��~uF;n[�<�򅽃�&>��x>�Q0>w�u�##�=^,���<a�a�g,u��>=�.<�i�=�D=�8�<���<�ɽ��o��u]=W�=�fH����<Y�;�s�=�eE�b4=�F>�'"=$/N<!�">��ƽL>�6�Ћt��7>�j�=��=̣��%/��� ���=�6<�>c>���-�8��f����/�g��i�yN+=��>�=���G��/#�(N=ᖾ�w������=��<�X���><��=1�<�$���jӽK���V+�<*r彝kh����=2��=NX�=��"�Z��=���ͷ�=����:������>�K��Z1�M#�Gꇼ���$�=n��=z{6<����	�hb=�=}i��g<�\�:��z=��z���F�"׊>�%�Njl�ף�=!) =��i�">qX�<��սر<�.>h:��������ϼg�>��=お���)����=�9�PA	��f>b9��i[�9�>g\'�@m>�����5H��߽�\>��E�=��'VڽQ�̼IX=�.�=�12=���=I��_=�>/��X�˽A���ۢ>T|���=�W��$2�����	R='[1=�O��2���=Z��<@j!>u3�{:&>�=n���a=V��<нm��~='��=И ���׽"d;���_=�1�=[�@>�9���=�=���!��=�=<�!�I>��L:���4�=t;�v�O�콗�>=�V�;0��>�Ύ=�L�<�<�/�=��<��>ݾk�&M>mx��`��Z��,l�<�M�=�2]=ͩ��}�=4�<����=���9H̼ն;�g���=�	>D׳=C�H<�������9q=\�P�> �=]�V>3�����=-S���=��K=Б��<��D���|>��/>Pွ��=~V���G�=�m�ϸ�<�Q�=�Ƚ�[�����:���=\�a�R�O��=�Y���v��R>됅� >��=]5��Q#���ƽO�j�TM<P��!ճ;d��4X6>�p)�U-=y�>�G=JBc�̧�=����
�=5=�$G�=��i��>d=�O>��=01����=b�=	�>�2^�k�<�=<�H�ԩ��Wf*���d���u��z�l	�=ߠ��� >CXY>4X>��=���z۾b�1��8���ý���=_7Ͻͪ̽�)ʽK҉>�A4�]Ms;K���aVR>6>�ۻ�Ѩ<8'>����<R�>BE��3>��m��=�r���?�8k�>�/>v�]�.Y���3>��#�>��<�m%>k¢��;����3�=�>^>Tc�Z�=D(>3	��w�=�� ���2�OpO�
�=W.5<���<(����wC>L��%��=
 >D.9=E>fpN>H{ѽ<~H=Q�d<vJ*=@�Y��f�����~g<7^�>&�h>��c����,�>���=B�R<�'7=GN>pֽD�ʾ�y�=��\>�t�=1o�>�.��(=,3m=��<&G�=��>��¾grT>14�G=>�]�=�2���X��[4=;�j>�z�7�'>x<����=U>'�3>*<S=�<>�d�=g�D��ډ=�k$�R��>���0����?<P6����l=���IWg���C>�T>�]���<Cm>��h�E�$�E���=�/=q�)m=">n��ᓬ=�W�M��=��A�G#���M���=?�	�y�Լ�y�=U���*��< �&>��=�z�Q¤=uǌ����>�7��>)>å�mR�V/�=',C��x��f�dpk�*�+>���J4˽�p�<F�ûu[��a >��	=��>�R�=���Â��7%��'�=��o���<E�Q�O�>��ɼ��}R�>��=��R�fм=
u>�D���\N=������>�}�%6���C<>dވ�DSu=6����=���=F!���P��U��@>�
>��~>n�{>�#>���&��\'��<��
��Ǆ>��:�]8�d�'=�翼1����1B��?�=��=̵�=XF�>���= IZ>�>�u�4�>8�;>�4h�k8>*W�I��=:Y�)��=?)
���=����]+�:�@>uz��G*����~���q��p�8>�#�<J���Ձ@>v��9��>dF�=�.h>>=��H�&>~�����>;���΍�=*1*��K̼��н��">°���ޅ�1�c�*x��cϣ>�C�rD���[>fk=T"�Q�q>�G>㧕���yX=��G�tB�=Q�y��#R>�嬽�x(�Oh=�7j���a>��=��<��KQ̽�a����������=��½����ƽa�G���v��tb��/g�=���:������>P�=�� �\>����=�PG=o���B�>!Y���,�W�=�m]<��� ��=�w=��	>���
i��,e��~a+�]
�<�[=~��~U������-r;\�iF��t>>u\�>䷛����;8�_����4 >jǀ=�?���8�>S	��Rg�˔b���<�Lt����=�P>{+��2̎=�,�;Q�=�3Ľ㦶=M#�=��>����y}�+Y��Փ��sl�=Cs�=�gR9G�ҽ��/��ɝ�=ŧ=�+����	����i��=���Iر=���:̝���޷��U=I>WI�>sSV>�N>�i:�c��
�u=E�>�VB��e�=(~Z=��v�H�G<J�!>~)�=�}0��!M>,�<Hɺ�=>(7=�Y���=�����e�;)�"3>��)��Zϼ��6>�H�2�Z>yE$�1)=S����W�<e;�=���=��=������� �١�<16�=M@�=Lh��-�8@<���[�=h��>��0��fD=C��U0��]F��-�=k�<�;ȼ�i=��� �B��3>u%���2����;t�>�������=ĒO���=�s��{��f�B���Ʈ��#��.���ͷ�}�=j��>�$�;Z��P#>8�׽�!޽V�=jPi=AQ����=J(��=G�\>6��?�	�y�=1��6M��u3�a�V�?�9>ǁ9>c2��XW/�U����?�O>=�\�=�ݤ=6��i >m啽G8�;�;���cG>N��¹=l��=�A��;>�=P�<�ʑ�I�����4R�<��P���O�v��<�(=��>ƹ�pd���7D���G�B2M�6v>qȠ�%zռQ�}=�^��5�<�YB=t���z��=˽�����J=�����p^=y<4�>4���<�=�,>�<�Ѓ=���=_y޼��s���%��@:�s3>�G����=��'����<�
@�Zr�=�>wp�=b�g�D.½9�=Fu+�Q�㽚�=��o>J�>����P8���X�;�������=�>CNy��۽�>\*�<�j�YV�=�*J���=�%J>�ʽ��=�w�zf�=�� >�8��I>��2�|���j�I=�/�<����
>�!�&Q=����.>�M�%�=��4>�ʹ=��1>o���+�9Y���J�aam>��&3��m�=�}J=�ց=��!>�ȳ�Aø=��7�⫦�3ŻGSD�y���[(��7����5>̩�=�9-� �Ͻ{T$<�`�>���=Ò���5��N�3�I=�4=��=���8#��s����<�t?>����=L�~���ݼ��Ӊ���	�=G<��]�@>�=6;E��0�xV;>@%���)\���=}ā�~����֋=��g>ߎW�7ʹ��9���>ݣ�=y��<�ǵ<��>�jC=0z�=?��Ϊ�=)p�<��*k�=�w'�t5�<����%�"<��_�JQ�%�e�|C[���N��H�<��p=S�ٻ�����9��>T
��1.������� =p��	��-�=7���G=�{���,��=%X�<�g>��I�i������<�FɼGa�<y�B�K�d���=���#>�9�<�OV��[>��=ӫi�?�=���=�����5>DݼpҼ�uؼ�<�'M�5~]����==JO���4<��=#΍<"�*�"�<�����bq>�H��rѼ;V��Q��=2>uN�<�P3��]ܽ�l�� 9<���w�\�H&>(����>���<f
��Dw�;/�dj=U~��������Q@>�:�n�T>P�)=;�������菁=�!���6>�-=��ܼ#�>a��=�^�=� >�hx�l9D=2���k�t�j���a>�-��=��	��'��4�<99D���<�_$�=b0뽽vy=<76����<,��1?�<��d>mN��2>n>)��<_��[�Y�P�G����>¨�=/����^!�=�����_����]3j��E��o>u�=�+=��߼0S=����rkx��<�>���=�j+����s��{��=n�F>n낼��	;�]m<èh�N�`=H-���>ڧ�=LM��'��=	����%��䐽�s����=3O=�=Ap*�
��=�7>�ӿ����=�ҽ��&���
���7�=�|c��и�@��%�c>-f����<�[���,=�T>�?>�Qi�����o|����Q>\Ү�ϼ��E�{��=�z׽S���B%#>3���l=v�=	N.�"�A�Jn<��<L�j>�҃>a��y��=d����>�s"���7�v��,"��GVN�P��<�x=>�{���2>���=p=����=j��=�驽W�;�af���5'>�9u�#�e=q�	��b�<���=)@�<>
�~�=���=��t=�p��5 ��5�=��>7��e�=%c>B�,��r�=�>�d#=�D:����Q�Q�BH�=�����(��a>� �&7<��EZL�»j=��=�e�=�-����V�?�=���8���u���7�=��A=�^νK�>�k�=EH=�(��(!={G��}�=>���-�:=pJ�Jg�<h�4>�h����"����=��=��=?ف�h��9a�<��޽��k��'j>mI	�����%V$=N�����9� ��8�^=t�=��S��a��y���� ν��(=�xE=+}	<�R��G�0q�<U=�=���NpG=8>��ּ�#>Ji�<Ѝ彦Z�����=&��<6�
�� q�<F8>����Uﶽ˓�=�����^�wA>�k���ۻB��<(�ڽ��2�[��=�8g>[��<
��=�ۥ=;t��"7�<�A>ԏ�L�N���=J��<Q�=�:�Rf�=���<�Uܽ󀻼6�4>�i��[�><>B��<�==g��<���<�e�=�(>��\=��=Q5=�3�=s�<�-�D>��\ν]}��m6�<-|���
=��=��!��n�=K�<�7�<EF�<�;��p=�8�=�~;=�,�==�0>���=��넼���->�/2>`H�=�-=0`_��A><^�<���<"x��<�>9i����m�vJ�=skѽ�c<��r���=�l�=��=YN<W�1>�A7>5:>5g >��j>�ޅ<P��=���=�2=�W=��=��=��*�g�`��>4��C���K�*P���{��h���T><�T �=��K�8x������9�=~��=;��<ҡl=��$��2�&ͽ��C�H��<�9=� �>�/=�\μ�> P�����QMM>�#\>F	�=���=#����f�=�`��A �<��4={1�;xǝ��TK=	�=��"=Sc �Bb�=�7<�y=V����=lA�e�=%ˌ�[���->?S���>L�=�v����ia=o!�!�=���a>d��.D>}0�
��哽�)�=(?�=����¼à$>�X�=%0>�N�;h:o���!L`=PtI>x��=��:�,>��|>4D3�"̽��=.����&��,���#�մ>�_�ca&>b�.=����[��=.��=M�'=�
@=�߼�oQ=��Y�j�Ż�"�m��=h����ӽ����G�=S�>�u[<gyڼ�1�=�E<G=¨_�#3>�f=��=��d=��<mм6?�=��!�|������b�(����<,1�ॅ�����m<%Ɠ���!=����yE��ꤻ>��A��=0�=����&�=W�J�|7��1)��7>��Y��\�>���=��9�s\��U��=�e����罴6�^h��L�H+�����n��0�h��~->���=0�=���
�=�#=ja>^#�<�=W���&��_�=�=؏�=.A����=�� ����i�>�l<���<_w� ��=�"��} <{��.A����=k�<��D�1��Aə�Mm�<$�Ƽ��>Ɉ;�G����=�2(�w��ib�>Љ
>��;ν=5쮽�W������A[>de���s��T��A�<��=��=MѽB�@��h'��	I>�y�<��8�Z�̿��ͅy=���=���c��|L]=��}���.���M=����Bq<�l= �'>�Ⱦ�꥟�)$�<�0=4X���,��_Խ��*�_�����=���<-��= e���^�=�qH=�:�<g�	�y� ��t�<��e=x�B=��"<]]=���=����<��=%7f=E.�=�ν�9-�ތ�<�	p=��"�� �c��=�W��]�2ެ���< p�=WNf>=���M�����=Bƶ=]�˽r�<rK>�I���Y[u=���^4�g'�=t�:>� %>�NU����=
�˽^ >(��]�G>Ǭ�}E>���=��?>���=;A	��7�<�3>d,�wd�����
fx;,9[>�����f=���B>D�>��F=�<�=@�S���ļ��P=m�=��C>��&�T�������Q��$��m`�6Yo>���Xy/�%=M�<�-��ٞ5=;i���=^"=b?O��==�J���==;�@��붽�D����.��Hټ֋ʼ�k=�;�:�nw>l�Zo�=������<e��9[ֽP�;���9��C��a��<��$�^��~&����<����T<w��m�5������ؽ3�ٽ�{B<� Z>H⌽�ٽ �˼/E0=��G�jS�<𣠼��s�g�=�'�=��<�6�;�9J��<4�6�b�M>�|��3��;{���޴S�p�>�qнA&��a,�y�<xQ�<k�=�j���=N��(0Ὢv:�V�=&��=QR�<4��<��y=��=W\c���==�u��OD-�Q�X��^!�c�ؼZ�=B��=X�*>}����K]=-"0>J��=�\(=��g�(]�=Oi=N��+C�No=X�=ee�!�V���=^}�=nZ���</)ܽ�����*�̚0=��=v#����Y�2@i��.<��=v;>�=�%�H��;��`>I�=��U=��e<;�D=v�r�������<W�<��4>
�v���;�������<S�N=h2�<[=���=ؓ;$}�=G�����>��G���>��=����E�u����;p�=���=�Q�=�����m=��>!c�=ќ�<@��r��=r� =NV���4�<ط�=<���艼��H����f��ŧ=t8�h�c=��ٽKʆ��L=��<����H��=�Y׽S�ؽ��H=�h��v>��>�)����<��>=W����=��=iJ��;><�Ļ�=���>��/=p�3>3&�=?
���㽎�2<?�轪Z�=��<���a=�Dֽ�*=�0m�r6>������>����[�~���b;3�,=kJ�<օ�=%�8���*�v1G���>G��;���� Ͻ.=�=�_N=u	�=^.W;��.>^�p�Q�>��꽪�5��1⽨����Ѽ���|�;�����B�=A�D����<������X���>v�=Ȅ���C�M=F��a��.uL<��M�rH�=��>��5=���=���=�z�=��=�x�=׈-����h�D��}�&=�x�٩��EE`=�G"�b=>�	4�.�)�7>��fm �!�\=�$�=��Ϯ�=�tX���*>�O;K��=�A$���<�ߧ��͟�%ᚼ�k�����;2�1Y�=�:vD�=�V=�½�[��K�<�z�=Ұ�W��=�D�����=���=���;&G]>Hp�q��� =	�O=���=��%={��=
���L����LG=�$h�0U����.���{��>u'=\��4%�=�㛼eo?�ܜr�*��=]"�;�'=Ǧ�=w�	�>�=���ͯ�=���9��	��%�=��X>�p=���&>�'����=��=}��<1���4<�G�����^��]�<�!'�|���`��Cp����H>8����<>�iؼ_��=�=1��=��?<==��'?R�������G�=�<�Y����.�tW�5x�=7�> �F��8f=۴����0�=j=:r�=�&=�m=c���˼�
���t����=x�>;��=Ub� ���a*=�l}=�״=�֠�K�,=�q:�"�3�̽���=&�n>����T$;>ʔ���0��q���I>��<>^D>	:��껽�]��W��=cGн>��=��/>��F=!H�W���d�/�)c�=$>B�;=ىa>���=>���G����}�do=��=�7������=mK��~;<M�t�}H�=�7=�>K<t��=;�߽Āʽcz���o>�`��Cf=��b=}�=
�˻O�)����=�.���$>#V6<u5�=�?��1��m�=+T=t�<��齶e�=��>�Z�z�Խϊ�2&ƽ�t=<� =�>�轢B��g�&=�ƺ���j=3�v<�(q=!�e���=?�������*>|Ɋ��#�V���[-�!�s>�C}<���=��F;i1�=��l�Mq�=w=5�8��H>mB(�Q��=R�<�W�� �H�o��r=�->�)>�%����;c����=v"f=)�;� �Խd�2>ϻ��'<����_����{=�O%������JG<#���[�V�p<��Q�.Va><=�58�����	�:�Ӊ����_�9=a��\��=��=�l<��@=Ax>�����1�D	#��Y�=�1ڽ����������J'��[=�Q�=�w>,]="^|��'��F6<Ie->B��u>#v�=U8��@/���n>릯=#�����>���ߛZ>���H>��1�ip�/�ݽ�/��N!�cI�_W㽪@B<U�&���/>�I�=	�>��;xJ,���:>��=��=�>->M4�'t!�
�>½�<�)Q��m8���>N�p��>ӕ@����_���������=��=M<�:SQ>�>���=*c�۱�<���m�=�<��B�=����:j=|����	�����b5�~)u<�N>�=���U��;W��;�� >|&F=��ռ�=��:�s>d >�$��w���TP��m������}����;� �>XPF>"8E>�! �u:�=~��;��J>��T�D�M>Ntb=�JU>�\�d�={�ٺD+/>�m>>�>�&��uȩ=r�����=s$f=���iJ=�r<ؼ���=�=�F>�>��q�'>�z���Se<o^�>�D=�u�=`'�f� ���ӽ<P���V��ݨ�==�g<�G=�,�<DA�c�=����u��]��ʐ���@>���ä/��E�=�'��Iv�<��L>�GP�玹��65�?[>u%�%��e��]�>J��N����<>�_�=Y���l$>W�'>.l=
O^�ȣR��Z��
ɽ)�����h�/Uս���;�4F=x�H��m�=�Ɇ<�8�_c�<���
t�m2A=|�>Ӏ>��[>�����9<�Ԩ����~�ɽv.�=�p,�����}Z��8]�)ɗ����=�����`,>�{��b춼�1U��?T>{,,�md�;�wC=S�P��)������=L.�>���=�<#;%�4=6��=�Z��"���x�=OՉ��=ҭ�t��=ޚ��,�k���=�,v=�,�=���=��-=�N}=尵�8�\��MA�W^>�H�ۄ潼�����=�}˽�f�m_M��t�=�=�t#<�����=��?�t�M�~���<��={�S>x���������=AkټuÖ=�#p��
��^7,��I�d!=!�����ɼ�$F��q���
��u�<���F�;LE;>w7ϼ�%�8=��?;�e�J<"�=���ܽ��=x� =8�W�:aA>�l<O|$����� ���1%=��A�;39>��qz�bv3>��G��?�=��W��#>'��{�'>�F-=���=|���<&��<,�(�� T����<�L��T�U=��W��?|=�)F�F��=廜�>	�
>%���A�=�V�=�����[ޡ�Y�8=D�Ǽ&8�=q�J����;�^ۼ����
U׻��{=�Y�AD�=��Z=�M�6�J:��ƽ4<�=f�)=�!*>�l`=Kɽ�d=�$>ro⽃�>��>�� �y�Z��Ò<�[/����=���=�n��,��m��=�����������E>d��4�6=�=��)=�C�/�߻R���-H>���=��h�=�6ʻ
e���ta=���=4J�ط�����}@<T�= ��=2��>'V�{/<V�=r�~�1���h���=%��S[O=����8mr=c>>Ω�<�=�=c>�n>� �<s1<E.n�a߼�~>4�M�$��=��=���.�H>�ť�
�\>��I )=3��5x�=��ü�>���l�0���<��=S�<x����/�<A=�>&������P�{>����_�=Id�����=C��5�Wb>Ud�=q������%>M ���6��x>�+ѽ�$l=�f+�SlD=���>�����x�������ѣ��x<���=��
>�UI=��<=P��
>iد�B ���=���<�K�F���Ԓ��ʃ<�)#�-W�=�����=Pm>&�)>�)k�o�����$��Kƽsda>�4=X�ݽ)	 =�-�=l�}>U�$=�}�={m=L��6�=־���@,u�=�׽�V>�d<_z�<h/7�/͋=t6=�]=�?E:mp@�p�q���${�`���c�� F�5e�=�������=�<� ��� ��h����(<�+=�K�<��<<#>��g��fټ�M&�h�B���`�X\����#=G�4�2=��=�N�mܽ���=+!�=v�95!>�o=�S9�ٷ$���N>�J`>�{�V�= �]��$=,��<��2f��Hd��<Ͷ=г��i��l�P>SO����= M�=��=&#`=!>�QP<7�?�����Z�_�oa�I�<9H<�+&&<�Ri=w-;>X�ؽ�0=
�'>vY�<t�<���=c��=�<�/�5�==>�a>㓭�RO�E�*�w?B=�t{�t�=��=ǁc>����B��X9[�?m�=��=R#��2��z��<D�.>Y�ǂ�	�;�x���@���o�=����q���,=½ս�=;�+�x�I>o�w<췽a'ཱི�G�]��<A	�b}�=f��<���>���Z=��=����<�(νy�ԼO㹼�<�=K�-���=�7���8q�9�>$��\
���b�:mԽPQ�=i��<����c�#>Hk=�俽AAȽ���<��S �TQ��2�:L`�=lW�<L@>B@��.�;�C=�Ƣ�}�= uȼ��'��Z>�<">��*>peK=��>Ùx��=3�I�sUZ;���=&����M �YG\��m(�Rώ���J�|�>��_=	�H�]��=��K>�茼o��=�.��i=�>N��&�b3���>�)���1�=Q>�=#E�-=�(���C=��/<�[���0��Q�=���A���4�@>�x>R'�=Ak��ɽ�3����;s4��<�=_�����]��
����=f�s>8'���<ֈ<���=yM�8�����l= nE�H��{1>�y�>1p��k�>I\Q����=u�����=���',��[���
ʽT�>Ƒ����D>��=�n��#��! ����=S��=�_7>#˽�>]�6>V�9�J���m�>X+{���&�#����(q��-�=8�����=�l�+�K��Z���z^=s�>�5'��3�Ռ;&bн����(U��;#=�%�$���z<8->�<ܽ�K'>�S:�/>mi��,݉=XD���ួYx�={�>0l�;��d��u�	>��R��v��3�2>:��>�<��>���<���6y���ĽS"M=d�s=��;|r>������z�<�C�=m�R>�VV�-�>�G=�����v>�s��|4�e��_��=��;n1��f>�Φ�K�>���=^��=�����=�z �۶�_����<�b��=ɮ�=
�G��ȵ��6���^K��g�<�� �>��=5��8މ;t�=ʺ�<�h��턣�AS==�н�� =�ӽ��=󔅽�9]<9y�>��>%g�W7=�>q>=�f->���<�g׼�i��id=�^)�5w>$���[c=����X�4L�<O�=�_>��1>x��>�g����=���=HǍ=�.,����=��������D>�s	>wq��B%���e�#���>^�$>�����W�=J�=N��=I;�<��<�x}>�y��j���{�;�.*>���ª~=�[ֽ"o���'�<����Z=]��l���Y���	>�� >�(>r.��|�6a��.�1��<[�o�E>t��;?��[���b�=�7[��;t>.S���>�ؽ�d<J�9��kX���1���@=)I>Jý9nR=t���}ڇ=
Z�	�?>�!����=�m<��/��.@~�{3>R���D]��"�C�U=o�E���<y�^>�ʽ�su=���>3�
������g=Z򒽧~�C�l>��=Y��<u&9�8���!�Ú�=���<�w�<���Y?='�>=`���[|�=���F<VH>> w=��>Q�ȽVR=��=�!=�?>��)=@���>0��=��R>�7�=���<]�=b�1=n瑽����v%N=���=�f�</�_�@� ������>Lʽ30�<�Ms<	hԽ��=����(�����p�)I�=]�ս�d�=�üHZ�<�c;��ϕ<�������\�O��t߽����!�=� ������yмI�	>,�>\Ԕ�!�P=	M�"s"=�x��`>"1�=OXg�$��=�;��=b5;�LGٽ������=J����b����D���漀7��*.�<�V�=[[�=c����|x=�������=-��0�=D�=e�9����� �>�T��<�|���;��?���]>P�<�m>�q�:�W�7����{�<��r=�=g�5>a�a=9�=�㺔��=V#�=�<Pw>�`	>xno���p<�p��~O=Z�:�6Y�=`�)���ϽC��<��'=��%��)z=tʴ=ih���)H����%dx=�X#�_��=
T��|��A�=�u�@���(�Ϡv�;��=bp+=��>�pp=�9�������<Ȅ�w=H�r>,�����ʻ��l1w=�*�>=뼹��=.˥��� <�e�=����e>ž��"��F߽{%����.�hM"�b|Y��z�%ν,y�;R��=4wӽ�8/>�߱��_���ʲ=��B��=�G�=��v�8�&<2N�=���;��=�8u�;�$�)���y5�VF��V�<��9����k��T�>�`ܽ��=�8���o;=����}\���ؽUY��S6<ʴ���̙=�ν�%����1w=��߽�*">˯I=����{�����;G;!��=Yō�+E�=�սm4>R'�=������ԣ}=b�<-�%�e���8F���ȼ�>o=�K>���f&��&m��������C�h/Z�g��˿��'S�;c0<7�I�;R�f�=W`�=gU�=�<��O�IG�=�ʖ=<ur=o�i��<C����A�́4=��νdڟ=�U�<Qi:�:��=O_=)"ƽ�wU�^�QDܽ?W�uC=#�=�Q%>7�������P��<Z$&��'��z�ɼ�O2:w�V=�e��a�<b\��n�]=Ue�=�9�m�<�Y(>��J=�z�=�괽� >�^A���Ž�U�����c?������|��в=~ϭ=��������匽�W+�C�����*=�Z����d�W팽����i�~=�N��	=ȧ�@�ӽ=+��
��z1�5��=+��=�c�<y�=����ʇ9��<�ۢ=�9���>>�9��&�9>���<�٦��1��C����W�,�<P��=�k��<V�|�q�=�g>XT5�.��=Eu��'���ዼk�>�8(>pt�1��=K$潲e����Ž�>М˽��|;��>��=9�B��<>�Q����=g���S�=WF���>R�<�=�p���"ǽ� >���<�-.=�T5��	>����Y�>�νH��>���=@dq<�m���Ƹ�z����2��=�=��/�y��5���;��=�0��%\�=����2,J=��'<C:��]o:=���=��=�؇����=��Q�9���+I�=
䂽�8����<����佋�n=����L�<���ì�<lT�?�^=+�f=�=7Q��-�:�����%�@o=�.�.k�='��=�� =��޽��+=�r�<��=˼7;Z�=�-�N�><�y����M����ٽڋ���9>��E�ʱ=R�>��J���=l����"(��aغ�����Q��>� ��\r=�2(�<͆?=��=��>>�D�%>��>�����A�=�o˽.!�=b��<��]=�ٽ��r�[<�/#>��'=|�G=(��=k�<sڶ=�>�&����U=i���w�����=�z����/����=%�;<!�"�>�ou=7Ak�$(��d�ӽ�R�>� �>q�
������G���Q�={#?g�Y����.�9�>4[��m���0'�������>J�>g��>1b> �%>�M>�i>s�9�_�=�S��I�3�<F��M�N/8=�k'�'��>{=̧M>�b�� ����i��|>�z >$xG�꾺��֭�,��=S"g=I��;�7��h0������)�i�C<��ʾ*$��=�<S>~�m�Y��>��˽�0>>�Й>��=�G=:	#�Β�>�ҵ>��>6~�>j>c�ý�n���>�6	��,��̗�އ>d�C�����h�� .�]�(� �{?�¯>wn<��Y>�[����
=ꞈ�g㦼_�'>Ө�>	uZ��}=yK+=v�U�ť��5�־?m�>>sS�>�p��ȾCNi��>�vm�w�=��o��Rv>L�>H��f�p�G�?�����*>��=�=� ��#��ͣ>C?$�n?�;ڱ*>��8�dĞ�:Jq�����i�>��t>�(#?F�=��s�GǸ>&��=�yü�Cս��<��k�3 A>��M�5&��j__���B��2E>ߌ�>�
?0��>C�>�Z�p&���<b����������ξ.���}s�XqV?O���m�<��b-�=�,^�����H=��?B����>��Ⱦ�@�> ����&�������m��j�>�"���|=g���!�=����k㱽��l=9v=�'Ǿ���#�>�b��>z=�K�>k8>�۽��)=��`�Lf���oԾ����(�>�*ξXU���x3>�?��2��G޾b��>���>y#�>��=�1�k>��վUD�>?�>��漦�d=�᰾`׊��	}��ȼ��w>;y�>b����=��=�{�>ߢѾ?�>���0��>���5余��<�>�O����0Q�<dԾ��`���>eI��}�>RI6�' �-M�����<æ$>�^o=�'?��ľmZ��}�=�s�>4�ٽ"�S=s[�O3>�	���?���c%��	3��x�6�I��~��ׅ>?�?V�н#ƅ����>�>ihL>>�H>��˽q~>�l�>L�`>L��>�P���*>�J��ʵ��ca>Up���-}�Ƽ��V�w�7���̾N?�+����I�>פ$<��>g�d���>�>��&>I��>op�>~��=��S����>*����jF�Q��>gF?�������>_��>� ��k�>';�>�K.�����Ֆ�g�>E7��E�oD0�N��>V>�=t�aw�>��;>��?��zQ�!\N=@=B���?ԣ�G�>R���l���!?�&�fUh=������>�ா
�¾�����_�>��.�L
�=�ϖ��%?7W���*-?"�=�u��Z#R��Y>�^��c�">��z�3�>4�4?䦁���ۼ��T#���u�<cz��ξ�k�=��P>�l�����<�_�>�>r�=���`�3�+>f�,>+Ɏ>�&f��]�>ܟ? ��<>�̾��K�Zޅ>^�">?8N�<�?�対aY�>f"��`���<��LϾ��O��a'��H�>I)��=1gȼ�ר�^���LȾ�>i�*>^�1� �׽��ū�>��=�T���ɽ�!�t��A���1����>�6>���=W�����>;��췱=}�?C�ǾmA���*�=�㽁x�=����
���\=1>�P�>4 ��Z�<��3_��0���N�{r�>�;�>%O�>�z?`�<=Ͳn�ݻ)>���=�k�>"|>���A�=vԋ>�y8�`��G�	?��>V�?H�F���>�Do<�!�=IRξ*�R<��>}׊>����4�?ಏ=��A>[ �>���>� �_�H>�´>�7c��y�>K�=��g���
����쾷�3=�p(�Y>!ǀ>����\�!?=u=�������n�<���n��=�=�%y��8��(��>Y��>�v��9湻��ٵ�ǰ=�_$���=�삺��=t��:����=
�l=G��>�ǻO�==�=�Ok=�ۂ=� ��$>�J���p���r>��<�B��h3>��V=���q�<�9Խ=Z˽a!����,&;����>��=�|_��U�z�={���z��O�<���;�n�K��i%��Fk�=�Vͼd�/=_��;�9�<LR��s��%�!�|�ؽ�7��=��
���&=�I�=�>j|6>�0H=.AQ�T�-h����F=y[�<T�b���<�G�������3>4a�=;!�:pk��>#�h���=N�ӽ
�=;��#��Ǽ��>���=������6�i]	�+5;�1�=���=�!k=^�?���2�M>�&Y� ��E�=<�<�|�=ȕK�Q�=�A�=YHV�D�=�	>���=��^>��{=~D�j�<����u>��'=�O\<��>s/�=&VU>&ȩ=���J)�=ǿE>�=>=�A�����Jb8=�#>S][�0dӼ���P�>�X=�.���I�=�G����<����;>+R��Rg���=)�R="�O�ȓ�Jr=�jF�COb��������<�=�c�=H��n��
�6ܽ<��*M�=���=�F����=�0F=��=��8�,%���6�����=j�>Ey=�ڱ�H�c8F5�����1B>_>½���=Uw�=�>=z ��ݒ=�������xzk<��ټ�u�(����a<{{�=�l>�^i��cE<��x>���u�= ;�=2V�<�7�<>05�]����>��=Q5=�7g�t����=� 0�`��@�|��"�;���=�8��`�=~Z���Mx=���k%�=��=<c?�)�=���'�Lx=Ɋ�=�Ñ�Km��������=�h��e\�=+�����=�� ==/��=7��a콲1���	����1t>��S��3�=֞G�f���c��jχ����r9p�k���LԽ��Ľ��<=���=g�̻,�&=��
�D��$��=o:�=�(�:RW5�'��n�?�S���d�N>�5��U�;=O8(��Wռ:��=,�J�&h>�?d=ϸ<4���
'>Eӭ<�mȽ�!>��[=y �=��E=����#����TeT��ɖ��/���LO<"M*�k=��<��>��b(N>���+��=S��7c�;���� �HWܽ�$w������&����=�=T�g<��ǽ;=�=�+H�Z��<���=WIս��3(��F�S�ѽ��0=��=Ϟf��<@��!�����<�9��u"����<:5a=�7��s��A[6�H-��l��A�����d�e��=0=\��^X�=2�i�,��E�:�ܽ媁=߄=7�����G�����D��:`H>N��=q�=�>	�����=���;�#*>s�=�R:��.����g�6���W���>K�ƼN3�=/W!>O�	�h4]=��=S6%�h�=B�h<�=!R�����~�=.�>]+��*�H8���<yŽ�v>���<��=��+>jMa>���#�<D������=��=MO>���=M��=ET�=�����>�R����� >n�=�����=�
;�pi�0A>S5>�T,>(��=� =�[:���=��/��
>3��=^ݒ��F���P?�c�P��<6�=��=�\ =�P�<��=�u�/!�}̼Az�=O�޽&�=XW��fX;�3�#=�\����=}Y�=1�=��ܽ�mp=��d=M�e>rҽ��<�}��6>X�=$�9�n
�=$h���/���i0����=[	@<9˞��?�<�:۽�=�+�k%�Sr=��'>Z���#>.ü�p�=,>~S�x��ff�=6��0�e�"�=�6��q�L�C�<�ڽI�S��=-4�=��z>�!)=�X_�Q<K���Ѓ���������<�yH<�J��)lｲ	�;O���G_�=��ݽa|λTL���Y�=z{#�un2=���f2>�A�u�;�|�ͽo���n�D6C=ա=���=`ƽ�Ը=�̖=�J=��m��R�=C�J=����n;=^�O=�C:	��=6�.��<�6<萈�f��<F�<ĩ��;�+��[Y)=l=��<��ҽ� ���V�K���=6�=����dx=�^�=ѼO� =��k>�x�x��<�Z�����=d����꽂�=�%���νO���tv�=�<!ս��j=_|s<US&�U��=�+�;/L�=���=����Z66=z.(>��O;㿬�D��=�rK=`Η��ײ��=�4U��nХ��:��X�ŻW�=�)9��8��j矽�*h�Nq5��z =s���k�=��鼖O�=z,�=��x;�	$��.=�ٻ=!�K�A*<��=O5 >�%=轚;�ȼ��B>Ϩ�=Vw=|Gt���C����<7+�<���<�f[�@+�:�=|�I�A|�=�l���k��O�)����C=S��1 =6�M���<��r���|>�&=��=�R>̹��!�>�:������9���c���<G��<B��A��<��>!�/=��@����b�>��%>*�s<��1��97=�s$>��� v���1����;��w=�$ٽE���z�="^v���>li~���j>h��P�=~S=S�3]�x�=�
�=��=����f޽F�>���W�=�砼�O�V�>�e���Q�=�ü��<D.N<����O=��%>��	>�`_�p=kUɼ4�R=>{f|=���l��l��������g�S<��>�e��~;�!�;>��`����=����;>�P��ͬ=����t�<�Gl���";�v%<b���#;����X=�=P������75�YD��٫�l0 =t�E���*� "�=� ���Ѽ�&���	�������~��=rL��TH�IH����=N�a{�=�Xo=��ͽ��>�e\�]P>Q̽�����=>�V5���T���<R޶��X������9�=�ռ���d����<���Q=�:��=�R�֌= ��=���=�;q�{+�>1�=|�V;7�2>Ĕ=��<Յ`=�d���G�_?��� 7�vi>>�̀=��8=���<?����<�����T�=�fy=d�<�л����ã�<�P�$� =.y'��;S��ge^��>g�K
k=���<�����B=(��h�
���d<s�=����;��=�C�<ݹ=�2`=����D.����3���F�A>*VȽ�7�=�!~�9)��y>��>+7=�>ՠ1��M#��<�+���� t���.>ۯ,����=@��+��=P�缷W��pE��3�E���B=I)j;�:1=�d-��%۽��+=^��=&V<��b��iT=����i>��<'g=��S>:�>�ų=h��<�VC��fO�lx4��0���#>L�3>�`����=���<�6½��F=��U�q����I=�r�<[��==���v��5 ����q=;�;����<X�
;E�>ߚ�<X͊���z=���<8%�Q	�<4���,+���&>)1<�k�=6�2��J�s��<Q<�Ҩ>�d�AmZ�+�$����=|�[=#�=���>��= D�=�A><�L:�x(=R�=CX���"s���Qd�<&5ѽ~"@��#\=#�����=��>��>p�~;T_�=�N5�/`a�;B��S.>��F��o���(*>����2�=��^=�A����i�&H>�d�ͦ>P=� L=�gh�&��=07��L^�N(> �����=lq�=�T����=9���>ݼ�ˢ=$�4����8����;0�ѽSŚ<�2��P>�^��Q��=��*��D�\y��{p���[;> ��>���	��=
g�)���#2�,��,�==)Q�=N�V��=-�=�3ƼU��=���=�[<<�R�-��<W��=�=�=E}0���A=:��;�;%�I('�/y>�+���-��8 ��@�<	�=Jk->��D>�'<��ֽ���=��<@�$��P1�޵�=��=:.O�h�>i��<^�_=�{�_�<�=؇+�m�=5��=QȆ=۫��pz=)'e��#�et}��Q^��s>ѕ��F�<3�Q�~�L>)�ּB�;,��n6�r.>=Kx����<�3=�-E>�T����>1��"j��$��	�%���>@.<�E�[�)q<��<�����>�=��@>-�m�|s�<��ż?��ڽM��=t�->�<�>Y�L���T>���=��-;7Ã�����S���=��=�� ��V���w>����/���)>�W�< �=�4�<0��+fz=l�><%���e!���.=�O$=G]'>s���a=wT2�La��M>�p��P>�&>�s3�d���Te��l�#/>+�+=KKֽN�=�= >L���=cl<��-��8<��>#��;|����r��rrl��<��=θ&��[��>fi����=fʡ=D��</= �?<.�Z���>��o���h>�ҽq�$=�E�=E;�f���D�'��=k��=|Ş>Ҩ�0��><�C>f]������c�l�%=��?=��=����B��q���A=�lQ�PT[>B��g��<�1����S>b��<$�7>9{=g��=���Dp=ݺB=?1��r3�
p=���=3-�N�=J��<yPA=f���W���� [[<�U��3>178<�@��C��=�N�>S.�<H�����,�M�=k$>$>g�~��j���3>,[��~X�=�Y\>Z�>�ѽ���w�>>��m���;�'�=�>UVi=�I���'4>_m>wm[=���<ޓ�;���d��=���~EM<i켼&�����;����g �TUh�a��=)���5��=.�3���[�ν��m���Խ ��=���A@>`=��f�C/}��-ɽ�Dl>d8#���=o��=�JG:aS->A�>���<a�=	>�n��Sn>���TW�׿�[^�=֚������8Ƚ�Ku=b�=��Ľ���>� �����<I��Wٽ\U�=b$�>A��=�ū��E~=~��>���=i=�|�>r[��MR=�T��kES��v�o�>�.��U�
>hJ�?�v�U2���a���U>i�6>˼��=�s;#����>\S}>��߼ H�=�\=������V=�.^>|y���>;-���m=c�T,��'o>�L�=�=�	���߽�ǖ�1�սx���O��>qǺ𡕼;B�=x1L�`�y=��=ܻ彎0d>�U3>��޼SE>�M<2�����8�%>�f>�{���Y=&�ǼA��:��n>3�(�!��'�<�䆽N���A����磽h�.�ʆH=B�>/����1�G⏽V���{�LK��P�R�h����=���U>Z���R�+�=��
�n���x��=�����L<�'o<w=P����;�	<')�0��d�<� ͹�N���>)�Q��G>fPl>��!����͍=`<��I=ҩ�}!>����˰=�O<�8,>��=<�Ua���ƽ�- �"ݥ��A.=o��< �=֔*�B�
����=Y��='�q>��=$�-��*�b\>�$�>�2���_=(염Z>����>I��=��׽-��ۉ=��)�S�����5>S=&�#X >9v�F�=�Z���å=J1�P�<���q>�p����=dT���ۄ�V���p���7q~��>s�`�{X���Ľ��[<;�>�T>i�<�of��� �!1=�����c�<-Ì=�R�\:�=_
��iF���h�wG�'V�~��|�<>?)�>��	�z�D>ђ�;#�8>�,���p�>��Ƕ���>��ݽ�a=dѤ��9>�ս�B��Y�'���8<�g���R�=�m�=�o�=5fR=vշ=����m���<���:�����5>���<lԞ��N>Bp��D�Cq�=�쫽�)�MW�*m>�"��崼ڬ��|"��멽:�"��oY���
>g�#�=��B2&<�Y��>�=����!�I>mW��>�4>إ�<�q>�U<�Ƚ.�����=�M�=�QR��콥�U=]�ʽ{悔��=�Y��*�&���!����=o�Ѽᗀ< y��c̽���=+��=)���ӽr9ǽ�D�<q�r=�潘�<��V=}b̼_�}��Ž�_��z��=� �=�l��Z\�K����;>��J��b���N>N�F�K~7���=�W�wuM>�G���=Ѕ3�v�>>��=��o=/���r��
����2>��=i�>�a@>w[���\ ��U��O���+>�b�=݆�<��ּ���<�w1��6h=-֑=!W�=#\̽�	7� ��z=��=P<����e�O�<v��=3�t=\〽}y6�h#;��<C��g܃=ݿ�=��%=@C���B,>�Dg=�N�=��Ġ=��=��/�2�ѽ�z꽜��=ِ���S=p�Ph,>bF�=��<CH�����+��QD>c��JH�=Y���<什���<n%�=�F�=��)=����>><�<<�3;H�w��һ��n��vӽ���j�=�����'(>�V�!;w>�sB>�13��$��d>B�:��=��b���E>�g��.����Q�����=�,>r�?>�>]9:�&J�=�X+=��$���ѼN�y���<�t�����=m�� ԗ<[a=��>��:J0��.=d�'=��V=����'�<�۽/S���O>�Z��%GQ������=��=7��>K�b���#>ͣL�b  >Fo�0�=�2��_3���W=�W3��]>g�X�?Ĳ��X?=���5��*q�<����K�>Y����>y+�<2A�=��ƽ�JW��bk��t��&8|��(��k��;s�p��N�/�E��%/����;�X<�2�R>q�=쓺��:	Z�<���=�Ň>�U����=�n<�˄�:��=�F��Q��=�o�����=����Dט��;ý�绋�
>�f�[c�=>��=�>CD�=��<뉗=�b*>���V�>��<	���բD>)��<����C'���潍������m��=c�ӽU� �����=ĕj������+=�o�=�������� >k��s	�=]<=h+��˵нjjȽ�;:�(�R>�K�=�&����������o[=���[��+!<:
T�=n�e<�w>��ɽ���Y�=���_-�w�?=({��i�*���=$�e>�D�=�_�����=�J>�\��=��<��Z =���=�j��{�*�g��>8T�<'8�hp�;ݼ�s�"��o2>&��;�'>�y>�2�=�C.=�,���z��&FC>��,=B�9=�H�/>a̽
![> �=9�=1�D=��;�`X��_5�|�|��|b>��j=�Ml�#�=��R>��<wy�=�T>��=�Y7=A��{%<�3A>���=6̸�9p�<�P{=�f�=Oj�:D>�B<��	>�o�z�=��$�K������ս��_>�Ӥ���=񩯽�$�~���%��=v�<�u���������l��;����3>�T<D(�"�=}d漒k�=wq�=��=7`�=�)=A�`=���=��*��=6^J��
m�T���he>�\=����t�<� =�l⼡�Q�e'=�9_���	���b='�Խ1�3>��R=��V=��=&�E�J:��倫��ET�������=���=M1�=��m�ғs>�c��D��=�X�m������=��m>Tȱ=�_%>岸����<)Ǩ=F�����r�x�Ǽ��)=�r��!�⥯�]�v>ぽ��=A�n=�7>W�=�1���m�:����н�ɽs���D!�����=�y�<�L�1dҽ �<φ�4��=-���b>�|��=i8=��=�� =k�8�����i<��H;���=�ǽ`i �Jpd��Ј=
����C����<>�����Խ��^>e(�<�<��'���D�ہ>vzټ���sB]>�Ҩ���%>��ݼ��⯽ndC�ay�;�IZ=��=�M޼�[�9��5	���g�Z�<~�/�~����Le�6s�=��=`��=���DE=�+>F��=8�!�M�2�B�#>G�O=���=�Ŀ�Y�(�_t9<�콜��w�(��]^��]�=;��"����i>��?=0_�=��0���.=�{�T=T���=�+p�k,��4=�^�=����=z>>�����~�9�th	�P�.�8j��kk�(>�A�=j*v��|�t]�=z̛=�9)���U<E.м���9�{�H��=�ϻ�	>���^�=Y�>D�>�ܥ=�h>V�>� �=�?ý�~z����ދ>�6��9<n��=׏D����=��1=�j�D���#���I=I�Ž� >nz��}�=9�=hSz��M�=iB�<��<)N��1���r>�s̼��/��q���d�_xC>�"����^���=W�C�=]!G=�9��|��:<v�I<��nb�*�F�	�>^����'>��=�w�=�����=�=n� �x��$=
�x)Ƽ�e��c�fW�<P� =8���vF]�[�ҽ���=��ڽW�ν��>%��K�;��&=����������Z%=*�=�Ⱥ�g{I=�#�=Y��<rx[>f��=�識�-��;��=0N<3~!����=�!>W���p=�=�1>��=>�������>�*���&��J\=��e�f�3�|�>԰����;.x��'A�4g��ސ;��"	>jZ>V7�<��!�=j->�9Z���C��kN:��4<���=L���活�����k�tO<��~�=�<H����==�/=�;�=,�ǽ�w�=�'!;@�=4�=,��<Ҋw=�g���=_��=��=��Zo��3���-�|Ș���<��=�=&����=>�u���=,�;��>Xd�=`�>=*Y��I��=md>m	=b)����#=1(�����,��9�>�sB�2?n�����%�=�h�>��ż�_��ټ�T�=1�&���Ƚ�5	>�\)>�N�<�a�<���C=��W�Ъ<8�N��������̽���<�-н��x��>�=+>h�h��<��r�~;=�F>���=�����h齖�н{C��v��u��*�G�*�=���=������E>��n��=�/N�Vs>ꋎ<�C$�rR���?���R�tR�=
��=�/>LC�ϐ/=*�½�ȭ�o���.��<��J>U�f�A������=��<r�'<*��=)��<��޸;=	+��I87=�=�"�=ZN�tL��g�=���p�	>��b����<��զ�<�>%T�]�=e��O���ׄ��ۇ=!�Z;���=�;�<8c7>��ս�-�=�:P� .&����=0)����L�>E|.=şE=l�>[��)?üŲ�<�^�=���γ�=�b��[�=��!>BҘ�����y<Э���>�ɺ��D<���=u�%>������n\=��=�6�����v��_h߽�M=�ͽ��.UI�fON�B�H>��Y>��=`�>�
]�N!�=I�=�̀�Xh���$ <�tX>,�	=T�H����=�vp�7<�=��>ok=�=~v�> v�=��=l4E�	�G�X&>A�<H�`=v�2>��+>N��ߴ!�16��M%����cJ����Hg�=G'>��A���սZe>�̰���ӽx{&>R�=,I�=ܭ>��<�#:��>H�<4�$�4�%<���Opn����=�+�=�<�Q>`]���>��L����=&Tj>(ݽ=?�;ʕQ���=��!�-D��$�Mt'>�턽�$�"������<6m������w3>�"[������Լ/��<�0��՘�J�>�Esp�R�M��V(>Y����>8䚾�=]�����������6���J> �1��l���M䒼x�q����.�~75=-~J=Z�W����;l�ɽ�=�<?>Cޅ>�*�NW�<~P���W>O̓=�0?>o���ƼP��kJ���0;y#½i4n<[cۻ�.=d��=�[&<*��^��<@&E>�޽F҇���=����{�½���;n��<N��p=&�=�a�;mx�=+��<O�/�������=�z�=g[#>���h�r���f>B� =�L>
)�r`=~��RE��۪
>P�J�x�]� Б>�h\=C�>�l>�=����<��K>���=�l�Ac�f����	��l�=���>81>{��8kʽe�k���<T�%�,Q>�&�=�>v�=4�<=��=��̽�JN��>�3>hQ��	�pd��p��a�[B�<�^��e�U>~(~=a I�jR�i���P ��½���>�=/>0~ɽm�D�Q>;�}��.U���1���>��>>��ʽZ����=^ߓ=�=Ώ��=Z��f�=c�~<,S��Z;��\=��&=��m=��A>b=� Ѻ_����(;��3�33���f>~�<�����QtR<�%��jf �)a�=�H>�OZ=����%��:�0�=K�	��x7��b{>�=o�w=qǅ�eL>N뼯1V>H���>� <�pF<��ὔT=��|��H�<�ɳ��"���'Z>*R��
��=�9�� ���9>�=�G8�KW=��j>�����K�P=R[�)���x�X$�w�E>6�ͽ�x��:Ta�@.�=}��=�!��0>�wt>�=�9/=��=�Kּ�<�ؙܽ����=����$>�!��� >�be���a=�B��<;�E�>�'��=�=�Ed>޾f�]�Ӽ<L�^ �c�M>�:=��;	[#>�ID��짽|�<96���2����=�ć=������<+ɼ,�/=tuu��%�ۮ��4�z<���i�>�p�>,.�H<�=R�=��=�+>����숽�C_=�	��tl=Sw�0N�=2^~����=��@<�AJ�!�W>��=��ɽDK�m.z=���<w�	��S�=:~�o�[>SS�=������=��z�! ��S��T��=��u��1��9���U��B>�\��=A�>y�;?�����f3V��m��D�=�Cn>�̔�v_�=� =��=�Ű;�$ <N� �z,ƽr����=��=��=�O|<Ξ꼇�ӑ9�I]��)>׳W;��a��kK��!kf>,�N�_�4�p:,�P<����&�a;�����<�8+��<>^��y��,>s5���
>�KY=�N>�l��]X�=3��Y<^\�>�O=�˃�-���X`��k�=#|���s���K>�����)����>�1<H�=
�>��X=$ؓ=c�;>�>tq>��a=`-2�4��=
n�J$�<-�>L�>��/>��=� U�����6�=�]{<���	��qf1���� j�����=?�*����=��R��[E<31�D�X}��꽨Z=�Ɛ��-b>�g ��QQ>	�����O�=zs�=��A�0üF�f>�w�=�=-�3=�M>���=c?'��(=���9�=#�J=�G�=�>�=k:�<^ƽkxX�e�����=7>�$0��>4����4렽{j�>�=G�����>g�>?������0мk��=�K>��!>�΍<�/��O�=��l�?<cQ*>)f����}>Z>s;=�>M <y����iz>�9>e�$>��<O�"=�ӏ�˯����<�q��bf=|C�=������o>�0��
�<d�+����==������a������=2>��>�ۼ���:�$>_��>QZ��Bm>҇9�#C����=9�`��S�:K	��[ݽ�=��_���c>�^p��1�E2���C
��1!=y���ʩ=k�Ļ%1�?`&��y�=vb8���<��W�� �<QS=f=�����㓔��`>P�I�v��=�ꏾ����!L��'�>�&>pG����6�?.�<B���V>��=K��������2>ڴ^����<���>M�>*
>�0>q�}��)�n�e=���=i�W>�=�z���1�>�����>��g�N�O��ߩ��u�=��&>[���7�">�a�>�a��&!d�~>[��=M�׾أ��P@���'�ڭ����@�Bsg���N��&���S>0��>Z�>��=MK���+�rZ���.#�r5��? ����;�h<�9�4>$N�>@����I�<z����S7�B�\���o���P��>��<��~�t=��\=��)��3=r���G�>��O>2�>�.�⾞�ӽi�;�J�ѽ*�㻞eL>V|�=�-�=�O�>�z��zh>�c>ZaD�/��=��3=��T�Z��>)�>yN>F٘�8X`��V��֙b>ӌ޽�>6��X�=̾�>I'�"�N>oG�>��>aI(��������>�Ɉ�?K���{��,�޽=� �>nv">�᪽?�>p-�<~����I��
�+��`g��}�>�v���_�>�ѾLw>��>�$�#��=)�>�Z�8h�>K�&>�F��b���
�>��q��>��>�N���=>�TkU�ۀ��c`9�u>�=0(����=0�Y���,=����|�j`���M3�,4o�2K�>����#>D��[�>$��ʗ��Zl>�E��j�=p��:+#>�K>�	>=+=v>�|�=�<p<|^>/��R��-`#�C�
��8O��!J�������4i�1_>n�>�;�����g���og�ʌ�<��
=Z�&��g��9 ҽ��>�|N��.�=�*��H7>�聾��O=���ݒw����!�׽s�/�5����,���,������L���=���=n�v���Z��+>�M�=AK�>��(��d��D�0�O�8���W\>�e�=�YG�0��=�џ�4��=���>���<�ł�����p��> ��>#ǆ>��C�⯧���;aa>0����н�v>F�=�X�>x]����=^.A���X����>G$>�zL=>�>���=�:;�~N�>Ю3>,�>Ʉ�̜	>��t�X&�>�)��(���#�Ë�=���<����rI����=�0ʾc�ҽp-�!�-?#&���.���R>��f�>"�t=E�����>s��;�RA=�K���d>�Y�%>`�|��t�=7ӂ=����B����(�_ڼ�W�C>�E��>&<��� �����=慡��ʽZ�h>9��=��=Ɣ6�!������>�?���=C�)?��>E�i����;=!>ݥ�=�¾��R=$�p=*�1=�\½����4��b�a�Ւ��k��=3���79�=ҧm���\��l�>�Gþ���3*�<w¾Z⸽�"%�e����se>8��>��׾�Ct���=���>�Ӣ�
W�=�E潫/���a��;����H=��>;^A=Rӳ��>��L���=y�=���7����>���>T�㾸|�=:I�>n�(�h�1��G�����(��=ty�����:�v��ڶ9>�*8>Vs����X>j-Y���>[r>Jq�=_G����(>�^�=�^���s>�Ċ>�9�=�==���<�#=c=�q�>�Ey�LY�U�ý�g���T��>�"C=��t=(�F>)L=߶=��!�F�>�1�>�.>R�a�9O�>ƾb��Q���D>V���3=>�<"A�<���XG�>��>��7>��;w����=5�V=��>n�� W?�%�<�����D\_��Vr>ܑ>�_G��D}>���u���\u�;�����o}��|>���%�;p/ ����>zg�=,��>X�ľ�B���'�[N9=��?]���P
=+�羇sP���Q>q�">�d�>pŅ�䆀�u_�>�"�=WjT>_�پڌ���>�8W���8���D>[)!�Հ��)=�u$�k�>p�����;��<�����>=7�=A̹<���=�f�=����L�=�)I=�r�=�=̽u8����=���=�x��SF-=�{Y����=�;=�SS��k2<XO�=�9�=���<e܏<�꨽���sO�!J�.�<om)�� ���ȡ=+誼[]y�t�������Z�;E��:q<롺;��X=����0N����[��_�=j�h�y�n=`�:�� *��m�=�����wK�{�3=�2��i����<DB�=ƒ�=��=F\�<��B�Y�>�.��=�4g= X>4�>�5m=ݏ�:��}��<|��<���$�ƽ�M�<}^���	x;�V�<̀Q�.�$� ���=Qk�=BK"=T�5��ϼ��=��ƽ��o<���;�� �ف�=}����=�{�s�<��L=�	߼Dd���+=D��=b� ���{�9�<	��<Ð�0����w<�6��-��V�=ʔ�x�= 爼��;�C�q�¼�)L=��w����<������=���Ӽ=;�<|��="m4=�u��g$=
�4����<���U=�e��z�<#�P�q�`<�2
�&e=�?x=�����=�T
�}#<�@�<g��< ��<�� �y�<
�;���=?<i<#ؒ�ζ6=�)��)��o�:�g��-= ��=�>�<&�<Ä���H��!H<�>/=�m��=���=8\�����=��=�l��nL���5�<NI滺�v=�ߞ=��l=m=V�e<��0=��Թ�ҳ=�,8����=�i =Z����=�e�!{%=��S=��+� &H�a뛽Oj�=f9�,�!��ü2�<�-�iR˼{����S��T>�/�<ɶ=����(3=<ʨ�]���o�x&=Þ=�L����}��}=w��=��-=ռٽ��=AB=���<'��=̝B�'@���<�ɽ�<@��D����ɼ�нS�>o�=f�5���@�|(���΅��$��!�=��=���(>��y���=���*�#x�=�L�<���EQ�=b
��+=��	<��<��;��ؼ!�»����1=�8��RP=�#���D󽼧�<�};=~+"<A	>���R�P��=lJ���s=��i�k=����e=��ҽ:�mjJ���Ƚp������s&�2��<���H$ѽ�U��[0��ڢ����w=�G�<$Wb���˽��=˽�)��Y��K񯽝x=lz&:/�ٽQ�=Pܳ�������&=]�t��7;�=n, ���<~��C��=u�<Q#^���:�*�����E==鈼0ؽ�O׽��H��h;�@�<�����0���>*�=cN�zt�<��='o=����=�<2��=�=�=V��=�z93�
=՘�4��=���<w�;=��M�;���:N�=��<%Jļ���^�= ��ֻ����=/�
�Uý��&�h���I=xr=Ș���=�G�=�O;=���;�?ͼ�T�
�3��4��J��J�;��j<�8T�~c=��<��`�E��=���=!<?��r�<���N�=��� ń��=�<W ���B=��M�Sg���=x����
�Aǀ��d���n�<�� �Zk�< j;���������y�<�φ��T�<�+�<@��@���=��=3��U�==��p�"��Y�P��=��ӆ<T��=)�5=�*4���N=:�кU �0�=�v<~�=�ؙ��j6<�lA|��T�=�%���6-=��P��:��Z�@��s=��>�6=�	������T=�J4=�<��[<h��<b�Y��'�!�?=�=��i��=�M�=�Ԁ�PN�=3p���h��̪<|�*�|����W� y�=g��:�zO���=�P�O�=����֐=���=�{���%>���jQ�='p������}�I��=����;I>��:r�=���D���x>��=���,I��V4�=����wa<��>�����u=�2Z=;;=yq�<��8���<���͟�<ޑؽ�iL����o�Q>X���#�*����=#63<p�߲�;W��;����'ܽ9P-�'�>(�E<5V>�ҵ=��"=t�U>ۼ>�+��G=t��\O���1>�O��>��R��d= �;xS�>=�6�0$f�w��<��6=��:���:�)����c����=<��=WYD>,D��H�=#3@����ּ2=���������9��L�<�6>=�����*�8�^=�x����XV>¾(<�+�=�b_�K�߽�;��<���b>z[��fF���l=�Ie��Vt�1�J>�J=)��b��	;<��z;�?����~�5�S�Һ>����DȽy�v�����>�͇= <�e=�)���3Ž��z�*9=�5>��_=���/�=��^=�����#��,>Cƣ�g����=�H= }(�Mh�=��@�/ǅ;l�={��=& >>,�=6+{<�	>|L�=�n$>v��aT���0>��=ja;��=���>I1=<�$>K�;��Q�h���4?��L��=[X�<캿���`�]���&M��k=��O>t�׼�i��t�;>���h�*4�=f�=�Q�*|�=��=o�罚1��r"1>�P���<"��R�󅡽1�>>���;�����ͼqNA>@q|=P�4>;��<�����Tw=i@h>�z1�TN�������<��нM��=P��	Gn�E�������i���E��(�=��=�>c�U=� x�=���6k�����d�>Z=�;�=��:���=���>4CB�'Z�=󃍼y:�mS-�O��#T�=򗳽�b<�r`�E	>n轉�E=l)�+�)��k(�X�<,[=�N�����;{6��/���e=Y�.<+n>���=х+>{�=�@:>��)��z>%��w�<z�=���\�X���)>/1>D!u=p�����H5>>�>��W��<�O�=Ɛ�� _>LFJ>MQ�ϼO��9<��U>��7��P]���=;D<=�\>Uah�ӭ��]$���C�*?�=K�=����Ka����%�q�=0D��P���Y�=����m� >�kh=�E�����8�r>/��=�:��q��=`9�`�y=<F���z�=��p��h��Ԇ,�f�ý"�a=c=��=^=`���;��8</>��w:n15=�>ݽO��;2�=bC2��G� 3X>�����Ǽp#��=>�<��>���<�>)�F�l�8>��K>�Ct=�3���D>�E�>�ɻ&�w=oo߼���=�<����
����H=>����B�L�߽4�p>�g�=�>�!�<��B=ҥ%����'n�<q�=��r�Hǽ=}���s� >f�����ӽ��5;[�b���=,����=F}�=����נ>;�9<FU�=�����?��_�ϼ薞<˻2=�L�.�<?���<v�d�9(=��>d�=�*�=��Ӽ�;������h;��>CP>{Q���5���=옢=bY�=�H<b�=>��>���=�m����=}~>�߼��<0P�<�͟=ړ�=M�$����=
�>u%�=T�]�A�+�!��>_8l�������=����P�<�-�}?f��6�=~6<}�D<��=���=�������8���e�=�R�=�PC���_������D�����R>�8a>��T>�M�<ܴ�+.���@���νSXk��2�4cֻ�Up��H>rp>�L�:ڊ=�zJ>o'<�o�<�*K�}id=Ja��|�������P�k�>)?�<J>
>.����2+>ע�=�S�=�����D=*������=����ւU�}�A�m�~��=z�<�G�;�F>u��<�=*`�����=( Ｃ�U>0#�[-��&��>�z�:���?��~�=�fs=�?ڻQ᜽x���j���J�=P�<��꼪��R�+}����r����D�;%�z�R>M��c���E��
R<����=X=�Hh�Y=.�#���Ui�=Dr���o�<�<��Qe�=Cr$��r�=�/�<��㽊[��C���u>��c=���=�s�=�����;�����=��"=�>d>lؖ<`����}�=��o��9�=�Fv�u��C(��9Z��C�4\>_B��P�r=�I���n�����`@���>Ph���9>�*=�y�=����~칽<�;P�='4�E{�]�C=a3ռCЙ�E뮼�E>�1@����=�f�=(w>��	�;X�=�;=���=���p�>%gm>��>�YV<ȕ>b�2�y;S�V3>g�߼����=_��=� "������w�
n�"��6=���9�{�����zO=�9�>s&,>�⬽d�7=e=\o	��F�s&� �P����=ө�= ��<!`E>��*����=<R�=�:ԽE{r���ؽr>N���>��w��Y���a>�;ʻj*B��m�߃�=J@>d�����f�f�T=F�`<�8F=`���>����z>���د�{��� )=u��<��ν��>n�A=��2<W���ʽ�;ʱ<ع�K�Žy�}�ݛ�<D��=�x�<M|a��*�=�xY=�n�=
6�hJ���e�=&A;=�����=���<d��=p��=6숻簨=�5��H>���=��M����);�~=К��;	��# v<��8>/��D��(�t=�����T�<�>>����|��fd>�닽uʱ�L���{��L�Ƚ�rǼ#��^S�=ۋ�=H�,=�+u=N�<�� �{�=;��;��<a��=S��
��� =�>��q=��=��X=n�ͽ��|���<���;�f=4��Q�h=n���N�%=��ֽ��=��7=ir�hD'�ip�F�w>ٽY=ƿ���5>�#�<�M<l�=F� =X�P=��=��0�hA��ZN�b$�OA�	>�<��>�d�=�ᕽ��C�V-�=;����ٹ��1>@�*��Ղ�����̗���>�͠�E��=����oý���c�X��/>��
�1{}����]�������Ǉ�=�cҽx��5������ �*�a�)�]>�� �'$6<Y=6?�QK�;�<�=�ʆ=�2$=�c\=��ʽ5K�=ѴY=���#���ݽ^6�]�M�0��N�������=b!��wg������I����8#o<PI�=y ���q<���� =�-=�f�=df�; s�=�#>'a<�' ;2E=b���\=��,=�ˆ=r�<Êν��>>��ӽ��2��]=���<�/���<�:�<iU���A�=H#�<e~>�r&=\�=�>��"=d,����<�t��3g�=L��N*R�K�=& �=��=�y�� �{=�W�|� >�=��&��G�ҽ˥>6��=��=�V=Ogx�	{��j3��t�=���=I�=L�A>����<���>b��:�=���=�� 巼4=42���=kľ��=�j �h�	>\����4�=��d�	�����=S�;<a�\=q����=<����>��=�#p=���i=`�|=��=���=N"�<�>58�=%���b��=���=]�뽢��<]�>Vl=|U�=a��T.k=���=P=�=��/��i>Z?�=����vOԼ��"�(��=[�=��~=6�ݽ�A{��塚��`�>��\�ѼY>��"=�R �ق�=��<B���=�(�};�4�=��m�[Y��M+>P˗�0b�=�8�=��8<}��������t�=rj>[�ýs,�=p����=&)�=��	>�ܟ=��|=�򭽯��t��<��=�5>a�6>nw�=�	��'��,8��A��r��e2<�Sa�Q�=��ؽS�'>OM�M1�=��={&'�);3�Ni��f�ܵ����P&=Y�<��; �ý�2��E�>�F<���=x�'>�S��V�=~�����-��dѽĿ=LO������ ن����*�=� �<�|���	��0�w7�>��O>��̹<D�����ϫy��,�V//>�A>��>R��>FP��V&>��>=�jg�h=V��y>E�:���\<S�n��Ω>�+/��}��!�]�.��>���=�r�>�eܾ��_<�3��{��=un��4*��.�껤�=>;ǾR��=�� �O�_>��D��۽iƾ:˧�7�W=A��d���l����<�8�>dL��$>J3�>!�=����G�G�^z�>4��>��}���=%����y>_4��3>�M�Kв��2=xx���f� ��=!ل=sp��	P@> $���˾^�=[�?��=%k
>�I߽»�>QN)>�&���t�S��=�x��Q�=>v��>��Z���>Gv>�I>���>�ǽ��g>tþv���p��[�=��=ï����˽�7_>8�<f<e>*C�=+���IǸ��N>�ݲ�������j��p�����=��>�Mʼ��澌��=TW��)`���v==�Y���O?�o����=��>���>�']��<�ev�>���{�=�B�(#���0���/�>
|���\<��;z�k�a]�>�Bʽ<�>s����,~��-�c��T�>T���g=rǞ<3�ۺ��>�7����[��+����>�߶q��E�(��>Ql���ɓ=y����|��PY�-�����>]Ǧ<��=��C���>j��=$m��^���.u���<1\�;�����00<��0��Z�>8#�����x�<����^>��>���G�ɽ2p=�䅽�=7�>�Sﻕ!�=�j�=ט>U<�F&>�~�>��=�¾ �(>;�b��>�d��0�Q>4">��
��0��dʒ>�[���d>8	�=�L*�⧉��=N�en���>O��rh=�e�>?��r�T�9���o��:��q/>^{t�{H>|�������Ǳ�υ�=s����7��� �=켁�	��>�8�>��<�i�>j4�>捚;�o>�諒Ǭ�=���=���>��ּ�-��F���gƾ���<����
>�S!�@C>x�t��jj��ľ�?����������:>\���~�=K瞾yi�"�(��lG���O>#ϐ�E�>���'�>T�)�w�	��٩<n��=�D�>��d>Xs�=ν�>[��>A9q�ۥ�>fY��O��[>~;^E���\>~#�<�������=̌����=j1�>�t �z�߻A��=L����*�=Oa�/�>�þZ:��R��w-����N��@$>�dn�-�=V��=5w=�B�!K���aX>�$��l��>o<6>��G�w<(T>ʩ>"��0T�
���|>)�B���8>݌H��-e������㾳����X��)��� 1<�-o�k�>`8���=央�^�>�6��(^J>
�� �#>W70��鿾F����U���5>>�R;B��>�I�>n~��b��gl->*?�����>�:?]\��@ݳ>�UJ>5H>��g��Ŗ=h�>;�>���>(>�R�����ّ�<q����>�����$==p��>Ṿ˥���<�B>�>\��<�O��#.�Ί�>�̢�������=�P@=�Կ>仞�����x >���Ls�>�q�>y�3�Zd�7�>GXn��r=�h��D�'���ƾ�Fx>ە[����6K���=�f�=^�.�R�h>G°�c��>K��3f߽d�>O��(O����>+ϙ�=�>�u�>,�t����Y���R�>��>�wv�.���{
�>�l>w��=L">�dh>O����U�>���|����;�B�����=��>8>�b���^��⁾����;`:0���4=�璽C-|>�w����y�D>�/��^���v�Yo߾���=�ռ��K�>7��=c	0����=/�O���>/0�NL���>!> >*>�b?�o��>CU :��^��Ӧ�h�|���ؽ�>���ŋ�2}��H��y�=��@>#*>��>�Q�zS>P�ϼ�Y��`�;�Yѥ�lқ��=�E��R�=����{��������=��]�n�<�/F<�:Z>����PǾa?}����>%^�<��=�J��(�>�>E־�,�R>����'=H�%>� >�l�<"(U=\r>�C��X�>�?:=�=f�����y�< �>�	-��2�.X���]��*��~�>܎��ww�>�O�'x����;�7B���⾅.	�4�>�q:�]<��h�m�@�G��Ľ7�>Lh�=���Ň��u�=쳹�㵉=y�1�"8��$�~�D{��5g=`b�<�=�=	���S�?�=Ͻ���>�<>��=�0�=Ib1=���=[0�<���>�)ɾ�I�����������=-}���](>"8�PZ�������~=Eg������,�<�gWD>�{�=t��>�8�=��>����7X-���ž$�\�"B콗᯾n��θ�� ������=EG��@�_�
1~�G���bl"���>ܰB�~m&>�I��d�=�� �>:��>}��%n?�V&>'Nq=�I>F�H�z�>��^��7%>`�[�=J�I����Z�>c����5>��t>�A�<�J>�[>����2'c�ۍ��[p��t��y5>Acj����8��_Ҽ=��<,`�X{�>�g�>N��8��>��K<�yc>w�=�V⽛�N<�Y�=uj>
ք��ֻ�|ӽ��P>�>	Eľ�; �|a>�0<�x�<���<7����ٮ>��v�SH�>����W���N��ws>m�k�^��½]n�=rwվ�k�=�j]>����$4��&��a���e>�ɲ���?�̏��)�ʮ3>7��>?��=����|�G��<��I>�>6�X���>Z�=�<"��n==�������w�{�	���>O;=�dӾ������D�(�e����A)�>��=�;�z��k���Q���F���s�#�:>PսU�>��=���=���v�,;V�>�p��o!����=#7�=���<��9>�?s��x>��>�t����ʽ�_{<�H�����<[�O��վ��+>�1 >gH��9+���>�f>�Kν��U>`��坽��u��竾8G2>����ٶz>���9Q���U��<���>P���� �=���g���It����tq���s>��<>�>]P;�)V��	Qw��_�=�z�>�ü�ɉ<�!��v���ݵ�>��>F��Qܗ���=ºȽ���4�5=4n�=wJ��#=�j�=nd�>�\i>�k=�bU���;��]>��=���<|+ڽ��6>�->$*;�f]B��>^���S>o* �9��>�,s��3,>�<``(�u���PJ���A�>��˽����e��>0C�K�m���O���=���>��Խ������o�4�=��=���=|P,>��P�m�>fXz���?>~�׽��>��}��:N>�-$>\oU��Hžy�_�𽀾�\B>��>�b>=�C�=�F�=&��="S>'��=��սh4,��=~��=VU6��Ll�yЂ��m1�*��]>=�v:���>�æ>QÜ�km�w���6>�i�R;��닱=S摾��N>Ş�>�*>>�g��,>��+>�g��w�>�Ѩ��=>�b�=�`�=��F=ʁ�=�w>�J�Z4�=S%&��ȹ>ģ=y,��3+�b`��d��=�A=$�S>?�>����>\��>��M��o���O	>��=d��>�p��+K>ƙD<vcr>��7�ߞT�������o>��>ô���e ��4@>�ԫ=�J$>>�S=/�j�իؽ��hX�����
>s�)< z���5��FX;<�:*\>`~=��4�Ʉ�=�G콰��B�<�Q���ݾ�\�>���>��<�Ǎ>��>�UŽ^��=s��)aH���<p"�2��� ����>Q��=�{D=ɪƽ37
>7G�>ㅽ���=�ڢ��Pܽ�F8>2d��kW;>�ə=�k�=~�>o�0��b>�����]���=�$��9]�>:���u��i	����<g�M>�K�>��>Xt�U#ľ�㚽�s��
MN=>
>�e =W-齒������p4���7c>��>&ܪ<#�ʼ�����>�`�=l\���B�<�\+���> �>$YB���=��=!x�=S�=�:��e���f=��v>3���.�>͒���Q;>�"�� Nl�	*��$�m>�u>L�R��؍<�%�3ǽ����(����>�^��
o��+]>�g�=�[>��8� 甾�#���ą=o�<]NZ>ض
>�y=oPd=X�E����=8)�=�����;o=[���z��(k�^�>�����z�$pR��f�>�z��KNo���������=�����)����;����Yy���ѐ=��>W�� �n>f�<8�l���|��L���r�?=	
.>,�ľ��ӽ2��̉q=����ԣ>/o������C&ܽ.��>�8u��R���r�>��/h �X'<��e��&�=N
v�hyi��T��h�@�@d� ��,�>g_���V>��>Kc"��2��p�P>�(㼗!�>��Z���>��(�O�S��o.��ަ��K>Ւ=����>=S��E��P�Ⱦ#�<�0$�{>0���`=i^M=L����k>2]���I>���>�(ʽ���>��Lp���v��cp`=8 ���u�kN�<u��=���L铽=���[�}��Ȍ=9�:�ft>�V���)�<߃>��-�V}Ͻ/�������B�>�=��b�p��`?��M�>b�>�)�>���=��5>���=���>������>����_�9�� D��L}>%+��v񌾉B>����s> �>0'><����*>�cp>�k=ji<!�����>,����@�Y���aQ5>K�<�1>(z�I��>��>a�0�tNA�����f7��Wr�>�[��������_�<�d���M>l�W��{K����>�Z><F�(|K=dy�=��>>j����Ҹ�G�m>�W�>�͇����3�۽4��;��<>! ����=$�)>��
�>ŬE>^ǽe�.>*#Ž�l���엾M���L>��B�>r�@.�=�0�>nbҽ�S}��\쾕�E>x���,J�� ���o>�"��:��=i�����r� G���.<���>	g��n���>����┾��T==��= f��c���>�ct>TT��{�V��?�=��y��I�21!��ƌ=��=�N�BV>S�>̐,>�>�M\7���P����=d �2B>��)>���>�6�=��M>��M>�w:>I�)�j!�>R�>N�������3�V�u>k�t�bC�g����N��O�=۴��>����3<�>UZ"������>�2L=>�]u=\ռd������;\�4<Ɓ������xQ������D/>�<�,�=��>�&��3g��xL�0\�>>�B>u������i=�b�>hQ�>���=��>/H>��@=����Y��s� ����>�Z��2���>����"?�?�D����=VB���=��=\~>G����*�'i=�܆>��}����z�e>z���3��(i=�_V='�K>�V��[/�br�=#y�>������<�i�>��v�6>�~�>�0㾶�t��v>���=
X���'�>�!�=K�"�S�->[`��Vݾ�E�������>������=q�.��
�=��>Z����<7�@>�Ā���˽t��>n'�>P���9>a��<,��qႾ�ܒ=<O&>"x��17>4�<�Ώ��0�<��5�p�>	���K>X�^����
U>�~�;�����J�>�+����=l[_<F^"�S4$���=m�5<�u-��>�Y��:޾�5�6�)>җ>|��<�Z=v^}>߭>o����R>��҂�>6��=u���,�>ߩ>���>c^[���!>���=�]��=��F���󽃃���9�>��>ȯ�=�*��<�����G(p�oQ*�7�>�����$���>�{�s�P���;�:�ɼ1�>b�/>�dT=�򧾀E�=�e�|��#k>�<�>���*�>u2�>���i�ٽ��=�0�:}���9��q> K���G�>�V�>T�{�A�:>�$I���W�c�`>����R@��_�����>��7> �ƽ��>+P���	��I��T���\��ф�%1�=FW�<�)���>j�2����=���=uJF>���=���={hU�V3��Ʌ��KE>(">��>�*@�(n)�'� �d�s��h?�Gq�*�6_=�k�ؑ��]ն���'������d>ձ�����=0�ѽmVD>f9>��:��r���Z��h ��z�ǽ�୾t�>�>��������W�=^NӾtX��mB��'��z��1��>�+'�5P�	�0���= �C<�I�<Č�>z���O���_��N��>yb>Gr���U�=2r���(>�ʟ� �4<�B�>7����k>P-��)���2>���=1O`<���>:���Se��7B>�Ǒ����;3)Z���">z{>Ј>�+���L�>�T^=.�=K���Vk>ۖ=��퍾tA7>Ns�>���>���Cs�>\���?�输���hW���=������<C�۽7�*�+׾w¾����F�>_d�=���>f=@W4��Ǿ-v�Gg>����\P=��>fW����=\^����=6a�fު�Ċ�>*]�>K�K��<�_��Q}�=�4�.(�=��������~�=�>�>S.�>��V=�|�>4�>YsM��ͽh�0��%=E>ߎ�=��|�S7���W����ܽ1��>��
<�b=��\�-�=������v>'�+=�ؾ�n��1����J=V䞾�*�<�!�>�A�s�����q�+���Ҏ��0�>dh�3K��D"��Ҫ=�O:�,LU��϶�Ԣ=����>���=?��>��C�Hǰ>��,<�U> 	\>h�s����>)/������G���:�>">}��>=2}���*>�s�=��>�Ӗ<��t�3��=�����$>㩾�}>���>���>S��<I}μ�	�=�0~>KԤ>��=��o5�>m܄;�h�>��>|	��?�b>��>�7�>-�	�ys>�>�~��J>>f:>V�g<��<,)A������+پ�i=P�!>/30��xS;�[�<kmX<���>�{�<o8�>ǜ�=.վ�꠽t��>\X��_�L�=�>�i��@x=;�8>O���m���s��=��>(k>���>�'?��žs�<��S���>i'�>��>��L>����=,R,>UUn��I/�x�3>ܽ�`e8�Ff���Ǿ�9�h�SD>Q��m��>�Y���żܮ�Z��>me�Z_;�p��;H�X!����=0׾��F��������+��>g��=�GW�O߾��~>��0>�
	>_s����v����j�|>�iC>��I��Xm��G˾t>d�����>Q.�?ו>�Zm��2>o��>�.8��n<6̲�Sn�>Ǧ�=.��>&��=N�˾�iH>�ʇ�XN�=�h-�Jgb�ǌJ>�ݸ>�k>�?��Q�>��>��> {V>��=�/>�>�=���ʖ>�d9>�~����)=V��~��.�缇G��eF�=[n�=L
>҉w�k��;������>�\�>�����t�=d5��'�>�S{=�ó���Y���ؽ?Җ��>���˥��rý�Խ��>���=ʴ=��C��婾̷��v�轐��l��>Nf�<t�6>t�����>�'>+�&�R�,=�8>�:�=:�=���>�h=�S�=,��4��H�3>�y�=�@]�0qQ����p �`w�>%�l���>�mμ+߸>�M������G�|t:�Vw|����=���\,=q�>���l>���>iq�>l��啾�x=�c��+�=�#�>��=�I��<�>#-���V��i==U�}������\>�d��q{��8��>�&�:����_(P>���4o��P�>ل>W�Ⱦ�^��,�L>�?�WC�>�r�>��=�G�=��?K��B�.#=7X�����:�b>�m�>��>L�9>��=.�_>���:�>�P>F��=�K���|>P(U�r:�>����j�>G��>uP>>$޾ �<�CE��>��1�mM�> �D>��y�{^�>����>�*>���>�-�����!�s�>&c@�%h���\Ž2YG������HM>�u�>;nk>�)��
L��C��c���i�>��=���ΰ>�r�>�&�>�$>NN��i/*>t>�������m�>���>U��=�}�>	�a�0|>p�$>(�"�/>_��V��Sꎾ�>Vա>A½�W����w=V�_��~}>ݮ�>�F�>��/��/��j>�f?녚>3�����>��>�ݡ�4��\���e}a��ٽ��C�T�v>��=�Bk�A��=ꤖ=�8�>����2�>_��=���=���1�b�Fs��
2�>_��>'�ʾ@�@�6C�> :�>�[�>ls>�X׾3B���"�H���b>;�����
 >�ݒ���2�(�%�땾Q��\��u�Lz�<�	�> �J��Ƚ��#��~i=T�>z�I>�SD>�҉��U>�E4�T`�>��r��I�����P�<T�>ޡd=�O_�Hm��>����-U�>)P�=oa>�S^>�&�>$%m>�T׼�4���2a>��>! ��X_��;�޼�x���|�+陽��->k᯽��`>;�>FѾ���>��X����+cX>�=Eҙ��Q>�U�>��6>Nuj>��,>�`>�q�=�*�����{柾;ʁ>�1�>�7�>,	��`-��8�4>��A���0��`�>����b��=�I�|�<pj�����=�}���_>}X�=�2>�u�W7k=5���5w�>y���~>%�x>�4>��<�#5>V������8K��4�=y&K��0[�Lǡ��{��i����=O�>#�,�;dk=f��=<>tt�>���=�oa�~�a��q�>��s=��">t�=�B >��=�㊾]?���>|<��1�Ȓm���þ�M��ӷ=f�>�ق>�Ʌ��p�=�6^�i��;#l��/���>��{>��
�jI>PT����`<��`>H�>m�!��cоS�ξ��>�];�B|M��m�>)�=���>9�G=���=�|Ͼ�*1���d>����j�>�n���*��E>��(��>����x��׾0d��O�=9QN����=�`O<�۷��0��;	r��qԾ�J�=*�޽��k>=Cľ oھ���=��{e�>���>��>s��>Jo�������z�i�>��>%���厾x�>��=����y�>Ցڽ�И�� %�=�>ϕ�>������>�M��Sp�l(�>���>��`�Wc�>���;�pA>�~�=��>��=�}=:ȟ>�ƞ�ޭ�x��>04�>Ma���_���Ll�t��>�� >�Ѿ�!�%M9>��_>}�>>;ݶ=0ľ��^���H>�x�����?s��a�F�r�c�M�<�
=����u|�=%��>ͧ�0���9��Z%>����[�>�J=M8��$?�>=�����>V8>������G>����.����=�Ӿ�@W>d3���2�>�t���2e>�ӣ=�:l=y����1A�8|7���C�M��>A����g>��=�v�>CY_;�e?>�R	�\^>�E>rV��bf�>�-�諂>�˺��N�>ϑO� X���2J>���>�������=Qս�ቼ����@��>=~�� y������i>,ڱ><���&� i>�8L>7�=���>fF�e����>=��>}O��*�>Ds�>
�C�aۛ�5j�=�d>���@��XvK>�D�=�Y�>�]O>���>��>#��=�ө��N���´>1�|�׶{>O�ֽ�'��$RF�M=�=�_G>�������>��j�v����̍=T��>GЍ�� =�*�>P	�W�>��=2��=������c�7���Q��7/�<z����T��M�|�=����̭��!ٽԂ�=	Q�޳���	�=K��>lx&��rf��KE>t�>s�d����>6N���O�=�b.�����VT�=l��=������=�p�=/SL=2N��{�=>}�轵	�p(��#�=���>�"�=���X>ʟv�����a<�1t <J>�˽5Az=۵��P��D���¾=��<��=ԫȾ���>��5=��=~�w����>�`��f!����>\˽���h.=?�=����3�=)�"<�*>��{��>�f>� ����D����U�\2�=:B�F|�A�ϻ�r&�Ñ�&�>2ъ<'����&��x��#��vx{�8,��b�p=g�f�8���&4~�0Y#��K�=(x1�J~�;IQ:�"��$j��M��>��J��8�=������4���>w�R�!$��g�P��y> EK�@�f�eAT�jD>Z6��}9>�zE��������=�ԗ>ҭӾ2���聳=&r$��[��1=�>Q>���@d��:�D��U�=w�#�fu�V������>��'>l����
=�d�>�>�<���>�������"膽7��Kr>Y��$=��2>�?#��.=�
U��R}>0��=)`>�u> �>�s�=���:���<%�=-���ʄ�1`#�?T���V�~u]��<�"u��LC���6���~�I�i�D�1>��c>*�$���T�t�T�m��=�c=���= ޽�Оֽ��~�NH	?|>�fA=յ��jbE��gR=Q�e=��'>^=Ir��~>4��=B8��z>�r�=��>��<>���=���>�����˩>��S���>�w�=+��C�;�qz�> �>6N?��5\>�5��&� �؝�>�>u�Q�=�˘�v2�=X����x>��0>j�E�@7�=��=;f�>2F��`��r�-��=
	�v(��f�W=�������Ks�>g>�'>D-g=���=�:a>����e�����!���b���=�����=p�>�qa� u�>��=toq��$�<�X�����=l6Q>�qM>+M����s>{�8����i��=��C>��;>���<�`����s��2�J���=>�k���:�� N=k�|>��S�ǉľ?�~>ƫ=���x�$�{����=���=���=n�{�ˋ�=���=P�Z��^�E.���	�I>�<-=J�'�&�z�ɧ�>4�B�z:[�F�<c�=ȿ�����>To>����n��4
%=<��<�f=�z�=�#�>Zn2>��M���o���=>ľ>��>(ۋ>�]���Fھ��[��a=����2�۽�6��ͬ�>���yw���>��>��	>��\�KG����/Ӆ>�Y+�y�:�߄�=(�	>����a�>[a�q�!>�<��.�m�v���\-��,z��������;M|�ᓈ=5�5>���>�}>��#>�T/��Ř�,C�x�>�-�=�ժ�L�>#x!;���<��*>�B�>��:���������������g��%��.�"|l�Z�=m�>}P>��=���=+�:>�Ġ>p(O�A!�Xe��	�$����M�=�
Y>@Oa�t>�V`��5J>�뙾/K�>6��j�~���S��u���7�	�½^���An��%Y>m[�>���>��սяܾ��P>�(���R�=���̽�K�>���=�
�.�5���������5=����F+���>�=�>~��=���=�el=��;��6+/=���> x >֘���̀��p>�'J>ٳ�y#
>���>t�=�T>��շ[>�Y��iH=| >�i�>=�=���=����k{>1톾Du�.A�=诋>\<�B�=�	�죢>�`�>D現_b�=���<���H4>�[�=��ٽ���=��<iĸ�.���̿���	�k��<5c�H�.>ƿ��a���=�>�V9��=Լ�����y�>O؍=� N�]轰����>t���=����gP��b�=����bO����_>�b����ֽ�ྼ~;&F��K��=�Qt��;g�F��>&����ғ>8�ĽWRY����=m��Mݬ>oZ���L=B[�=�A�����!O>��>X���i�=��>w"���M��:�=��>�ɽ|:�=3+Z=W[=F��V���A���ݾ�B`>��T>O�=�8�>FN޽��>;hy�?�>��>�q�>\��=l�>9W�m�h>����A]"�q|a�?�9���YeD�F�ɾ���1�����ڤj=@�˻�0'>$�.�V:)>ے>C�|�>Կ�=�$=-��TuZ>�C��1t="g��w���]��d���F�B�e<x�>1/�=���=���>rP��H�P>V���?��!ؼBԮ>%����\=�����ߋ���
��͡�56h>hG�<�Ǣ��A�����)=�H����>n?��W<���<+�>��w�%������(��X'=��+>u����?<�C=�^��=���>�۾J���u>
�=�$�=��4D>5�L�I�<��z>�#$�}�!�-�E>G6��j:%>a����F˾�<�>QG�:y�<��ނ�����7>�����%Ľs���7�=aߔ>Pv>7�>�^I>Ao�=�ח�	������Z�=�:�=9Mt>�n>m�`�D�a=�Bg��¬�=_U='�>�*��;#>E�>gӅ>�¼��I>ed�>D����SL>|)v��װ>�o�!�>qf�>��B��ͥ��p>�c>9`�;K1��h�35@>��>\u�;$ۼ�@�>�?�<�8�=rp>����=�pS>��2�})�6
�=G6>���=��E��r=/N>
�>�V�>�U���V�=
vN��Ŀ���A>ȧ>��>�V�>��g�%ܼ���=����v�<���d�>��=)Bq>���<����逼p!?>*g+��h��Ip�=���>���=8�>h�v>�n>ѭj>І8��A>��k<�#>� =>��>�3h>�_�N�g>����_^�=�Ͻ�������=4�=�L��ѯ>�#�=,D�>��@=�/��R&�=tSB��@��w�=Н�=�В�d�~<��O�X&���9����~��=G��؎	��C�=�����<�ʔ�������W�����7�E��Wþl�P�2�>��>D2#�?d>��޽�!�=/id=�:�>域=���=%��=g�ҽed�t􁽴��C)�����;�>���=g.f����=݃���"������	�>�D�=b������<Wڀ>�;5�s�>>�U{�&��K���A�2�U>�F�O����\k?��=��d>Y���U����=d}=dꚾ�ټn�,>���JE>�^>GL�&d�ؙ�=�qr>g}F=��%>�>(-��=$,�<�#���S�,|ǽ��&>���=)�d��N� �E�&+�<�D>/��=���;��>N5���,>��<���>� �>�n�>�,k= �1�]>嘆�BT�=�>w��<zH�>D�G>2�˽�O�ED=>��-�>���h?>4��=I��<4?��eMh>bGV���_�x�k>�^k�����onཚ��ó���>�/'�bj�=\���G2��'���ZO�E��>1P��M�a����}>Z���h{�>�g"���>�����<��oP���V���v�=�5>�=4>��G>�C�P�	��N
�2n�>��>�Q�>�֑=�mr=�E��F�4>����.q�c�����~=��w�E(�=a���uJ	>�u�0�H>���>{�^�x#�=I�=��>��=�]��5�,>�#=�>bI�� �=lI���~�=�lK>gA�=�cν��"����Ӄ>?,n>���9	�</҂>\*���=��J�EJ���zF�J]>�B >f��=�W�=��<%�>�J�>��>:�>ݪ���C<���=�н���<�y��7�v���-�<���50��Q��EC�rh���AX�ު��.���b�>c9<J��=F�>@2��t��sչ=$�D����>�f>��P>S|>2�=<�u�Lb=�o�=/�=B���wo`=P녾�ż����N�¾cF�����i�^��W�x��т��N�>�ۘ>�s%��#r(�"Y6>0ׇ>��3=����G4�>�3T>`葾*-.>�.����(>�H2>��C�Mx��İo>tw�=�#P�k��>"T^����>���=)�=���=���<p��<.>�q�>��n�� ���ݾ���?�>��>S>.&�<�d��1��?�3>]Iݾ���> 7�^H>vw�>Ҫf���޽e�v>�8�=[r�жB���8>�/���tM=��
����@��>��>P9f>ޫ�>eV(�A8����e>	.��w�>۪6�%��>ܽ����;>PL���D)>��������~���'�Ӹ�=�P�>��>)��̮�>rt�B(������_>gQ�;��ۼ��c��?=XN��SI��7о�У>e���l��=�=r�3�>[J�=�fx��٢=&�꾖��>�/����d>,4�o��>7�;�>s�4S7>�Ǩ�(��=(e�=u�q���=
P<��������_���������=�d��,%�>�@�y�����>�ҩ>o8@�eF�i�<��u>�V�p>#��p��:%O�t�F��/%>��Z>3p���t=e�-��J�o>�3|�>������v>7���A޶�� �>��F��1�>~-���D�<�p��Xo�mȀ�9�G��HH�W,Ƚ���=�]>:�>�#i�'�Y�n>����s�x>m>�˒��P7���o�>��W��f�
��;�Z=/��g\;�ʒ��i��ՋL>��U>#��5������>]�N�C$!�P�E>ÒQ���=�Nþ��=�?�< *��u�5=uU��҃=�/k=��>�i��W�=>v�=b(������2͠� �=��>>��>0u>$������=��>,���*<�l��;4�&����;�$�>�遾[y=_�=�>*G=aֽ�M*>뮱�r���ӵ���b=9X�>Ƴ/� �m���>�i=q�8����/,�=̿y<K��j�>_�m����q*`>;>�=�H�=Y^��{���y�_=�M�>�M�=�&�=�s����a>� ��!4c=�J%�� ǽ
�.>J�|��߰����=�i0��˛�+K���ټ���=Kg�����<�
�'��<eDѾ�b�=��>'s`�`�=��>(�T��|�>�=t��m!>՝�2y�>����G����H�p����>�Ƕ=�m>�擾��=��p����>~h=�V6>ҕ�>��>�~ͽ��>��>qf��i?�="���	Ͼ�$J>uI=���=�_>���`��=�Ž��j>U������K=�1��b�=C�	>�">Vb���9>��L>ax��;]>���=V9��U���Qc>	m2>Ё8���=��&>�b�<���>z���
��ŏ���^�:���و�F��q��lR����$=\�l�+Z��Ģ�=�te=���c}q��>>��>��7'�>;|k>-��=��3��'�>P
�>QG[�Х#�ߦ�>���>$�f=�k ��uq��H�>�� �[8�<�!�ޜ���E>�C�='Ǽ��<eY8>�1�>�}>Hhk>&0��b���7U��Rn�=���=*�>,����8̽-�w�����͊>�X���}i�y�3���G��̎�_	�>�>:ԯ�=���@-��s�;>�v�4m�N��;��^�iO>�=�'�>�z&>Kh>=��@��F�<�*Ƚ�>�<�x>��A>�7Q���cZսx\�>����@h�WHｱz�=���}%$>Y�i>�f>8G�=�F>�J>�,��)�Y>�Z��� L�U��}i�=k�q�>�>�g`>�w������/�>��>N$j����,٣�na>��<Yx3����nż=:Ҿ��=N�f��{�c�p�|X_���D=5HI�zC>�4
�ˌ�>0�4��>6��>̍6>�=���k��	�>[�>>+�>*ى���>)j�0�*���ͽ[3�=K<��/�>m-��*�=8x��lƽ�]�>�4���:���P���6��s>�s�>sï>8�>n��;i=o�!>���>g�=�m����;��掾��꼘�X>�8K>_�>���>�z[�Q�M�����@�>g�=9�>�!`�d"�=�lO>��=�9�>�!%��fg>S��m��>�k=�w�9����>�e���� ?�fx=f�*>uT?>;l
>- h��Wq>P�<������>�`�fK���N�xq|>�
��ȥ�>�5r>@�>�!�=am|>G"���L����u>��4~���q��3q��<��*�=�"��T�$>���7Z���6�>�av�~0�>��5��>BG�ggL�>�k��=e�>�D_t�Ws�>����Zr=�t-,���ּ�����	�>�����u�KoL>��>�&5����>�x����>kO����tz#���8>]y��u�E>�9�\��*愾y]����>�~6=ã�>�w5>mp������Xl�>�\�,�=6y��(�>"����O=�b���a>8+��[�<���>����p�U>�Zf>�d9>�[b�q�+�ht�>'6�����A�޾DAQ>�I�>�w�=Dح�����"m���f�#�����Q�Q���.�>��>��>�>`�j>)�ؒ���K>Wǐ>���=����Z�¾x(�=���>�9��|SB=�z� l�>�>>ZB�d��>�d�>�I<�+���=�>�mӾ�ܴ��hϾ��ƾ�)�>���<�;J>��p>�J>/h��#>���'n=��_��q�>�8h�Z�K>�A�>��5��p�>yL�=NY<��2=zc>eb��UV�1E�U�%�F�}>�U=`��<j
�	L5>��羋W���Q��LǄ>��%�ʃo��o= .��(����žɎ]�i�о-�>j7�<ؽ�=S�>�{=���s=#�Y�{���k�	>)�F>k��>��>l��E�j�լ�>:)�>����%��8��#s����"�$F�=��h��˾�"��.��>Ɯ"��Õ�n�0>\KZ����>�C-��� >��=	�8��>�۽{�a>����1�h��mn>�o���j>���>D򙻃�>>�>��#��R��>�<��]>+�	�'΋�W�u<Of�>���� !=R4>ʴ=NF�>���=����C�==��q��!<��e=:�@>%����a�>��Y>�A�<LH+>d��><�N>&��>)Bj����=����Vbw�T?>l��>qSE�¥�=r;�)`��<<PC�	)���#�>�,�����=}O�=��.>Z*>�5�S�m�86�=p:�>��i���
�o"�=�j�>�Z�� �=u:�>�P�=���>�J�;�|�b��>�_��vfľa�����d��V�%נ>#w�p=�V,��VB��@�0���>�]�9}�<!�@>��v)��c�> /5�諭CO�<�M������=l>�f�>�)���:���>��>�7�>7���>����}��C�=DB>S4t���->�*�<��/>�  >l)�:_e��}�?>Z��'lD����>�{�=Ä>�M���\��OX�G���8F�>2`��0*���Wo>�5�>z �^�D>�x���սu��5�>1�;�����̭�J��
>41�=�X��2��>_��1�:_�=��5�!k'>�9�>ZO��i> ��t�=m��������=�� �EU�>߃�=VxW>�D�;��=Ҕ���	=cW�>�hؽmi����>�G��'%?C>mU{�F"��K,>�}>|>�Ke���^=���<�����TW�EBl>'΁�q�*>!�>"XI=]^>
A>��ټ�1�>�ⶾ�Ō�:>��%.�Z����y��޾����-o;�s�=���7m�=<���F�>}�y;I�+�\>R(K>�D�=�_�>q1H>��E�����yk�>y�(����I������p>� >*�>��>@:e�6�;�)�=���=��9�ek��;�6�/�I�z���-�j�I>F��=[}�=m#t��Oq��������8���J����>���4�=����y7���>��	.Ӿ�!��Ù=�_>05S��L>тͽ���>T_׽`h;����J�;	��=�՝�}[?����Y��=ָG��(�=�I���j�w�<�;��L �ن�i��'���Z>��">q��94/>�p�>Ԥ�>�!>��ʾ�،��f��ʽT2\>�N�y�=Y>��T�Fb�>�ո�f�@���>�dR=b��; ��=��^�v�>�����$>V�Y����=>��c�����2�T��=��<�����(n����<d�<�ހ=�@�=���=CN�g�>���a$�����,�=�=<��"�x�4��&>�(���vg����=��i=|��ފu�&V�>��v�7�=�|�=G{ν}�|=,'�=d�����=��>�*"�3+=��{�Xo'>)0t��P�=禍���f�U��u#G��#�>@@N>c�+=Y�6>�q�>~A�>@,?��G�Y�=�+O��0��v����=�  >��<�3>;���&r�<�E0�b=��=�#>�}>*�>�s��u���ٽ�'G�[m>�sJ�D!O�y�=���r3f��GW>R(`;Pr��W���;u�X�����>�mk�n���l�P>�`>��C>	�>�>/>����>��x>%���gC �|ے="
r>�7����=Xe�=L�>��=��`�l�=�Q����=P=�<>g+=�1�<����m�> cx�Q��<�.�A[��6\�=�� =�W@>����{Q�=Bz�>��=*-%>�#Y>S�MR[=���<�a��-�Ѡ�m�m��l=P�=��M˽<:�����X�[�����0=��a>%�	<�ݔ>Z���C�= �.>�����=M��>�X�=��e>���=/���L�=�g�<6�������=~�=��N>�����G�>�+=tA�9t>c�@����=��5=">(��y�=W4"���=����HX=iZ����%���=�G>)�����9�A5�X�=2�l��ȩ�l(K��O)>��>>y�<C~���&@>��:��;��9>�`�>�
+�V�t��D>��Z]>D��=��>v�J�Y`�=��M���*=�ެ;�۽~<?>kr����;��0�k��=���=3�ҽ�<2���E>w,����=��J>�4�;/����� ��ġ��'�>���r)½EZ2>�1���8�m ʾ��>n,7>/~��2=���>�'�=)��;�f_���v��lU>P����~ݽ�ϒ��i>b�
��v>D`=��>m��=�M�<F�c�(>�	��ܼLv���l>�B�j�k>�־?J�=7?>h��_E#>���>Zt�<a��< ;���1>�OܼPZ�=��=?/��V�=8֨=���/���z�<ͷ�=Ւ>����jx󻢂�=������=�нnp>0!4�t3�>�h<s�<�xO=�
��b���K�1=��E�,���SV>£�>/�/>~��=�	�o=�>n"�<�k�>��=|{��t�^���=�B�>]B�<Ш	�����&�<�s�>���=�@��p�[����=�P�>��>$ϐ>���=w���:<�3<�ٜ=���<��N>d<�aq<������� Jq=�o�_5l���߻�9�>�$<.y�>6�q��}p��u��.>��>'	8>�n�˶;���X�	�W<�<Q�>.�N>��4%>��r������^�\�>r��&]�>���o{>.#6>��=��N�>�5���A>���=���f_�<<;3�1�8�ҕԾ��=<	���8� ��=a���:^�K�Խ�ٖ=e��.ֽ�7佩���Ş���Q�:eh��,H���u�<��O"K�{�='䲽����=q񠽉牽�F��Q>~朼0٤<M�C>��*a�=\���=��{=$����3>P[<�!ݽ�;����#�}�= �o;@��<�+V���a=�=�{>�TQ��7�v�y>_�=�C{>d���"�=��2��w����<�Iv���%�����K�-c��p�=�`�>�>�Ek=X��>�Z���{��ޥ �~4���L��I��P[=�۽�t�<F�'>u�=Vn��ѭ�{?2<�=>,{�[uA>͏	=�᡽��>f�����=�H};���=�w>0�`��3�>^^L>h9ʼ���(���z��$}G>#I�d�a>V>\� �F��>�JμJ�߼-���"�H=�\>ي���>�J< ���#���0�>2֯<�������>�އ>^0> 5�E�"=z�>���=���%(�ލY=�{>��y>L�!>��'�84�;"�Y>��>#'�ڈ>�����e>��>u{�>��=�F��z�=YԚ>�Q9>ǚ��Q����=�n�%و�u�������=v�$>&:��e,��K�>'��>`L�>V�)>�c����7>"D�=�O5>�t�>�␾�g�>z����.>�h,<Li;��S�L��s+> g�=��:>궷9�����9g�fA��5�T��3$>�5>��|�a�Y��@�;]]�Qޖ���>W�~>ʃ���Ⱦ��/>�r>\ɛ=�t>>�a�=-oA�O�>9GR���*����m� �\>�\�=m�=}U�=�ɍ>#�Z>����|�q�?��>}ʛ>%��>��b��=>�篽��r�٢Ҿ��?���)>���>� �GD�=�'��M���w��ݡ	>Pd��8D>�l��C&>���_0����N��>�DI�Ys�G�����=�ξ W��_�ve���=>qb>�.�=�B�>_Y]����j"ڽ�c>�~�4��xz��<�>����nK�n�<($8��97��?>�O�jr>^��(Z=�n>:;=dz9>mR���+>3�4��� � >��e���=�">D3޽�����ڳ�s��=�U�<�	��/F�>���>c�>�F�> "�X��-H�=݈>7��:��*�<��4�
��m���6���J>ߨ�,n�&�F��B���b<@�=��=��C�=(ٲ�/�=�f�>z�=ٸؼh5�<�?���,>��>��<�����t��G��/�=u���9>���;�⩽��>K�e=��=�ӎ�1 ���.��]>��i��yA<th��=�楶=�R�=��S�SÜ;�)�"�h>��x�Çk�Y,J�N=U�ֽ��>>Ď�;W���e�[;.�����>�#���a���\����>���=�T>5T>�G[>(�ޟT>@�=;h�&�����=>[�"=q�=W>�-��=��ݽ�&>f�B����>J�=F~�>	0Q>�>^���>��<o$�=��4��=<o$=���=3_�>�>�{>��==ͱu�y�T>�:�=�8�">U��=ſ=��4�k捾�{C>�=��ҽ��J=7�6����(%��y<�_���ZϽ�n���="���αV�Ӫ��k?�=-���j�n�3n�>h'�=�BV>b��>�!N�\FؼH����<�q��Ŗ��bg��f��͂����>|�=��	>����Y#2=󷏾�U#>��<y[>���=W� >�>ZU�>����G�Qx(>��o=�˯>��O>�D��T����>lt����>�����M��D>��u���g��K��vzɾ1�~>%��=\Hn�����>wn����\>��� %6>e�J=����f½\��|k�=C'�����AI�=���>��>9�=����*��:^����)=2�L�<N#m��`����G>{O�/N� �'=V���&j��7����=��>R��><^��X><�Q�>�;>�愾61>��r��C׽�m�=Ƣ>�?�>���=�>��[>#������;�����T>��>�w>�u�>�n����=�0�=�A�>G���� ;�v�� 2�>��=��ڽ���=mI��' ><x��	>�m���>ݼ���N���Y>�A��_4>��=���;7����>�z���W>	���Y�<���=aV�>�����g >�$�>��O��K�>������>=DȾcr�-q$��-���g<�k��=�[~>�2���ŀ=�
޾#��>l�N�o��>;��<X��>��=Ž��i�=5��>��,�|:�>�x�>�[;�wI�>�׎���>[Q@�C�>���>�I���ͽ�i->��g>Sx>{�a���I�XIe���q�uZ�T�=������N�;=\U`�yWd>��u�4�>���>���=����iǽq��O�)�[N�>@i��#�M�*ֶ�����>{Oм��$>�B�aT\����=R
?���?|��%V>��_>@"��\<x<�� ��>|*'����⁻�k��=)nW=<>)X=��9�پ$����-�=S^�<;M����p��<ؽh߽��~>Dj�>�c���_�����]�8>��Խ��?3V>qc��!M�=!S!����>J73>��1>�a>��i�է">T-Q����>����[����v�<9mn����=볽�hP���Kh��,
>���=u �O��=�+6=��<��T�(�Ѿ6�о�p'>����>�>��>�L=e�N�I]�=�~>�qW�q��>��׼���a��>�옽o��>���=�?�$bb���m=�Pq���+�Q��<1��>��L=���>����ؗ���={��Q_�����~�=k5�@L�NRq��{	�]O��L�	�|,<[ʽׯm>���>��>~?'�KD��E߽�d>�aj>i�%� ��=��V>$/�xJս̼�����Ĵ�>�S�<@ ���>�R��y&ϼ�=�86�U1�>�֓�� L������!?�ܐ�~O����>��U��9�>s���Ə>u�>ÉϾ�����B��W0�ߚ$>��W�G5n=��G>n��>��T<�?�/���q�5ӈ��?�=�?�>��k��s��d�>#��O[;>B*��dk��7��>9�=��T>>W>���<j�>��=tp����<g*���ҽ�>>m��=�S`>?m'>늛>��k>�~m���=��Y>�y����>!-5��i>P1z>S�s��s[>,�{>�j���I˼nB�>vP�>�e>���=b�>`3�<f�>��>���>$�k>��*���D�~�����B,���=�꛽]��=4G�>�N�a>P��d�>�����.�ٵi=��Ծ���<?��>�:��.s��J>�A7>�HֽLg%��8�>`%}>�=�>̰�{A�=�G�=�.>���f5���>��>Fվ�KE����>4@#�&�F��@�����L>�0��>�Ok��LȾs�=�>k܁�����h�6>����q�ž}9��{<�� ��=�|���E��><r�=H�>��ݽ�*_��l�>�д>�>�(�>�\x=��S��=T�P>�����3>Ce!�����=T=��Ͼ�&6>|�)>��$��o@>F!�>��<�'�����nF�>����S>�O��6S�@��CSg�TO=�]��	N��1>��>�GI�J����+����Y�=���/�>��S>pJN�"�	?���=3-�>[>W�8,>�U�����=ٚ�=��>���>U'�}��.M=S�T���G�Vݲ>88V�Mgt���=$#���{�=�#C>������<�e>�/ƾz׉��{Y>����]�=�νZ�n<�`�JO>L�x>��s>2T�=I���W`#>�j/=s�>���=pR%��>�{;>�>I-�/�����>:н/�ή(�����?�Y>�X7�.g��j�w5�<X��>�Q�ZE,��j�=mN�E�*>�%��o�e>*�w��m]>�8s�تE�݈#�yN��m~L������;�a>x6��Q�}������yV>S�1�&�����P��Y���L��MM>�־�E>�ɽ=r�=�4}=�	>�F$=(�)��3���ݽp�=&���V=!���͋>@=��ͽ�<ڽQ�B>�C>K��/U�zu�>A�>�s�=ѵ��f)��=�������>r��>�]'�͗=�#�>��{>�8�Bh�>��̽��=^k˻���H	�P5�=f��ٕ�=RV|>cB��j�:J΅��ܾ�f>s��Zҁ>b
�-�>^�Y=�4�>�i$���Ǿ!p��=�G=B=;��=���=z��E��$ɛ�$o�>�T��P߽�Q.�P�x>"�L�cx%>�a3�Gd�;�q���^\�>Đ=���>U��Q��?ꩽ�>Ů>���3ӽ�zw�nd;˛�>��Z=����=��Iĉ��H�=-��>�z:>�A,��<�>z�_<��!>s�X>A�">�킽����Q��=�N�=�mf>��z�{�k=v~��lj5>�쀾�ݐ�QD�>i�K��6�=���=[��BDY��M���>PՒ=�W=dڌ>�S>��,=������f_�>���G��y%p>lS���־��s>�l���0=!f=3X�>�Q����F>s僾`x-����=�T>��O�܋8����>�%�=I�O�� �<"z�>��0��˙>��>��=�\]����>f������i>��
>}4y��O>�o�90
�!v�ݽܾy�=���>���R�˻���>��4��BK>���AT==H�t>?ҧ���u�F�Խ��>s~�K@>�
�Nt>��b��0���������9Z>C�v�:�\�y��>�3S��~���B>Gjm�P&>F�_�������=)<zv">�����ߠ>�J��s�=E-Y��2��֤>�La�P��=n��YW>����͌>x��=-�y���N��{>
F߻iL�>�4;��o>��Z=΃*>@w�>.���"�����4��սb�޼��>�ʳ>j�<�^�=22����=h_7�^۲��+>�Z<Le]=�F`��1�=JTK���d�/��$�>ص�=D�>�d>`^�)�<(#�>ހ>x�ʾ/e�<��^����ž�v>5�����e>_�ҽcO�>�@}>�|~�o$��?��۽[���v�������r���=�ۊ=�𽚤v��v(���n����<���>�o���7=�l�<Z��=�>rk�=-��o��=��>8��=�J�=g��<��#�J�,<�4�>��N�v�>_�Y�=d��"mb�R��>Vg�>Jzܾc5�>oIK�]u�=�y7>�͌�z굾�o=Ȳ���9#�cT0>)E<�y�8>����6%>�i��t�=J�9>{^>�����,>E��e�r�0�>zA�X̓>�W{>:�������=�wq�������(��>�>�憾k\��/J!�m��>
�=����b�rn�2�w>�/;��SCͽ���>�$�>�t�=�"��@_��7���^�Ϳ����=�������]/>��O>�������*A��/=��9�x#���߽w��>���>���=�E̾��;>��d>��>��Ƚ�|�>�BH>��h�^���m���:�{=ڀI>��S�f>��j<�0?<m�;>S9s�J`���>G3>Ede=2K��rܽ�	㾚�<�潧��=��N>L�>�Lн�">��>N����`=i�6����;��>�c���<=n�>�T��f���\��>.���>��Ts����g;�-�Q��%�<�=l� ,>Z��=O�y>��A�� Q� z'����K�>o�>槙>/c�>��/�^b"<�K�������af
>�im����>�\�ˌ��:����u>��>b������� �>'Շ>&\t�Gj�|�>�&���7�I�=�=O>*�=QK>�/��FYJ<��q=pe�=�[�z�+���>%f'�X��,J>����Շ�<�����E�=�@>K��>ꬬ�{����>��N>~���K?�W=��\y>-'1>�%?������<����i	=������y̾>)�>a�>�N���v>��h��a���JM<w�m�a�P� ��<��=ʅU>밼>-�(>�o�>� ����������>�y&V>e�e>a��:f%��Pq>�l�:b�=�̽  >{:ּ�I�>o���~q�Cw��E
>���Ԋ==�u>�涽p>�F;��3�<�%=�+s��"�4�I=u->?�O>�Z�m�}��O>擟>K�=�>�<�(>��(�a���t�=�m�>4LQ�Fԟ���>
->�b>������=���T�p��/>�ʐ>o/q�w��=�*a>ࣧ�U������׾)���#k��z{����>G���������>2^�>�{c�O���]�=�����ۻ��[J�ݏI�P�=��3>�w�<"P�<��<.�M>�%���#�3f=`�輒N#�&� �Puk�Dl�>��<�>�>�|>��>��#��ħ>��t>��>5�>��v�'5�𛃾LR�����=����g�Z��=DJ�>�G>�����i}�Y@+>����t��O>W���낝���ƽ��ܾ�c>lP���K����=�7�r4����>�Z�=���ǁ���BO�T#�>"��>�^,>�nC>�.ݾ�n<>��9���-�;��kK��λ���=N�9�B^{=��=o��1U��z��J>O	��P����k>,i����<I��,��=�~>��O>����R�=�#�^u�=4,�>�Ek=��>��ս�ɾx�>��7�m�=�!���a�>H�<Y���:�-=�c>�����b%>�&�k��>4���B��'G/>��>�2����x/�>L����Fs>���>�;>t�"�z/��z�<�O���;�U�þ���>��->������Q82>; �������c���Rc��菽m�>e����?}��)(>�=��-�}k�E�E�>nke��y�����f<*���>��=&�P>��=�.<���>���=\��>������>&�I��0�e��=�`�VɄ>��>��>��>��}���N�E��;Y����
>���>��{�-ɷ�qli>9X߾�{�u7�l�>�l̾G^�<�����'�>���=���;��_>�Ʊ>¤���M���v6> ����=�b��k���Ǿ��	�`>@��՛>��I=�Wg���>� �>�>z��>��<ǣ>K����F'>2Ze��믾�T<�T�> :�������Q��T�c���ޜ��z̽oq>�IL<	f>H6�=I�Q��e?���/�
��>��@;E��Ȥ��Pb�R嬽C�l�N��>��>b�ļte/>p+(>��ͽX�e�V>�^����=�������>�6a�%�>W`�|ph=��={>}L�g>c<7巽�U�y>��q=���>��3}���>�y�>Q���%�=��,>�� �R>�G��-�6W�>-��U��l���oV=_�k�$�~[>T�n�� �=��>�Vm���ƾ�=#")=�5�G�S���&�O�L��>!g�=���Ң��0#S��Q���p�>��~=�����j�1y�=o58>�OV>� ��;�>X�>A/�:V�T��P�>�f8>��=�}��y�<	���C��j��>�}>�n�>���=���>��l=)p�>��kư>���d�	�)
B>9*���?���>�0b>֤���=*W	>@���8>P8>wZ2>�Ο�~���[3�^z���L�>+=ui->����X�� !<]�g>��:>!yq>SPX�}��_M>+����>��;3�m��9��}���<����?Ծ���>���<H*�>.��>4>���K�{<�=��:>$4���,����>� 4=@��4�|>�h�>����y�2��*�>1%�_�>0�j��j�>(dӻP�S�u�=%>��r��<��սǤ�>��>;s��0������=��='�=��?�O=�����9=�C&�L�P�>�A=�J�¾��>�w�>��=�!>��=f��Vj���*ѻl�e���_��/�>�7��:->A�:>�d�>�C> m��x1��d��V�>^�+�<m���R�j�H�l��=����<���><����)����>@4�>|o��U$�� �彵��>�Q`>)@�=BJ7���>�&>����ש>6M�>���a$>�c<�X��(�=P��<�C�>�4�=R�����>��ܘ/�e.>�ľ�==>��?���=�ȏ>�7�g�=��Ɍ�>��7>�g>�k>�:ľ�p �~��d����*�I��=Z���+��~�<K�\>ڨ��`t>Vx�>����_�>�Up�������=~�b����=립���>t�¾��;���=��¾�i\���>�`�>���=h��>:PC��T<�8>ŞϼJg�>�g]��X�[7z��X�]��>s+=�t�m釾2�2>�A���~��5D�=��>歗>&/ͼq$�H��=�����0>]m*�5*ﾶI���=���<l\��Ϻ2>@d����_�P׾>�z�>3y#�����Y3$>�a4�<�=��|�F��G8c>�	�Wd7=�#=ya	>`��>���=K<F>�U���2��fo�>�ܓ>D��V��;��>���>�#"�U�>�٬>V�>"8>~$�g�U���>�iZ��|�=�e{��>Bz��c�ҽX�p<�>1��|J��7�=��B>�D>>Bu=8S>��c�^v=��O=�$���ז>���>߹���|>�E:>5ȶ�p�V�>��>_�P>$G�=�0}>��>ё�>�ˎ=��?PPe��:��Ư>�=>��Rڥ=�S=&�L>�go=���t���c�bg���E>��^�v�r$�=����w>8��=/��>rG7=,�>���T���BYS������5�9�>��V��>W|�>�>�[^=w�Dz�>=ʻ���\��о5Z=��.<��7�x{7�;���a솾�kO�c1K=8Ӿ���������=1L�E�+��>,����M>λ��e�>��_>شR>���>$��>�^v��6���p�>�����>bdG�E���#�<���>�=�=��>����>}7E�WϽ�u��\�=<%=m��>=�=
��>���<�w�������{L���p�&>K�þ~��='L�=,�>�
�>�Y��C��*�=u�>������M�"�@>��>�ʡ��5>�����Cǻ�6���̚>�2�>α�>!^>*օ��� =�ݢ���p>с�>f��>"у>=�p��_=�8��>?�B���*�L �>c�5���>^��>[,�;�C<&�B��
*=|�E<�=�<b�罭�H�S>� �<���=���>T�>>6��>Ă�>����b�:���ֽSN`=O��=�&����>^ž�]{��.��OP��U�/A>��>��d��H̼F�> ��j��=	�9�L�¾�d�>s^�<A�S���>�>P��eNo>yO��>�S�<�A>+���Fؽ��|��>�[s��i�=�D�I�=p&�=x>ʽ�V��Y��G��[em�S��>A��\D2��L�ݳ
���$�o�-��ɿ>Ge+�K�"�b
�=�z]���L���/>��$=����WO�����=��H=?��=)�G�𽷭m>VB����>��>@N��������&>~Q;=�!�=
̾�z��3�e<�N+�
y)�z�V��k>���>�R>��A����=�L�<�fO>��������Ⱦ��{>�3.���=��f>粽�弾�\��s�Q�Ҽ>�C�=��=��=P">�������>2�=*>}Kٽ�1��>�z�=T���н�
>k��[��=w�ݽ�B��o\>���]������>&��>��B�"���C�=y�:�7�>AKO�\�ֽ.n>��6����7�24<a�=,�뽂�r�� �=eޞ>��=g�����>�ͷ>��},������ z= ����<�� ���P�"#�>���,Ӻ<#�<5&�=�=v�R>+�>�v]>.5q���=r�>`4���(�=p��R�����Խ�+�_�������<>��O>N�j>�R=��<)��=+*=�����Qp�jӾ)3>�<�>DL�Uܽt�<r�v>�}�>n]V�qG=<IG>�EG=��>��>�?���M>㚉�J�p>�6�=�gP��D>�����>M6>�h@>l�q�����W���a>����+Š����mL���
�<`�>l={Yվ�=@��������=m�ѽ�bX��lU>:�>i�>S��![>��,��~�v4��1u�:��=��پ|=͢߼��=B>Zp >�;H>�G,>����\>:J	�p�=�����>�9������Y�n|�>�/>�0���GW��:�>+��;V#,=�C��?>�>c��=\��=c����NW�7�a����>q,>R�]�  �`jͽ�Y�<:��>rvo����������dZ�b�|>�g4���ὒ<���g>�W[=>l�>�D=��>��䲽L3����=�������>ſ��b�=t�;>�e=�5�#[q>���馋�*�4���>����5>I�{��1�=;$�>��ᾊ��>=�����==�>�"/>T97>%+a�ؗ�=��:���k�=2�2�B��=�*q��g潊E����>���>z��H����,�;u�,�$8�>{� =��>H�1��:սJ�<tL��e�F��VѾ#�y�j[�>��>'謽�c�<�����N���^<>D�;>KV��q�z>.&>��������/�����.=7���4;��; >�f���>D�M>�_l=�&>�tc�ԉ�<�KL��˝�
����Q�>�Ҋ�
@�>dR1>J��>^R8>���=��\�E�,��5�>�i��4(=�%�=�)K�W9��ݐ��
A>��=~���8�=1tJ�~��=��>=,|>vGc=��=D�=�p>`ʗ�?w�</�b�
<�
%�L��<p�<G��O�>�羑�G>*IƼ8�D;ﾝ[?>�0�>H�þ���>?]�>�8����X���#�5�6>| z>7��<����C���w�nq��j�u>��>/gs��q���	?>��=L¼�~��=<��=+0�<�|8>$rI��K5�����������U>:��=��>�X�>��>r#ؽ�;��P����

>m��=c P>҇f��k.���f���㽜l��/�=3�Z>{��(l���:.=Ś�<Z���>�@�=��<��p��;���>`�W=	g׻���=�}">9�<[��>w�=	R�ӌ�=�����H�=�TY>f�={�c���=�����n��?������w�>�/%�R�<��7���,>�����{H>9�[=H�'�y��>^$���X�Ż����>��>9�X��!�ܯD>	�G>��<�&4>څH>\�=u\���>�������:Gc��ڂ>bI�>��F�ƔͽM�->̺0>�3E��#�_�<\{��2�;�=����3\>�e�o,�=�/�<L�d>�k��-�k�����R�=V�>ʚi�xq�=�g>W&����=�؝>�sC��ߺ=��<�\�V�`��`x>^yg�)]����j=�"<pQ2���\����>D��*)I>/9:> g�=�.}����=����8>6��U�&��4�ٟ�KX!��#o>&�=�
���O/��o0>���>�����>�kW>/e�z�v>Ѥ-��=����
���¾�*>2�=e�=$�W�g��6�>/��>���J�=�<v:�>��=�؇>em<� ;�`~��\�;Mr�Y���_=� G�\ہ��A>��a�!�������>m1���\z�b�
�B�^=� ���?�=��!���=��@��<�U,���i=$&���Y">=��s������n>��վ���l�u�V$d>3-��1fC>�q�=$^=�k��G��>[c@���N��$ �y��I�>�;=wn�=�@t=�u�=v�h����=�7E>,b�=L��=��=_ d>���=.!��y<}<���>��d=H./>�RĽ���=�-i��ꅽ8Ȼ�7��FW�9g�;�eS=	���,�>T ���m(�%���X�=3�>�">�]����؞>� ;=vި��:����p>q�&����=���<I�齹|E>��=�3�P觾^;Ⓘ,�s>z�S<�I��	>�z����<��a�R�!>d���׽\>��>+����(>Kዾ�Y�<񬪽yO⽙?�=��v��9P=R��=�Ч��]��_d�H��=�>[� >b]��
�=�`������>�팼�k1>@�����&=���=5ϱ�C��=@v�<�R>5�>X=�v弗8Ƚ�I=���=5�þ�����{'>*A�ˬ�<�=���=��6��Hf����=�x�>�X�lV�=�kH�M�=��y>�1>����j*�c	D��q>�"��d/=�o�x�;�e�<���=�J>��B��Ğ=�?Ǿt�ͽ��>��<�]>����#!>s@>�c>�'��M�<���>�I����x�;>7�~=R�@>W���a�9=z����>�ؐ>(K�=�^�=�~���t���JJ�(�-�\g1�S	,��^J�d�5>HD>��l>�����i���w�c!����C�4�Er�=�a�E.	>J+���ƾ�<��K��SS>K�<=
'ɽ�$=��}>u�/=nA�=�h����>{ɠ>�^�
�3�������n�Dl�<�G>�ͽ6��z $��w��I�����	z���\`>cQz�c�s>WI>��>yc��L^>�~<=]9�,��>3�e�.�>����tʽ�����=E놽��W>d�=����->{�$�7&�d�<RK=<k�����=�ƾ�Q<y���-��yhJ����!:<>�z>r-��g;��@����$�>{��>	jp�����f��>q�$���>|޽�xýW@ �V��>m��w�Ⱦقپڸz�S��=P���ڇ(>�ꂽ����=�<�;�=� �>���>��P�Wѧ>Uq.�l�ǽ����uإ>�}�=>)O�7���㿃<၍�)`>ы�� ���3K��l��^!�s�����>�[�������v��!���)h#���;U��>��>�ψ�̑彅Q>�z�=@>6v<�<��=�f(���:=�0�S�*�ӯ�=�v!>p��<\'��;�=@-ܽ��6��˭��ٲ=�s'�ƌ̽i�+>���=�&��ܯ=�D�1��=f�1>��v�k�>��9Ÿ�@<��pF5���>������\>�&>��=�/�>��!�%�N��g+=����Y��>�<�>��>��ɾ�E�_�)���\���%^��^��J8.>�0��f^���"�����ڷһ�o���`��L +�y�N��A�=@=X�P�>yĽ�a>��@�b�>�˛<��>I�Ҽ~ϐ���=�ȉ=H˳�,>g�4�����>�|o�x:���>�d��pn>��%�&�E��2��<�Y��!}>���>4�.��ް�l���L*�O=� S��J�>q�o>��Ͻc_�<��v>&����>�*���i��5$]=a<���?7�����=���=�zi�nm#�9u>�Į�rc>Jk�>�/���>��L=�f?��Խ�=T�*>J~f>��=���<�8�����>q%�>�C0>ߐ��n�'���=\N�<��~� >z�>����Eھ��j��>��;���+�0��=�9=�
�>���>-�<��w�=�u�<�����}��~H�>͑]��� ���>9qF>Ch��D=�D@=]�>o2X�Ib4>�<��V��~>>�4=O� ��΃��g>�i.�^J�=*�=�{`R�O��<�P=i�n>''�bͬ;м�������O4>���=�>����$-X>�>x�8=�d=���}���
`=���w��B����$�>�	��4,�>/����Q?�矾�����Zr�m�T��ڪ�$Қ>b��SžQ��>[��>lн��*>s>�>]c�>ڿ<�VC���E��\��a!>5X��<J�=K�=n�>/.(��z�>9��<�)�>x���ȸ�S �=��> ���3\���U=C2���>�����zʾ��y>g�h>V'|>�u��j�>,0>^ >Nt����=�e��8�����k=����=� ?XP�:m��Ц���پg/�=2x1�}�ϼ��>oI5>#��egI>R���`A>���>�E<c�x>D޽NN�>��� J���!�ڽ�׾P8j��偾Ր!=S�>�!_��ۅ>��q��`I��r��#)=�T�<I�>zX�>	�x=�H�1�վ\;��ˆS����=�4��{�
>\\�� �Z{���žλ>=[%��1�>�@_>VF����|���.>
Y�>g>�x?��e�߄�>^���T��>�\��s�=Tq\=4� �ː�>m>�h^4�R� >K�>v��>�;�Ѕ>�m>I�2�� Z�ꆂ>�K�>�]ڽ�>����RH^>�|˽"�R�E��;�>�뙾8s:JT��t=�վ�^_�(w���T?>B
�F��;=�<>�H��&�׽�٤>s�ξ�Zq��.	>��>3�q���f�y#����>��>kX�=s�"�ML>j#�Dǧ=����b�>�I�<g��>->I`K�����m>I�a>���>��>��=��g���C>EK�=�P�I��=�T>�X�>��=x���4(�>8:�=�¯�*T����>UmȽ�uG>L\�=��_>8t��󈾤�5�}ʶ��9>��6=0�q�Ʒ:>���}WL���n�S�׾,��=�v��=K����{>X)�QĞ>G{=e}a�`"`>䰖�t[�>�O�>���P�s>l�S>[��=�I"�k�r��č>�`A��O�L0��5�>�� ��6uY>����O�l>/�u�
G>�L>Ȭ=ݖ{�eT>�m�>����d��a�پ��>��>4�˾*p?>�>������>��I>��,�,�'>�m���5�>��!=Ȕ��~tY�'�==��>hÖ��m��X���L��g��>�*P>�P���"�>b�c�p�����>+���H�>�)>Gu�sd�>�x�>ҝw>��KD��&.)>��
�Ld>���,�9�+��	��>���~	���E�=������f��h>^V�e��l��>%���`Y��ֈ>��f��4=F�=�>��	B�=#L���=1��>+5���ϗ���G��*{>{�0>E��������2S��	C���.L�(Fo>�U9�|���'�ѽ ʋ���������0J�f, ���>P��<[Wr����<�G�<4Q�Z>r�ٽ�����ٗ<��o<p���)�{>'�[�p�`ƽ�ܯl;��=:\+��+=���>ގ�=�c�>�G>����y5�=�8�Cm;>w�>Pw����:�O�<�j�>�r��&��?��>*�=�|u�w�9>
���>�.>��n>��>�&�>)��>���>�̾�Jg��kk���=1�
���c=�\�9|H[>�&���>%1�>=���;�����̟����=�rp��S>��̽rU��T�)>��>�R��0>��>�q>20=��5>@!�>�>|�,>�<�=Nj>�)4>l��sYd>nl>l ��b�Ӿ��h��-����ʧ	��tH>�!<���>ZB���o��^%¾��g�ҙ>>�h�襁��?2�佼1->޺�>�p�>0�X>��w>���l����i=ޑ,� ����T�jM¾P�/>D=j=Z�6>���)�׽�7E=1g�> ;�>.��>���<~l�>탾�C�=������>��>q��<zN=��7����>��E����=�O'������>Me�>L����В>*�o>�� ?u����	�:o=�%�=�L�>�b>�#<!�!�>�4�>��h��[�>�~���Z޽NXP��(>��=�Ah��<b>zc���f����>�o:��q*��dn�^�a��Jľ���2��=wߏ��Q������yO|>��>q�����,>&�=���V�nz���y>��i=^xo>A�k�փ��!E>�=�+�>!��,3�Y/�=�>L����A>���=�2>9��<ȓ�>������h>	���{=��կ>,��=w5˾�)r>�<νȾ�>}ʾ��<��p>��>��D�  ]>�6��>ŽȪ�>DJ¾p]X�婫��)F>����n��>1�z>u�=]���S#�>}W!����=���>��@�%z��{5ܼ#嵽n.�>��0>���Eh�>L�->2��"�F���o>yWW>%Ƿ=x�>�2�>�M=X�����/�"}�>Q$�=��*��D>[����ؽ�X'>O/>��L>�!��_#>D��=�	�F�>�ɲ=#�=����ԇ�=��3=�ž�����,�>�UZ=1��8"<��2>���=��>[�s�|���}����n�>fϞ�2 '��j����>v�>k��������>�m�M�>^���uM��
�����>G����휾6v�ȑ�>��D���@���ܹ=�u&>"�@>ͷ>X�M<uL�K>�G��"�=!�X���>>I���V���>`��>�n��qkD<�ꩾ
k�>����f��>�yӼ��Z>��>��{>��l��|X���L;�h��p���FsS��b�>;��>SF!�:R�<u�>�<����=���6$)��i"�JS����I���=h̭�R�4�;8t�n��>�q>s����w�>�?>Mn�bBu>ŋr��iz=ȷL>UL����<�ҕ�;�>�=/{����>^��=�\+>�Ja����<U��i�z=Bs�X�:��o[>� =,��>�饽`˜>���=P't�z�<=�3�>���=m�>2M>�
=��I��ʑ�_�d=LS�|�p>EZ)=r6Z>P�W�1L3���7��>gӥ�в����f>��=>q�v���	����=����č߾^b=�!�=��=4B����_�d���>'�U<�J�<�C߽uΜ��	c��rἫ�;����>�<���=(?��_�>2�����;6
�hߒ> ���Z�����������V�;H���`�>��Ǿ�X2��錾؅=��輴�u��3Ǿ>Kt>���㔊�Y�#�F�r�&yC�{�=%�w>��>%��B�׻?bF��<>�\��*��=E��=����PϽ��Ǿ?���=���>����E���>bZ�����k��dp׾���<�þ��,��=1>��>�v?��&��=j�$����OY����%>�A�yN��K�*>Wɹ���A��%�=RX>��� -4>$�U���I>��þM�޼P�>sn>`7���"��"��#���dX�O;�>� >?����;<#�>w�:�b[�ަ����?=�	��"&�>�h�]r�>2��F�!�Ng׽D����O���R>֊/>��)=���>�p�=��J>�Qe�N�̽&2Ľ���=0$>S�W�W"T<��:>��_���>��Q=��f�>VY�>v%�>�ZW=���B��>�gƾ��ս��<7Q��-�=�uM��F,�r�x��S��%>�	�q�'�W;ӽ��=j&�;�s��|l����>#!A���]>���>��=��?�=.���=�&����������>@~����{���>I?����e����=��>����e��>P~�>��W��~�>������>�o>.š�P�H�R/��؀���c>'��!������lw>o�>��=��>�=�0��^ȳ>8w��ْ����ՠ��/ �:�j����>�|�	 �<:!#>[�i�)��	�:�-�������������SX>f8��;I�>�hн�W��`b<0<I�3�%��>��=ۓ?��i=%�/��>�}�~
>*���m>�{�>���<��<->F�>�f�=OOi�?�S�76��z>{/����ܾ�n��H�>ٜ½�>ϊ�v�+>-,�=>U>�>�Н>�&���$>}~3>R�
��)�>�ڻ>H�=����s>��<G;I�����  >�G��6`�=�_��`/��8d½���>�*k>6�>>_5�>P��>>Ƞ>.i�=L ھ\w>��ͽ�<���=+e�>�Y>J@��ž�Ӽ��l>��>d<6��l�>_�>��q���8�Aْ>v�1>\O�,�˽����=��N>&3�>MTZ>��$��ya>�I�>=��=�)�=�R�=0���>
��I�j>uQ��J���{>s��=dI]>����1��>�������=`��>�F���̽C�����6>A>��&�U�Y��=�r�>��	>�J�>m0�<��>*��>��/>�󽩈<�{����H��H>�������<;�=5���~ӻ��5�=X�=��=���=9�r=�~���|�>��l�,�
>����"���T=7�!�Y���]#��YZ��|K���a>2o��p��=;����=��$�z>����!n�>�U><���jѽ��;>�F�>$-ｲ��>�X=�y>Q��>����\_��&���&Ǽ囝�Il�>u��>������>�+#=��=g_>�S�=+�>���߽�>]����l�
=��R�!{D��߾[����^ƾ�X�ذ�>K�/=6  �;���@��3PN�\4@�R>4��>QϚ>n�_>}�>�Hy�?��8��>S�:>s���ʦ�L����W��F�=[~�<�>��3��Ͳ>�x����K��㊾��ʾ�	�>�N�==�~�O��>93�>@��%�=tM�>蓭=l��>[p�VN��m)�x�.=���M����P���	>u]�׉>��P>/�=���>�( ��*��> ��t�P
����>�y>`��>]z'=�(��z�>
2
>u��56�4�c>û-����UX�>7!��=�u> 6����=����E>���=s[<(T=�k�U���-¸>��T�-���w=�{���=gF����z��G�=bZ#��(s�7�>��3�>�-E���>��V��t�,&�>Xm��>�a5�ܪ>�{]��5��6�E��썼W��>(��>�|�=~��>�I]�AM�>]<�=/��>P#һ㹣>[�������A�V>����0Җ���&����>
�@=��ν�"���*��?�,���0f>���=	M�s�=`��>����񥝽դ��`�l>�������3����|=�]s=�
��=��;�>�I>_�>Nr�>4�>
I<�뽏I�=�G��d�>zY�=��?���Um?>�
A>�e�Wt=G#��Z�2���t�򃮾���>��:>;>%�{>K8>��O>@�>ޛ�>w��B�;}8M������<����=l*h>V��C1�>��¾���>0�.>��}>6PᾺ|�>.�C��(�>B�<;��=T1c>t�?>A�*>Mon�ɭ>��r�{�2>�*㹷��i=Mi>7��<A��=MR>CҐ>�d��Z���,�=M�[�7�2�TK���L�>X�/��M�>�>*�>D�=�C#>�[1���Z>\�T>K�N>�j>X�>�:='г=K�d� ���֢>�.���B���B��Au>}?��r�>�X>גT=#	�<�_v=��q�����A^@�c���𖾪ͥ>W!��05s:��M�ը�%@^>���AO>�'+���=������H�>�{��#v�=!I��(��<X��<"lľ̦�>ߪ�>] ��� G*�V)���A���<�>��)>�ki�m~=|:j>!�����>�a̽���a��<��y,>�	N>�L>y��>5�>=o�>�=+�3���M���V>�L�=�ò�	�<�� �=$.�>
)�=��{=����/n��L>����:C�.,@>AaM>&(���2��.>�_��y2�dOt��⻞/G>�?�����>9�=rs	>˗>F�>�tr��;q����>3���{�<�Bj>ڎ�=N���c��>@w>���՗��w�����K�� =AE,>�j�=Z�U��?=��*>u��=�a�>�ɾ!Bl�9�g=a｛�#>0����z��G�,=����7��ӏ���l��X>{C>�y��#�+>�\>эy<���<�?<>G`˽Z���I��������=f>�`��BwƾA>*7�>5&>wb뾸�սׇ�
�����>z|=>t�������!���D�>[=>�}[��\�f�C��"�Q���|{�����G>^���_��>�,'<�*¼M��=�x������AFV�O��Ǖ��7q��P.>y�'����>���d>@�����=�<ý��=�>��K�̙뼮��r�6��?=�|�<���<i�=ޕ��0�>��3�F�>c8���2�>�H�>�۫>����wv=���I>�U׾O`���<B>$��=�7�C�G>m<;[�">*��/�V�A<3�ɨ�>8½�	K>�!�\?ƾ�=��>�&W>�-ν�r>�?�۹E��M�>�ҽP瑽JD>�F"����RdA=�@f>��(�7݊=�k��t���V��7X�>~�)>��ԾE��=I0=?8.�ţx>j�>.��>��>�x�>�E7>O�̾���<��h>��>ut���k>a(y>�V�<� �=���>�.��5>$�Ͻ�ى����l��=j��Η�>��&=�%�;¥���#>��i������-�=�3�ɴ�P��=M.d>��h��L��Uk���/5�y� ���D��I�o���J
p�J��=~2y�Y̝=�5��in�vH2����=D>��>:N����]��7�=a��=�7���K?B�?5h����9>f� >PEy��*%>@ͩ��eZ>q՚�p�>�D>8>�}>��>?+�=�cA��k���Ž�����HS<��>!��ͷ��	�I>m+>	N>�-�>b�>Ş�=C6�#�J�8=��������&���形�>�M>�X7�D���O׶��g�>9�;�o�E�N>Yu�>���?��>d �<��/>�a��Bi�ib���|s�<">ڨ��4<�>c��>PT�>ocX�YRþ��S=�����ͼ��8>h�j�־��[���]�n��d�"����^>�=�g���i�X>�>�>,x�>y3<��%�9`Y�=�A��HF>�Js�>L�u��7k=^|̽V��O��H�>"�D���=���>Ҙ>�۽>�ט>�N�>Ԇ�������6<S�K>�=��lMA=�ӆ>�ϼ=��->Ϯ@�v�>in���R�#�(���,�ۭ���u�>�z�>^�a��y߼>����g����>�+����>v�A���S��#><�ؾ#��>�$��|�l>4E3>�<���_���<���h?���&>��f��p=��|�9q�>�p��A�>��!9w��/���׈>\܇>ե�������Ӎ�>���%��>$�y���D����>z8پ�7?�����G)~�o�I*�g�̽&=W�����پӇ��X�>V̾��C�$��>'<>J�>�*>��Z>d��=D���_�}�G��=S	U>;@�=@�>���=��pu�� ���Ф�˴��t/�Q;FC�=2g��%��>_��=��Y�gQ�>��?�v2>�í��N����ƾ'��=�ڽ��e��j+>�⭾�D,�Qu�>�;z>{�7��>�Ȋ�iӽm&o����=�A]>7[,���û)�O>�t��J��^X�l�>o<>X��Ru�W3۽�iѽ3쌾��>P|쾋�z>��8>�^>n�0=v_�<pѽ�z���
>d哽r{�����>��ۛ�>�/A��KV���>��*>$�=�}���7�����N<؀>�7�>�>}��oY�c������=D��=�r>�2�����0k=Z�5���W��D�K2i>K�=ȳE=��<+,�����UK�O��>�R�=���τ=����y��>�$�>�_U;�y�>�=���>~@c>�R�=�z0>s����$~>��?W���t�`�ׁ��j�>"b>�`�>Ȏ==M�=�s?�:9?b�A?�/�>9��>�������Z>Y=��� ���c=%rE��L>�_y?�%�>��==H�>�"��XL�.w���=��??I�X>1k��뛾 �ľf=�=�`���Q�z.>������l�c8=��?;|`� ӊ��B�>L�S>���yE6���c��P�`�ͽ��<�8+�-���G~����5?/�����<g��>���i�EtҼ��;���=3�ͽj���ԙ?t�>� ���>�}>���>����P�z�l?��Y��Z�����!�-�>W�M��I^>ic�����>��ƾ��=����Z�CLe>��N=ۈ�����:�����Nh��9�H�*>�_T�-Y�ڛ���mT=lH/?l ����)�0��>sپ���=�>v3h?5�B?iⲾ3m�<��<*飾�gνGH��j>*�7�w�@���>3�$?����f�\>|̽�A���=��=_�����>�#�>:N?�׷�b"�0��XH?� �&r�>�1����>)�>�� ?%�� _Q��v?��E>[v�>�v??;?�B%�:?��!?�� �p��>��>=Y�>N��=^p�7ے�d�>��t>]������!���>��v����>���>�ng>
?�B��~��������>�M]�k>�$�>X�=��=49��t<D�)�̾�r�>� ��ї>�Z��ef?��2?��=2��>�:=�o��S�5>��辙�����}>�c�c�����> �>��ýQ;��dR�z(���b2>*ľ�^O����>4��>"E�V`����2?����F�>���>�b=E��>��?$H�{AO?�u�N�'>m�;{�?:��=��������u<�.�>����u>6�>����),���>�\���� ?����P.����=�k2?������>L\�>�q>���>�4k�=φ��҈=a,p?['B�=�c�^5?�2>���v��� %뾢^ɾ�F`���>@�t��j�>���4�[�.��~߯>�`�/�5�=�>�#�>?�?�+�>��]=N�7>���=���[:�>�����>����yM�W'=��ؽ��¾q��>�#���9��g�����ܾ'>M�5>
��>_�#�K��&�^��,���`�lh?��=;Ծ[�̾\��H��>�A>���P�>y�'=fe=?H>)�����>DyF�@�=��>۲=�ھ����T�>@H3�\g�=��-�"��p���b�>�>Z��+о{�?g��=9G�`RN>�V�>�U����>���>�13?UA)�ӵ��I��kB�D�<�����vɾ��a>Ɉ?��оw�=Y >�.2��{��0�Ѽ�,�����=p�?���>�������KM?)s�>��>v�z�� ?~��=ï<,�?���>��>��=��?��>m�����>�y��"�>���[ )��&?;�L�{*��>[�����>�^=�;P�[��Mt>��>�e�> �$>�E�=3�z�%� =�6<M�?�Uт���=�U�>G���5��>7��3'?Z9?���>����G&��ZQ?��R>��$?���8�i_>jt�>m�~=��.=)�>���>&���p�����|�D=q����?.I�>���f��¯��(>@j>�vH?�⽽=	���>t?U�=Z����=�>=kC>�/^>�*f>��>>���!�?Kc?{�ռ�=��f��;�N�<��l�ŷ�~1?����/�#ɾ�?�?o`��.Ŧ�g��O7?�� =m��j��[LC>�w��j�=e����#�>�5��#�>������.�C�O�4��>�׿��aȾgK���E�&[?�\�>M0�>d�c>.p�=�P*>k@	���d���o>*l�`<b0�>�:���+��>���-O˾��T��䐾Tb$?��_����9[��Ht��;��ipܾ�k�>�,����=�����w�����a����j�W��-5��5>I�0�!��=��	��A�v�.=�	<�>����o<��]�?->�Tg>�G�>A�F>�ؖ�ل>r������<�1̾w�+>`u/�X�r=:�>��=�M>�>�8M>�T���=xx��Km�o3��u�=S�i���&f�=d+7�5��=��r=�]y>���>d�޾�~�=$J�=�z���ѽ��}>S��;�M����<���>�����C>Z�_�f��>�vn��g��ៅ�M��}��iЄ����|.�Y��=����+Nݽ��;5�.��"��\�,>3v�<!�弳�&�=5i������<�w���!i�aV�=�w�>ަ�>�O�@���/˾���=��>�	�������7���l->{~d=���%v*>c ���Q�jj<>@�=���1�����L������o>zO ��M�>ЦR�A�=|�>Mz��	���vS����%=�_%�/�[>���*:w>�ñ>��b�V�>�=n���>!?
�L~� 
H>��<�c%�.�7>	�k=~��=��9�=>�+>L�S�Dz>�#����U>k���K�/>�P��Y�|%���?�����/������=���-F$>�K%�Ԥ���=ͽi^�<M'���4j�M�&�f�8�j<w>,�S���>>��ʽh
>-�}>����?q>��v5>yJ��@��=`fj>B�.>��<د<ϟ��=U���2f9�R2��T��>��>�Z�<�E�=�=z">9��=��`����
3 >��*�Ƌ�=J{��\/�>��ݻ��<���<���=��>tC���g`=o>�"F>vh?>�L��1gn������_�0*�<?�b���̽�P<��нl�!=G��>G��>�ܾ��M\��H�e�;>5��>��>�W�=�"�<�^�=�\T>�	��H�>�����D�=
S�)Y�=%��<��f1<c����D�Of��z��m���p�:����.�,�W�E��x�D{���>��N�<F��jr�<j��;�h����>&.'>�>�->1�N�")۽�%��G��>p�:���}>��|��S�ਜ਼>}L�>�]�=���> �>㪩>=|����G>)W?�����#'�=�C�=E`��:�˾�b��h��XTI>TϚ��U>��\��U����>*X=#0'� �=��9=�$->k���2�<��y>}ж>C��L�ҽ�`���N�>�����R>ؽ�\��9">h�A��	����7����=a�o�>#2>�`<�tă>F�>� <cr=)a�����zZK�d�>�=�����5G˽�I�.�>�kn=�>�=��">��ܼ�P>v->�IN>+y<�z�lbI>{s�>����!�>Im�%܊�lc+:E�>��>o4�>�D>�_�>7��=vɾHB��M7�>����ʰ�=�jj�H�����>n��>�@K>���G�N>��=�Z>@��>m�>� E>M�A��!�)i׾��=Q!=�-�=��E>c@(��\�=���<���=T�c���)>�W.={S7>~P�=���;F'���>��V�=
���i|�=l�>8A�>,����Z >o��B#>NM�C_>�">����;=���,�>6�&��-�=(�"=o�<ll>CF=H���Oo>�w�=l]�<@��<��=;�=�/��A�>�z�������'t���<�-K>m7=p盾z�R�z�6�5���%=EuP�f�>1R����>(XZ�k�����4�<'/�=끑=k~.=މϾ��߽�[�=ʍ_>{���`>z;F��L�x��[A�>�F�>�oB���̽���=s����g�<kR=S�њ����W��;�=$,>&���fOE<pd�;������#>�@>i�X���k��f���
���E>��?��Kּ�%�g�>g�w�#=�=O`?V�b>͋�>`Ib>�F,>�VԺ��S��j�=Il
>��Ƚxݽ;X�=�c���M�=f��.�:�1^�`�=�95����<�`=���=�1>\1�=������	�M���G=�RY�\��=�'\=�]�<l�W��R�:��h=A=J��>i0;>�`��ҕ�M��8Sf>�1k�ŝ�=��;�]>��`���p>����EE��w�+=����|4潧Ռ>9�F>�pT�/c8��ѽ䬅���STg>q���c�������/�:��
�ପ�����潭��� @<>��=:�R@�fOX>�aݽ R1��26��ȓ>Ô�����<^�3=I�н� E=ڛ>D��������>�	|=�>G��HB1>��O�:H`>��)����;W��> u*>5�彆/2>ka�>P�ϼ a;�ͨ;[����;>�t �ޠ�=i�Ƚ14Լ�ԇ>�`�>fPu>s9>>���,=Ӿ��9���
�8�k> �&=G/=���=Y�;��.�=�|#>�L�=1Ě>�̵=k�|>E{ʻ߱�=wt>i�Ǿ�¾�䟽Űu>�zK�?����ۼ�g��|o3���i>����=�*���/�;a@�= G"�%�=�(>�d$��]�< �8��>w����p>�_�>�!x=�+>��=!|�7�>�g�~/ɽE\���>��r�=�D��].�]B>6&��f����i=��-�]����*�𞎾��=�y<�M�������=ҁ�=}�	=4���uǾ��>t�;B��=�~��!@�Ɲ��B=2�C�[]=��c��&g=�&�<�l_�É|=��>�~��(�=G'��a#=��T<S**=^(V�K+.�K`��]�߽IX� ��>`�>%,�k;׽��=Spv����=F��<8��>[���i->V�W��o�>��C>��&�	y>��B��)=S�	�4�4���=B$����B��<���&�<V�a>��=�?��ς����νʐ���0�=eT�!m ���=���<uB0<��=�H�.A���Q�>a�>A
q�
hM���6>WK�<@M�9���b�=u�ѽ�'>��Ǻ5/��������9<SO�[Uʽz���w��<H��=�s�=��h> �h�C;w�:m��f�<��o>�1|=�#�=S��X;�=�7 =E�lbU�2�>cЄ��k��4���~$��8����_�ϭj�3��>UF<ʹp���	�����\�=����W�P�(f�=��L>af�`a=߼�=�%<�`2o���+3C>�o
�EU����0����=�]��G�I��W�=W��s�=��7=���<g2[���=�?�;[��Z=.=�A�=6X�=#9~�'����>���<z2�<�&>��<7䫽����9)��2R7��7>�G�=Z�=Y�W>!E�;����D�A>�<�<T�3���<C}�>TS>�#��q�U>�(�;�n=>�� =��>>��<�v�>d�����@��G��=^�u>Zݐ>�#���=��g�"d�=�G=%f	=i�=t�2>��F���������=�LP�^A����B=�;�����</ׂ��D*�9@=>v��u" >m��=������;!�P>�>x��=�J�~�>�/��cA=�.��/>	�:��$=���$� �9LĽ������=-b(<��=F=罶Y��>>���}w>�3�=Đ=���I�>(�=�9�|\@��tH�����c->H){>��ܼ���j#W=��>D�1�U>���c1�Z+���q���Y0>�	�ֽ�K�(��)�=/!�>/���o�n
t�d�I�6�]3,���D=���>�,�{q:�7�h�R�=흦>���=��\���@�%���xx#�d����=��E=�NU����=�"��<���:��3>Jw{��uJ�%��=�̯>Hf��k�.>m�>�	3>����>fL$��׵<����:�ͦ1>;�Y�����M���O���N����>Td�=ʯZ=�>��A�,�ъ8��� �w�;����4<�<�i3�*�H������~@=���=Y���?���>��׾? ʽ�yG�+};�w������L|�=��6�����P<��ER�=�g��߾�����}�=@�>�8	�l�9> �W����<a�>�ڶ>�rW>oyj�I�=�\���X
��k�=�^潛�ν������O>;�����=R��J>���>��%=`+!;��X>}��>w��=F��=vl����Ct����5������<Ə�>5$��n��T7E=Y�?><�!�l�">�+����=�Q��� >(��>Lk�<��;�ܧ�>p��=�J^�����7��=���!3e>��=���> ]Y>ez��M�>�T���O*���<�>���wz>�l>c�=��=����K�>�#t>�>3�>b�>j�-���%>v�T�]�T> <�>Q)�!����ぽ>�<N�Y�'�:���=����Օ��4��u.�=�c)>��-\=�E�<P����������<�ѾOm��$��b"���q=�4�<�ig�,�m����>Nzp�&I�=I�@>�͛>9����#>jhm=D�>��d�<�G>}��2�s>9��=o)�<�Va��Й��/�>1�<�җ�>�>>��7>Y2>~!=�h}���>AՁ=�<�>��#�3��=��>p?�>&�>:���=D��>�]��ת����=��>Օ>Z�2>-�>>Q9þ�

?��%>eBٽ��<
n��g_�=�_�>��;jΙ����>��[=����J�S���ɺ9�<��>��ټ^�|>8ػ�����;4� >�Y>^wͻ5�8�~��k��?*�>�1b�\���N����>�>�!��h96>n4E>�ih��A��?R�U�#�d�Ӟڼm��>'%վ\��>�I>ܞ2��Y�=H�?W�>--���,��VK����u>�6Z=y��>Ϯ>�E��h��ӻ��E�\�dƻ<�.��d�~���.�>뚇�$��>xH�>�P�=j�=Vp���>��o����>���"ӽ>�	���|>d����ga>߃>��>ޓ�>٫g� �>ܑ��	�=h&�=*�!����>%M���=�[�>���>${*=�&�5e�Ij�=5㫽��>�/�>�?�=�Í�C�!���<���\=E���sF��Z�ž��>�c<���>A�\��W�=i�>T�$�&����UT>3�G��ؘ<{�ʼ:�̽=XQ>�D�>+U����=]x\>UtL>Z=�=ep�=��>�j��S7�[o����=�F�}�>�YO=� �=��M�{䒽���>{���p�[> 7e>���>��%>߭ݾ�W��g�h=)�i����&Fu�����N�>�GO>'�x����[BѾR�W���7�S��JZ ��%�A���v��<� �;�J>m��>7镽��ϼ��}�����v>U���G�C���Q�>%���$o�b�M�H�>#���׬���{��ʀ>ߐ�>9S��:> ���<� �;�}�
��^�6\1=8�/>}���%=�Ir�S��<�Ѣ<5�����>��=s->O�>f =;%G��.�� q>������=�(����Ne���1��}#7�6�ɾ�b�2��B�[>!���c�=A�>)]�>oB���z��9���:��>�־!��=#�>��5=_���h��>��>�qS��M�=�F�B�B���v�E�3}��Y<>��8�d�3>	�?�Ĵ	��(�#O�=����@�F=�ɒ>&�+=|2=ģ���I{=��?�Ɇ�>�Z&>GB����̾#|ؼ��D>��<�~|�<����c4Q�S�,��x>�j!>D���Ͻ.w>��>`ρ�n濾4Jܾ�(�=ʿ�=m ��>�>R�h=�S1=��f���Ap>U�> ����>[�P��h�wm����-�,�����<�g�>C�B>��־�EM>\��>���=M͑��Aa>���<8���i����?�[���v>9�	�,��>p�,�o���ө>�Q�>-e�>�$�=��X��1����'�%�
�*>��< m >
�@>I��e��T�ž��l�>F�99���x%k����> �A>�k>�-�>Ȼ�tXg>�ϗ=H�s���}V#�V��=� �5�>����ɽS�=����F�=up=�$&>E��>4i4>�?�<����=*X<-��<�ǁ�?��=N������F��툪<�/��Y�>�=��l>��!>'�<��-w�g��:��>�Ĳ��7�=dn%����<�&��U��f-M>�����f>!���߽6���f?>n�,>S�0�T���@Tǽ���P���1��(�>f�j��	x={�>�,���>�;>E��p��U��=��X=�qսvg>�"i��`�=�]�SM>�>� >�kǾ��b>߾}����;�ؽt�	>�S��ZֽL�>��#��(N����=���=r����>�G>{=$���|U!�Ō��[�=�:>
t���/�<҃'��NH>%4�P�=�$�<�}�<UC<Mɣ>!"c>�|B��vʽ^���T��=&Jo���������=��h>D%B>����I�¼1!�>gӠ�y�<>lI��F�B>�=lQ�>4����2���� >с<�DR>�仗펽YR�=���<�i�=|�=v;F�>I�}�=ʥ-���߽ʪ�;3��<3+��j��>�|��������<�=au�=�W���껼��>�X�=A�>񉍻7@B<�
>c)���	=��a�j��Ў��	;>ü� ��e�ͽ�Y?�o�=��Q��.=���=T�C>�ƽ�}>ܗ�=왊���q>e��=�:R�<F���{�<��#W>ܤf�Խu> ���Z��J��Խ�G>HV�緿>k�=i�>p�v=K\v��)>�
[>�L>�m�=bh>fH>!#�6��z>���<�:�&,���R��/=q�1�<l.>���<��;��<4�c��->��#>1`�=%�f>f4>d">=�ʽ�9,��j��O�>��1>��>zW�>HF����>�̗>�t��=�=�=��R����>(�&�籑�$5�=m>�-��s��<��6�G�=_���d�j���@�=r�y�ڗ=lf�H��=�Ʉ>��$=���g��>�0�;��:�A[=��f>{���rT>{�7�S�=��ؽ���=�{��ʬ#>���dJT���?���=+�>�>2>��X�#I)�m��‾�x>w�=޸�������=��'>�(s<�J��R^��H�= ����C��;��=U�ǽ܉�=fV>�y�=�m1��n>��ǽ4�����=92w>!�%���<����s>C�[�9��H�=�8޻SW>T�ʼH�9��5$�e����(�=�%�h�=�~��â��E�O�i>PR���M�=���=œ��v�>OI���O�=���m>ݏ�SQ>`�=wk	>{�R����<�da=���=YB��ٌ�����>O��>�8���;D�*Gl�aE��"�ܽ�r%��Z�=d�9>���<�X�= �ܽ�3�;�@���uv��G��G�@��>>O�=
�0� r�Wݙ�v�>���=Jd=����ݬO>��>�؜���/>.4>�LϽh}>#�|�����S>N;:�ͨ=Y-�����ӽn��>"�h>Ƌ=K&��?p�%.>"����V>�rR<���1�=�պ=9�= ���A�	�\�&�н���=\�Y>$DS�ɸ�CcR���e���=�`=}�>؟���=4���҈>���=3}{� ����/>(S�I�B��}�>�&�=�;û�P3����;#�=�>q�G�)q�̘�۬�$��>����U������<�}>��F�b{�����=N���u��g���\����۝���μ���)�L���.��=p�D�f�=�|��'罛5��}�=>�������>�p=q3�=;�o�I���8���?ɼ1�R>g�>T��{G��)R�>�v4��Ա=˵�>�=K۾E�Q>�u����&��i��t3�=��W���9;�|��,���Cz>���PK��P� P� PK                     0 checkpoint/data/43FB, ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�����<�,2����c���R�;�W�R�0<�Js��0��i����>��������07���%�����Dtv��A�R�s<����"l��A��k{��̤�_Ⱦ����D����<l�	�f=��9q'�=
Jq�W�2=��<���<%��<��<|��©���*=���<�<	a;Լ=X�Ⱦ��S=6��=��<�<<�������Y����=�ӾPKW@|�   �   PK                      checkpoint/data/5FB ZZZZZZZZZZZZZZZZZZZZZZZZZ]`�3WL4�Am4�`�3}�(4�8�3�4�s�3O��3^k�3;�3l�4��3�c4�d4��4�)�3-�3�f-3�¦3�@3��3]�3��4+�3�O�4��4�K5i��4���4��14�"5uy�4�`34榁4h�3��.5�;�4�#�4��4O�4�P4�=�4a/G4�/5���3(��4 4��4��3�>�3�4)lI4�J�38��3M�3��Y4�+?4U�3n[4��3���4�)�3���3��3��-43��3�U4�Ĉ3|��4�0l3�<f4�aI3�^L4_�_3��3��!46��4�n-4�734)��3ϓ�3��14U��3��3۹3AH<4�&4�[4��3F4s�4�	4���3�Q4�ԋ3�f[4).;3�)�4I3	4
4�!4Z+y4�lB4�k�3-N�3yRr4�i=4���3��24E_;3N�v4�~�3U-4�6�3M4���3�G4Հ3��4��3��+4\5�3[d4ң�3�X�37�4�I�4��h4\%4��3e�p4�^Y4��3��4�]�3���4	J�3u�i4^:�3�˄4+j3�8�4.#�3�*�4��3�l{4� �3���44:v3t�3�)�3�4���3�l"3�93L[4���3کT3�`y3�3E�4�.s3+F'4��q3��4��&3�@4�83	��3nf^3B�4��2E{24�=3���3x\4���4�=�4��3���36O4�p,4葪3Ė�3;�3rv;4��}3�&_4���3�#A4�F�3>�a4���3b;y4p��3��Q4@��3D��4�	�3Y�949�g4!)�4Bȃ4�C�4���3�¦4,[4R�,4�y34u��3���4��'4?,�484�6[4�/�3W�e4ɔ�3�}E4�y�3�405�3��4��3^5/4�x>4��4��94��3l��3	>4}Xk4A�3��4N�3�ť4e��3j�24e��3( 14R�4�6w4��>3앋4_`�3�jR4ӿ�3�2E4� 3ޢ�3#�4�Y41X4{L4	��3(4:�4�A�3R�?4��3x�y4d��3��*4F��3�V 4�i�3�l4n<�3��4y��3��[4͹q3%H4��B3؂ 4��j4m�y4�g24�)4��3���4-��4}��3V$�3q�3�X�4A�3��4�N�3���4t��3��4��X3��4l~:3��34$�3��4C�2k:4?��4ˁ�4��4�4v�94�>�4@��4Ȓ4e��4���3̖�4C��4�" 5�64���4�9)4�ך45�84�$�4E�4��4��F3s�5��<4�3k�34s�3}|�3��33�;�3��3gR3��$3��2�&�3("3��3�=63!��3�_�2��4���2��3n#3�v�3ݧ3��4��3�U4=`5Q�z5��5��>42�4)5���4آ�4���4�J
4ME`5+�c4�=5�e�4K�5D;4|<5a�+4�v5!4<�15��3v�(5�0�3��v4��W4z"5�B�4HUp4r|@4��45��44v�f4C�3P��4�7�3bs�4r�L4K�4��"4��4�4�+5�/ 4GX�4V��3_�5ѕ3��?43�5!V15�~y4�V4Jҵ3� �4)�H4C�w4H�=4m�63*��4�x�3�,m4���3n�o4�޼31��4H�3��4��3n#:4��3�#�4�L�3/�$4���4��4.�4��4. �3��4�К4�X4�E4&]43��4�K�3[47� 4�A�4ί�3�y�4�c�3�.�4mϐ3��4
Dz3�K�4G73F�;4��T4K7�4a�A4��4�`4��4u4�$ 4�"(4�33�-�4�L
4�s4�|�3d,�4��3�v�4�O�3<!�4��3z��4�r�3��4̴�3�4@C�4���4&'u4���4]b�3�C�4նl4
�3��$4���3�5��3z��4�a�4�Ĩ4L'v3�� 5(��3��4���3���4���3��05�-�3���3�:�3�+4�ú3u5�3Ie�3��4��3�3U��3�3�	Z4�:�3�A�3�VZ3�M43c�4�m3ȡ3j/@3��4�g43��{4֣�3ҩ�34˓�4[�*4l�I4��3�Ձ4JW,4c�3Y�H4�/t3��4*�!4�#,4ȧ�3N�E4o�4ňJ4��3:4�Z�3 |4�K�3<��4���3A�'4e"�4���4,�4}�^4�H4=j�4��]4�3�3S�4��4���4�A4�K�4��3Sq�4�4oW�4>/4��4��45��4���3$`5cW
4~�3s�4R�5uR�4T44=94;&�4���4wr�3Y�4y�3� 5���3��4[�4���4e,�3a�4�3��4��3\�4��3�F5ٳW3�h
4!��3�\|4��3Z'4=�3i�*4�I�4���3D)C4[�l3^/�4�R&4~�4�D�3�Q04�.4��d48��3�uW4�P�3THI4[R�3���4��r3j�4x�3�X4��^3��4OO�3xf�3;��3���3nH�3�,?3r�i3=H4�E4�\�3"Y:3̪�3�3:�{3��3��_3���3�.3Id 4�!43�!�3��	4�g�4�� 4��4��3��4���3yn�3���3��v3���3���3qe4 ֽ3Ϗ3��]4#ԗ3�2�3|ۥ3�a�3�]14t,�39�3p�S3��"4�M4+_5��4�ٓ4���3Xox3��3�@34썷318�3�	�3��H4��4���3�9�2��3$��3C�4f^	4^+�3�n�4Bn3��>4[�t3I�4���4��*5)c�4]:�4	�84��47]{4�s�3J��3Gk�3N�74��4	5wO�4YS�3ê4<�44��|4/��3���4��3q�A4�;�3I:�4�/�4ۃ45a>e4�]�4��4�E4T,4�I�4
�4�44��3g}�4�5�4YZ�4B�M3��$4�>04Xx<4�Dx4��3�C�4f�3�4��3�'�3j��3�k/4��3-b�3�C�223�YD3׈4�K373y343�r3�y�3�ˇ3%[3�܋3�jE3�
3��3bfS3|��3�a3/r�3FkA3��{4$j�4/tJ5��?4�4P4F�4�<94«X49ڪ43��34
�3��4�}:4d\74��J4�:�3F=�4�P�3q��3��;4{��3
�4~g!4��)4���3$]�4��4���4%14�@4B��3�O4WF4���4�:�3{�3�@4%=�4�U�4pw4�}4 �4P[4_�3"p�4a��3�x�4��4�9 4x�3ph,4���3L�5ی�3�u!4 Qo3���3���3�44r�3��3"��3��4*�,4��44�+�3��4#��3j^�3�R�3�@3���47��3]��3���3b��3*�3뮌4�~�3�ȝ30�f3��!37�3Ȱ�3cm3��;3�:�3���3
Д3G��3v�'3�^\3��93B�2���3��^3�4b�3c�3Zh
37��3K@4#o4CGA4���3�O�3���3jL�3s�y4��24�V}3��3.9�3
�d4(�3�͸3b]4:��3��3,)�3�:�3���3>�3�Y�3���33��4'^5F0(5�o45e=5���3��4���4ì�5��5K�o4��4�m55�5�Z�4�oJ5�8�4 4뫭4�=�4�a�4�R�4���4�y4��C4�Q�4�[4Qå4Q&J4�)�3q��3=B4�+�4�v�4f<D3XA4��#4Cv^4�x4x?�3�ݍ4��4Z�r38��3�"4�-�3fD-4knH4Ɍ�3G��4o�P5Nvk5
�5Mm�4��3+�4 �4�p�5�Q5a=4�Ă4N�5�5ON�4OѨ4���4�=�4��3�F�4�H�4�Y4���4W�4qUp4��z4J<�4���4�Sx4�0	4�G3F��3�{+4̤4��y4E+�3�}3!�4�tU4���3(#4F�4/��3r;�3c�G4���3ť�3�A,4�)4i�3(��3j��3N4b��3Z8�3���3�H4��3]��3�#�32 M3wϥ3�EV4,��3et�3�kv3�qj40�3��3D��3_�4|":3���3֫�4	i3I ,4�QH4q�M4��3vl�3`l35��3\��3-�4��3-	+3�s�3��04s��3ѷ�31�H3v+;44m�}3`�3O4���3��3�M�4l��3�.Y4M�4_��4���3Ç�3��w3_CP4� �3�4oe�3]e3M�4��L4�4���3C��3�Z�4�i�3��3�64d�t44�m3!��3~P�46ZE3��=4t��4��5f�4�4)�<3E.q4}��3��4�l4.�;3��4؟4�=�3&�4V��3҃4�K
4�R4�hG4��k4O�3pN�3���4��3���3��h4�:5�T�3�L]3�	3F��3r
3v��3�i�3��2,�Y3�M14�Ծ3VR3ާ�2�3i-�3��&3���3�+W3���32�3�	 4`�3���3�3���3��46T�3�n13�^�3FQ�3Xj�3:$�3��F3��3(^48 4�3p/l3���37{�3[�%3S�3��3]2�3�}`3��*4��>3�_]4��39A�3�4�d�3�ݧ3@i�3K$�3�`�3�B�3m�]3��3�3��3. �3+�;3O��3>�`3	3�[|3��h3�M�3�7D3�3t�3�X�3��3W:4�}#42/�3Xn�3�M�3�1�3�$�3��3�kR3g��3�t`4U��3���3]Mq3z��3|�3͍=3䫖3X�4�ٙ3䴪3h 4�W3���3|��3�� 4ز�35��3�3}�3��Y3�d�3��3��2톚3�04q=�3���3+�=3 �3c�3w�p3�Fp3��3���3SOC3H��3�3,S�3��4ŵI4z�4�4��g3���3��3��G4V�]4n�3=-4��4&;�3T4kF�3X>4�4���3�48�#4$P4�?�3�!�4��37Wh5�_T5 76�R�5��5}��5xX�5.�W6��>5'y�5:<�4��6��i5�c�5"r5���5PS�5�W"6T.�4S�>6de5���5m�95��m6�4�47��50�5ܯ;6�<z5&�5�
6W�6��6!R5.9T6+��4~��6tL5��56L>5���6	�:5|D�6��5��6ǻ&5�iZ6��5k��6`��48�75�h5�J*6#�L59��5�:�5��5��6���4|>6�g�4�xt6�=�5[��5z8�4rg�5��5׎+6��5�|96r��4Á6��4��}6���4`�w5i%5�6�́5��F5���50Ҵ5y�6K��4]U�5EО4w�t6l.^5�޿5�@5�l6 (52C66��4��*6Ӏ�4��6���4D˙6�ߋ4k�e5Iw5l/6�`h5���5���5x_6=Po6c�52�5���4(#�6ɯ^5��6���4��U6(�s5[��6y!5~D�6)*5f�>6���4	�6ҁl4�g�536@��6��66��5a�963��6ɻ�6�ֶ5�6��4�T�6�Ɨ5�ˆ6�35b�6�˅5��6���5�A�6��v4�<
6��55^��6�z�4�PS5���5�߆6�x6�*U5X�y5`�$6I�,6�=y5D�75�S�4�\J6@*5���5�5)�6�]�4� 6?l�4�z6A�4��5Pp�4O,6�y�4B|�5|܂5�5���5��r5�F6Ӄa6��6s�]5h�5N*�4�t�6��c5�td6G��4N��6m5L�q6�	�5zT�6΍4^�d6�5�n�6]�4��U5N/`5��5�z�5ZLm5�y6)n	6z](6�`�5��6�4=Z�6 �4�f.6tӂ5�B6�5x1~6�85#4E6��4L�6N�5nxk6D�!5|(5m�5��85�|5y� 5�5��R5Dh�5�C)5�i5���3i��5a�4껙5��4���5�C�4f5u5JD�4?��5Ŧ!4�g�5���4X��5��c4���5��76^��6��6c^6��6[Փ6�'�6�G6�H�6
#5�.7��5��n6܁d5�6��5��6j5���6���5]�D6#��5��7c�5Ιh51�5�fe6��5�5���5_EL6�p]6���5},V6��4"a�6���5�Q6���4a�6,^5�y6�5��6&�5՞�5�c5a�6n�4�5{�,6���6@#�5˒o5 #�5n$�6<�6�+�5��26K�\4���6��5���5��5�hM6I��5�W�6�O5���6�h�4S�	6�e*5��6�ѐ4��b5���5kg�6='�5	&�5d�5u�@6�&6�J5�66�74���6��5]�5�M459�6�%b5po�6� �4?�6�)5�1�5e�"5��6y��4-�&5���50$
6��95L?5��T5T-6��6\%�4"ݮ5�4~�e6�a5J��5�>5=��5L5�Y+6~(�4��Z6
��4R�5{��4ڏ;6I�<4��u5��&5�O�5���5�e5�6d�6ȵ�6�516ȸY4M�6���5oi6�Z�4�}m6�25gz6�05 �6�X�4P�>6j!5��6+0g4O*5��5��5��I5P��4m j5��5�e6�D!5Nn�5�74�t6��u5o��5�s�4�Q�5�1�4�36�ـ4�96d��4)�5 �4��B6Ƒ�4v:5��4���5��5d�I5]��5X�	6�76C"�4��6���3�~�6��k5�P�5^l�4��5"(5mk-6���4�[6���4��5���4Ռ?6��y4vyy5]5x�_5�H5D�;5i�5�#�5�26:uo5��6ϩ64�Sd6��5�5��|4�]�56a>5��6�1�476g�4��5<@5Wi	6y��4A�h5��45�n5��55��g5;�6x'6%�6��4�,6�J4�w�6Rz5�T86}ײ4�-6DW+5�Mg61#5ـ�6�n�4�-*6F��4��6*��4��=5
5b5�5UV5ߌ�5̴�5z6U6T�l6�e5���5�P49e�6{�4&�5v�50�<6n�5��6�A5�;v6�Z�4��6���4w:�6�D�4�,�5��!5X��5��F5�G85�`6�@&6��c6���4��68#4ɞ�6֎n5��6���4�[Y65V�l6*�5��6�`�4���50ѵ4�u�6]�4zS�5���5IV�54��5�ڋ5��5ݪ�5EX6��i5���5�R`4���6��e5.߱5�ڌ5��6( e5�4F6�+5U�6�&5�c�5)�5��W6J��4���5@��5]��5ݍ�55b�5ýh6�:l6��6��Q5V�k6�r�4l�7[Tr5kk`6��5f��6�U+5�1�6��c5���6���4� s6�5��6���4�;V5P�5���5:�d5��5c9�5m��5Ma6��~5�5>��4�RN6*�5�}�5F�5���5>.5�6��5���5s�4��6��4M66$�4PK��ΕL  L  PK                     5 checkpoint/data/6FB1 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     = checkpoint/data/7FB9 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ|�~��N�r�?6��6 ����M58u��)�(6�K��6�o6:�����lMʵf��ls:5���5Ӈ7B�������:��f���i7�s�Du��&���_7,FI��Ь*�����ʪ���+�� X�*0��������d+�'*͓�d�+�M�,Q�<�r��,y�+(:ȫ08����JZ���.���f�,��8"��6��ŶL��+)�����6��/5`�&6�٤6����l��<Y��%����6�S�7�8�d47@���4��i�\6�A7ld5�b)����{�LH�6PK��!,  ,  PK                      checkpoint/data/8FB ZZZZZZZZZZZZZZZZZ��u3{*�4L��3V��3��3GC457�3���34v�3q�3�@4Tmw4`J3��4@1U4�C+412@4��4%@C4⣇3c��3)M40�D4�}4��u�k������/ȷ-�;Ɛ�h��4YeU hY�p�YT<('��J����?�)J�4Az�A�
��Pd�9xC$��5D�O6���5�x�5�"6�f6��5J�?6'�5�l5�X�6�6�gC6��6���5�XH6{i�5�v�5?�5�$6>(6�"'66�5�ދ6���5PKB��,  ,  PK                      checkpoint/data/9FB ZZZZZZZZZZZZZZZZZ @�FPKos�      PK                     < checkpoint/versionFB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ3
PKўgU      PK                    ! / checkpoint/.data/serialization_idFB+ ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ1696559397809954828100142202874921287156PK˵\�(   (   PK          r�?m                       checkpoint/data.pklPK          �=�                   p  checkpoint/byteorderPK          os�                   �  checkpoint/data/0PK          *���D  D               T  checkpoint/data/1PK          W<љ�	  �	               ,  checkpoint/data/10PK          �5���	  �	               T6  checkpoint/data/11PK          os�                   �@  checkpoint/data/12PK          ��˦d   d                A  checkpoint/data/13PK          ��%kd   d                �A  checkpoint/data/14PK          os�                   �B  checkpoint/data/15PK          4�;� �  �              C  checkpoint/data/16PK          w��V �  �              �� checkpoint/data/17PK          os�                   0� checkpoint/data/18PK          H�EP�  �               �� checkpoint/data/19PK           �JD  D               �� checkpoint/data/2PK          ��Q|�  �               �� checkpoint/data/20PK          os�                   � checkpoint/data/21PK          N���  �               T� checkpoint/data/22PK          NR���  �               �� checkpoint/data/23PK          os�                   � checkpoint/data/24PK          D���  �               T� checkpoint/data/25PK          e"ڼ�  �               �� checkpoint/data/26PK          os�                   �� checkpoint/data/27PK          Q���P� P�              T� checkpoint/data/28PK          A.C�P� P�               � checkpoint/data/29PK          os�                   �K checkpoint/data/3PK          os�                   TL checkpoint/data/30PK          ����   �                �L checkpoint/data/31PK          �y��   �                4N checkpoint/data/32PK          ��ED  D               tO checkpoint/data/33PK          V���L  L               f checkpoint/data/34PK          �,  ,               ܃ checkpoint/data/35PK          Y9N�	  �	               |� checkpoint/data/36PK          $�Umd   d                �� checkpoint/data/37PK          ړ�� �  �              t� checkpoint/data/38PK          ">�o�  �               �1 checkpoint/data/39PK          �gHL  L                : checkpoint/data/4PK          l���  �               �W checkpoint/data/40PK          P+���  �                ` checkpoint/data/41PK          ��P� P�              `h checkpoint/data/42PK          W@|�   �                 & checkpoint/data/43PK          ��ΕL  L               t' checkpoint/data/5PK          os�                   E checkpoint/data/6PK          ��!,  ,               �E checkpoint/data/7PK          B��,  ,               <G checkpoint/data/8PK          os�                   �H checkpoint/data/9PK          ўgU                   I checkpoint/versionPK          ˵\�(   (   !             �I checkpoint/.data/serialization_idPK,       -         0       0             8J     PK    @V        PK    0 0   8J   